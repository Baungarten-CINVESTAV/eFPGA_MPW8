magic
tech sky130A
magscale 1 2
timestamp 1672417657
<< viali >>
rect 10333 37281 10367 37315
rect 15485 37281 15519 37315
rect 17141 37281 17175 37315
rect 18153 37281 18187 37315
rect 23673 37281 23707 37315
rect 26341 37281 26375 37315
rect 32321 37281 32355 37315
rect 37473 37281 37507 37315
rect 1593 37213 1627 37247
rect 1869 37213 1903 37247
rect 2881 37213 2915 37247
rect 4169 37213 4203 37247
rect 4629 37213 4663 37247
rect 5549 37213 5583 37247
rect 6561 37213 6595 37247
rect 7849 37213 7883 37247
rect 9873 37213 9907 37247
rect 10609 37213 10643 37247
rect 12357 37213 12391 37247
rect 14289 37213 14323 37247
rect 15761 37213 15795 37247
rect 16957 37213 16991 37247
rect 17969 37213 18003 37247
rect 18613 37213 18647 37247
rect 19993 37213 20027 37247
rect 20729 37213 20763 37247
rect 22201 37213 22235 37247
rect 22661 37213 22695 37247
rect 23489 37213 23523 37247
rect 24593 37213 24627 37247
rect 25329 37213 25363 37247
rect 26157 37213 26191 37247
rect 27169 37213 27203 37247
rect 28089 37213 28123 37247
rect 29193 37213 29227 37247
rect 29745 37213 29779 37247
rect 30665 37213 30699 37247
rect 32597 37213 32631 37247
rect 33609 37213 33643 37247
rect 34897 37213 34931 37247
rect 35725 37213 35759 37247
rect 36369 37213 36403 37247
rect 37749 37213 37783 37247
rect 35909 37145 35943 37179
rect 3065 37077 3099 37111
rect 3985 37077 4019 37111
rect 4813 37077 4847 37111
rect 5365 37077 5399 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 9689 37077 9723 37111
rect 12541 37077 12575 37111
rect 14473 37077 14507 37111
rect 18797 37077 18831 37111
rect 20177 37077 20211 37111
rect 20913 37077 20947 37111
rect 22017 37077 22051 37111
rect 22845 37077 22879 37111
rect 24777 37077 24811 37111
rect 25513 37077 25547 37111
rect 27353 37077 27387 37111
rect 27905 37077 27939 37111
rect 29009 37077 29043 37111
rect 29929 37077 29963 37111
rect 30481 37077 30515 37111
rect 33793 37077 33827 37111
rect 35081 37077 35115 37111
rect 36553 37077 36587 37111
rect 1777 36873 1811 36907
rect 2513 36873 2547 36907
rect 3249 36873 3283 36907
rect 6837 36873 6871 36907
rect 11897 36873 11931 36907
rect 19533 36873 19567 36907
rect 20269 36873 20303 36907
rect 22477 36873 22511 36907
rect 24041 36873 24075 36907
rect 32505 36873 32539 36907
rect 36093 36873 36127 36907
rect 37565 36805 37599 36839
rect 1593 36737 1627 36771
rect 2329 36737 2363 36771
rect 3065 36737 3099 36771
rect 7021 36737 7055 36771
rect 8125 36737 8159 36771
rect 9321 36737 9355 36771
rect 11713 36737 11747 36771
rect 14289 36737 14323 36771
rect 17049 36737 17083 36771
rect 18889 36737 18923 36771
rect 18981 36737 19015 36771
rect 19717 36737 19751 36771
rect 20453 36737 20487 36771
rect 22661 36737 22695 36771
rect 23581 36737 23615 36771
rect 24225 36737 24259 36771
rect 32321 36737 32355 36771
rect 35081 36737 35115 36771
rect 35909 36737 35943 36771
rect 36737 36737 36771 36771
rect 14565 36669 14599 36703
rect 7941 36601 7975 36635
rect 23397 36601 23431 36635
rect 35173 36601 35207 36635
rect 9137 36533 9171 36567
rect 16865 36533 16899 36567
rect 35541 36533 35575 36567
rect 36829 36533 36863 36567
rect 37657 36533 37691 36567
rect 2513 36329 2547 36363
rect 36737 36329 36771 36363
rect 1685 36125 1719 36159
rect 2329 36125 2363 36159
rect 3249 36125 3283 36159
rect 7389 36125 7423 36159
rect 36553 36125 36587 36159
rect 38025 36125 38059 36159
rect 1869 36057 1903 36091
rect 37381 36057 37415 36091
rect 37565 36057 37599 36091
rect 3065 35989 3099 36023
rect 7205 35989 7239 36023
rect 38209 35989 38243 36023
rect 2329 35785 2363 35819
rect 23397 35785 23431 35819
rect 38209 35785 38243 35819
rect 1593 35649 1627 35683
rect 2513 35649 2547 35683
rect 22201 35649 22235 35683
rect 23305 35649 23339 35683
rect 38025 35649 38059 35683
rect 22017 35513 22051 35547
rect 1777 35445 1811 35479
rect 37197 35241 37231 35275
rect 37381 35037 37415 35071
rect 38025 35037 38059 35071
rect 37657 34901 37691 34935
rect 38209 34901 38243 34935
rect 1593 34697 1627 34731
rect 1777 34561 1811 34595
rect 37749 34561 37783 34595
rect 37473 34493 37507 34527
rect 35817 33609 35851 33643
rect 1593 33473 1627 33507
rect 5825 33473 5859 33507
rect 27353 33473 27387 33507
rect 27629 33473 27663 33507
rect 36001 33473 36035 33507
rect 38025 33473 38059 33507
rect 1777 33337 1811 33371
rect 27169 33337 27203 33371
rect 38209 33337 38243 33371
rect 5917 33269 5951 33303
rect 26065 32861 26099 32895
rect 19441 32725 19475 32759
rect 26157 32725 26191 32759
rect 19349 32453 19383 32487
rect 19441 32453 19475 32487
rect 20361 32453 20395 32487
rect 30665 32385 30699 32419
rect 37749 32385 37783 32419
rect 1593 32317 1627 32351
rect 1869 32317 1903 32351
rect 37473 32317 37507 32351
rect 30757 32181 30791 32215
rect 9229 31909 9263 31943
rect 12633 31909 12667 31943
rect 38209 31909 38243 31943
rect 1593 31773 1627 31807
rect 5733 31773 5767 31807
rect 5825 31773 5859 31807
rect 9137 31773 9171 31807
rect 12541 31773 12575 31807
rect 13185 31773 13219 31807
rect 13277 31773 13311 31807
rect 38025 31773 38059 31807
rect 1777 31637 1811 31671
rect 38117 31433 38151 31467
rect 17141 31365 17175 31399
rect 7573 31297 7607 31331
rect 14657 31297 14691 31331
rect 16957 31297 16991 31331
rect 25513 31297 25547 31331
rect 37473 31297 37507 31331
rect 37565 31297 37599 31331
rect 38301 31297 38335 31331
rect 14473 31229 14507 31263
rect 15577 31229 15611 31263
rect 7665 31093 7699 31127
rect 14933 31093 14967 31127
rect 25605 31093 25639 31127
rect 4261 30889 4295 30923
rect 13001 30889 13035 30923
rect 22661 30889 22695 30923
rect 15209 30821 15243 30855
rect 10977 30753 11011 30787
rect 11989 30753 12023 30787
rect 14841 30753 14875 30787
rect 1777 30685 1811 30719
rect 4445 30685 4479 30719
rect 13185 30685 13219 30719
rect 15025 30685 15059 30719
rect 22845 30685 22879 30719
rect 24593 30685 24627 30719
rect 11069 30617 11103 30651
rect 1593 30549 1627 30583
rect 24685 30549 24719 30583
rect 12173 30345 12207 30379
rect 13185 30277 13219 30311
rect 14473 30277 14507 30311
rect 14565 30277 14599 30311
rect 16221 30277 16255 30311
rect 17049 30277 17083 30311
rect 17601 30277 17635 30311
rect 22201 30277 22235 30311
rect 29193 30277 29227 30311
rect 12081 30209 12115 30243
rect 13093 30209 13127 30243
rect 13737 30209 13771 30243
rect 16129 30209 16163 30243
rect 23581 30209 23615 30243
rect 24225 30209 24259 30243
rect 25145 30209 25179 30243
rect 26341 30209 26375 30243
rect 38117 30209 38151 30243
rect 15485 30141 15519 30175
rect 16957 30141 16991 30175
rect 22109 30141 22143 30175
rect 23121 30141 23155 30175
rect 29101 30141 29135 30175
rect 29653 30073 29687 30107
rect 38301 30073 38335 30107
rect 13829 30005 13863 30039
rect 23673 30005 23707 30039
rect 24317 30005 24351 30039
rect 25237 30005 25271 30039
rect 26433 30005 26467 30039
rect 10701 29801 10735 29835
rect 15393 29801 15427 29835
rect 16037 29801 16071 29835
rect 18705 29801 18739 29835
rect 21925 29801 21959 29835
rect 26801 29801 26835 29835
rect 18061 29733 18095 29767
rect 25237 29665 25271 29699
rect 1593 29597 1627 29631
rect 6653 29597 6687 29631
rect 9137 29597 9171 29631
rect 9321 29597 9355 29631
rect 10609 29597 10643 29631
rect 13369 29597 13403 29631
rect 14657 29597 14691 29631
rect 15301 29597 15335 29631
rect 15945 29597 15979 29631
rect 17049 29597 17083 29631
rect 18245 29597 18279 29631
rect 18889 29597 18923 29631
rect 21833 29597 21867 29631
rect 23029 29597 23063 29631
rect 23673 29597 23707 29631
rect 26709 29597 26743 29631
rect 38025 29597 38059 29631
rect 6745 29529 6779 29563
rect 25329 29529 25363 29563
rect 26249 29529 26283 29563
rect 1777 29461 1811 29495
rect 9781 29461 9815 29495
rect 13461 29461 13495 29495
rect 14749 29461 14783 29495
rect 17141 29461 17175 29495
rect 23121 29461 23155 29495
rect 23765 29461 23799 29495
rect 38209 29461 38243 29495
rect 9321 29257 9355 29291
rect 22017 29257 22051 29291
rect 25329 29257 25363 29291
rect 13093 29189 13127 29223
rect 13829 29189 13863 29223
rect 23765 29189 23799 29223
rect 30941 29189 30975 29223
rect 31033 29189 31067 29223
rect 1593 29121 1627 29155
rect 9229 29121 9263 29155
rect 11713 29121 11747 29155
rect 13001 29121 13035 29155
rect 15025 29121 15059 29155
rect 16037 29121 16071 29155
rect 20913 29121 20947 29155
rect 22201 29121 22235 29155
rect 22937 29121 22971 29155
rect 25237 29121 25271 29155
rect 26249 29121 26283 29155
rect 27169 29121 27203 29155
rect 12357 29053 12391 29087
rect 13737 29053 13771 29087
rect 14841 29053 14875 29087
rect 23673 29053 23707 29087
rect 23949 29053 23983 29087
rect 37473 29053 37507 29087
rect 37749 29053 37783 29087
rect 1777 28985 1811 29019
rect 14289 28985 14323 29019
rect 16221 28985 16255 29019
rect 23029 28985 23063 29019
rect 27261 28985 27295 29019
rect 31493 28985 31527 29019
rect 11805 28917 11839 28951
rect 15485 28917 15519 28951
rect 21005 28917 21039 28951
rect 26341 28917 26375 28951
rect 6377 28713 6411 28747
rect 10609 28713 10643 28747
rect 30665 28645 30699 28679
rect 11437 28577 11471 28611
rect 19533 28577 19567 28611
rect 20085 28577 20119 28611
rect 21465 28577 21499 28611
rect 5733 28509 5767 28543
rect 5825 28509 5859 28543
rect 6561 28509 6595 28543
rect 7297 28509 7331 28543
rect 10241 28509 10275 28543
rect 10425 28509 10459 28543
rect 12909 28509 12943 28543
rect 13553 28509 13587 28543
rect 14289 28509 14323 28543
rect 16129 28509 16163 28543
rect 16773 28509 16807 28543
rect 22661 28509 22695 28543
rect 23305 28509 23339 28543
rect 24593 28509 24627 28543
rect 25237 28509 25271 28543
rect 28273 28509 28307 28543
rect 29009 28509 29043 28543
rect 30573 28509 30607 28543
rect 11529 28441 11563 28475
rect 12449 28441 12483 28475
rect 13645 28441 13679 28475
rect 15025 28441 15059 28475
rect 15117 28441 15151 28475
rect 15669 28441 15703 28475
rect 19625 28441 19659 28475
rect 21189 28441 21223 28475
rect 21281 28441 21315 28475
rect 25973 28441 26007 28475
rect 26065 28441 26099 28475
rect 26985 28441 27019 28475
rect 28365 28441 28399 28475
rect 7389 28373 7423 28407
rect 13001 28373 13035 28407
rect 14381 28373 14415 28407
rect 16221 28373 16255 28407
rect 16865 28373 16899 28407
rect 22753 28373 22787 28407
rect 23397 28373 23431 28407
rect 24685 28373 24719 28407
rect 25329 28373 25363 28407
rect 29101 28373 29135 28407
rect 6653 28169 6687 28203
rect 8401 28169 8435 28203
rect 21281 28169 21315 28203
rect 15761 28101 15795 28135
rect 16313 28101 16347 28135
rect 17877 28101 17911 28135
rect 18797 28101 18831 28135
rect 23305 28101 23339 28135
rect 24869 28101 24903 28135
rect 25789 28101 25823 28135
rect 28641 28101 28675 28135
rect 30113 28101 30147 28135
rect 30205 28101 30239 28135
rect 6837 28033 6871 28067
rect 7297 28033 7331 28067
rect 8309 28033 8343 28067
rect 8953 28033 8987 28067
rect 9045 28033 9079 28067
rect 10517 28033 10551 28067
rect 12081 28033 12115 28067
rect 14657 28033 14691 28067
rect 16865 28033 16899 28067
rect 19257 28033 19291 28067
rect 20177 28033 20211 28067
rect 21465 28033 21499 28067
rect 22109 28033 22143 28067
rect 26249 28033 26283 28067
rect 27169 28033 27203 28067
rect 27813 28033 27847 28067
rect 7389 27965 7423 27999
rect 10701 27965 10735 27999
rect 12725 27965 12759 27999
rect 13369 27965 13403 27999
rect 13553 27965 13587 27999
rect 14473 27965 14507 27999
rect 15669 27965 15703 27999
rect 17785 27965 17819 27999
rect 23213 27965 23247 27999
rect 23765 27965 23799 27999
rect 24777 27965 24811 27999
rect 26341 27965 26375 27999
rect 28549 27965 28583 27999
rect 29009 27965 29043 27999
rect 30757 27965 30791 27999
rect 11161 27829 11195 27863
rect 12173 27829 12207 27863
rect 14013 27829 14047 27863
rect 14841 27829 14875 27863
rect 16957 27829 16991 27863
rect 19349 27829 19383 27863
rect 20269 27829 20303 27863
rect 22201 27829 22235 27863
rect 27261 27829 27295 27863
rect 27905 27829 27939 27863
rect 9965 27625 9999 27659
rect 17601 27625 17635 27659
rect 12357 27557 12391 27591
rect 30481 27557 30515 27591
rect 7481 27489 7515 27523
rect 10793 27489 10827 27523
rect 11069 27489 11103 27523
rect 13277 27489 13311 27523
rect 14381 27489 14415 27523
rect 16313 27489 16347 27523
rect 19533 27489 19567 27523
rect 23029 27489 23063 27523
rect 24685 27489 24719 27523
rect 26249 27489 26283 27523
rect 26709 27489 26743 27523
rect 27813 27489 27847 27523
rect 28181 27489 28215 27523
rect 1593 27421 1627 27455
rect 9597 27421 9631 27455
rect 9781 27421 9815 27455
rect 12265 27421 12299 27455
rect 17509 27421 17543 27455
rect 19441 27421 19475 27455
rect 22937 27421 22971 27455
rect 23581 27421 23615 27455
rect 29745 27421 29779 27455
rect 30389 27421 30423 27455
rect 38301 27421 38335 27455
rect 7573 27353 7607 27387
rect 8493 27353 8527 27387
rect 10885 27353 10919 27387
rect 13001 27353 13035 27387
rect 13093 27353 13127 27387
rect 14473 27353 14507 27387
rect 15393 27353 15427 27387
rect 15945 27353 15979 27387
rect 16037 27353 16071 27387
rect 18245 27353 18279 27387
rect 18337 27353 18371 27387
rect 18889 27353 18923 27387
rect 20177 27353 20211 27387
rect 20269 27353 20303 27387
rect 20821 27353 20855 27387
rect 21833 27353 21867 27387
rect 21925 27353 21959 27387
rect 22477 27353 22511 27387
rect 23673 27353 23707 27387
rect 24777 27353 24811 27387
rect 25697 27353 25731 27387
rect 26341 27353 26375 27387
rect 27905 27353 27939 27387
rect 1777 27285 1811 27319
rect 29837 27285 29871 27319
rect 38117 27285 38151 27319
rect 1593 27081 1627 27115
rect 9781 27081 9815 27115
rect 10425 27081 10459 27115
rect 11069 27081 11103 27115
rect 33333 27081 33367 27115
rect 13001 27013 13035 27047
rect 13921 27013 13955 27047
rect 14565 27013 14599 27047
rect 17141 27013 17175 27047
rect 17233 27013 17267 27047
rect 18797 27013 18831 27047
rect 20545 27013 20579 27047
rect 22845 27013 22879 27047
rect 24685 27013 24719 27047
rect 27261 27013 27295 27047
rect 28181 27013 28215 27047
rect 29653 27013 29687 27047
rect 1777 26945 1811 26979
rect 9689 26945 9723 26979
rect 10333 26945 10367 26979
rect 10977 26945 11011 26979
rect 11897 26945 11931 26979
rect 15945 26945 15979 26979
rect 22017 26945 22051 26979
rect 26065 26945 26099 26979
rect 29561 26945 29595 26979
rect 32689 26945 32723 26979
rect 33241 26945 33275 26979
rect 38301 26945 38335 26979
rect 11713 26877 11747 26911
rect 12909 26877 12943 26911
rect 14473 26877 14507 26911
rect 15485 26877 15519 26911
rect 17417 26877 17451 26911
rect 18705 26877 18739 26911
rect 20453 26877 20487 26911
rect 20913 26877 20947 26911
rect 22753 26877 22787 26911
rect 23029 26877 23063 26911
rect 24593 26877 24627 26911
rect 24869 26877 24903 26911
rect 28089 26877 28123 26911
rect 28365 26877 28399 26911
rect 12081 26809 12115 26843
rect 19257 26809 19291 26843
rect 32505 26809 32539 26843
rect 16037 26741 16071 26775
rect 22109 26741 22143 26775
rect 26157 26741 26191 26775
rect 27353 26741 27387 26775
rect 38117 26741 38151 26775
rect 10149 26537 10183 26571
rect 10793 26537 10827 26571
rect 12081 26537 12115 26571
rect 14933 26537 14967 26571
rect 18797 26537 18831 26571
rect 27813 26537 27847 26571
rect 32689 26537 32723 26571
rect 11437 26469 11471 26503
rect 16497 26469 16531 26503
rect 25237 26469 25271 26503
rect 32045 26469 32079 26503
rect 12725 26401 12759 26435
rect 13001 26401 13035 26435
rect 14473 26401 14507 26435
rect 15945 26401 15979 26435
rect 17233 26401 17267 26435
rect 19809 26401 19843 26435
rect 21281 26401 21315 26435
rect 22845 26401 22879 26435
rect 26249 26401 26283 26435
rect 26525 26401 26559 26435
rect 28457 26401 28491 26435
rect 30481 26401 30515 26435
rect 10057 26333 10091 26367
rect 10701 26333 10735 26367
rect 11345 26333 11379 26367
rect 11989 26333 12023 26367
rect 14289 26333 14323 26367
rect 18705 26333 18739 26367
rect 27721 26333 27755 26367
rect 28365 26333 28399 26367
rect 29009 26333 29043 26367
rect 31309 26333 31343 26367
rect 31953 26333 31987 26367
rect 32597 26333 32631 26367
rect 12817 26265 12851 26299
rect 16030 26265 16064 26299
rect 17325 26265 17359 26299
rect 18245 26265 18279 26299
rect 19533 26265 19567 26299
rect 19625 26265 19659 26299
rect 21373 26265 21407 26299
rect 22293 26265 22327 26299
rect 22937 26265 22971 26299
rect 23857 26265 23891 26299
rect 24685 26265 24719 26299
rect 24777 26265 24811 26299
rect 26341 26265 26375 26299
rect 29101 26265 29135 26299
rect 29837 26265 29871 26299
rect 29929 26265 29963 26299
rect 31401 26197 31435 26231
rect 16957 25993 16991 26027
rect 17601 25993 17635 26027
rect 27813 25993 27847 26027
rect 30757 25993 30791 26027
rect 31401 25993 31435 26027
rect 11989 25925 12023 25959
rect 12541 25925 12575 25959
rect 15117 25925 15151 25959
rect 18889 25925 18923 25959
rect 23121 25925 23155 25959
rect 24593 25925 24627 25959
rect 24685 25925 24719 25959
rect 26433 25925 26467 25959
rect 29285 25925 29319 25959
rect 29377 25925 29411 25959
rect 9873 25857 9907 25891
rect 9965 25857 9999 25891
rect 10701 25857 10735 25891
rect 13093 25857 13127 25891
rect 13921 25857 13955 25891
rect 16865 25857 16899 25891
rect 17509 25857 17543 25891
rect 21281 25857 21315 25891
rect 22109 25857 22143 25891
rect 25697 25857 25731 25891
rect 26341 25857 26375 25891
rect 27169 25857 27203 25891
rect 27997 25857 28031 25891
rect 28549 25857 28583 25891
rect 31585 25857 31619 25891
rect 34161 25857 34195 25891
rect 10517 25789 10551 25823
rect 11161 25789 11195 25823
rect 11897 25789 11931 25823
rect 13737 25789 13771 25823
rect 15025 25789 15059 25823
rect 15669 25789 15703 25823
rect 18797 25789 18831 25823
rect 19809 25789 19843 25823
rect 23029 25789 23063 25823
rect 24041 25789 24075 25823
rect 24961 25789 24995 25823
rect 30297 25789 30331 25823
rect 13185 25721 13219 25755
rect 21373 25721 21407 25755
rect 27261 25721 27295 25755
rect 14105 25653 14139 25687
rect 22201 25653 22235 25687
rect 25789 25653 25823 25687
rect 28641 25653 28675 25687
rect 34253 25653 34287 25687
rect 10885 25449 10919 25483
rect 13737 25449 13771 25483
rect 9597 25313 9631 25347
rect 11621 25313 11655 25347
rect 12081 25313 12115 25347
rect 24869 25313 24903 25347
rect 25421 25313 25455 25347
rect 26985 25313 27019 25347
rect 27629 25313 27663 25347
rect 31769 25313 31803 25347
rect 33701 25313 33735 25347
rect 1593 25245 1627 25279
rect 9505 25245 9539 25279
rect 10149 25245 10183 25279
rect 10793 25245 10827 25279
rect 11437 25245 11471 25279
rect 13093 25245 13127 25279
rect 13277 25245 13311 25279
rect 16129 25245 16163 25279
rect 18429 25245 18463 25279
rect 19993 25245 20027 25279
rect 20637 25245 20671 25279
rect 38025 25245 38059 25279
rect 14381 25177 14415 25211
rect 14473 25177 14507 25211
rect 15393 25177 15427 25211
rect 16865 25177 16899 25211
rect 16957 25177 16991 25211
rect 17877 25177 17911 25211
rect 20085 25177 20119 25211
rect 21373 25177 21407 25211
rect 21465 25177 21499 25211
rect 22017 25177 22051 25211
rect 22753 25177 22787 25211
rect 22845 25177 22879 25211
rect 23765 25177 23799 25211
rect 24685 25177 24719 25211
rect 25513 25177 25547 25211
rect 26433 25177 26467 25211
rect 27077 25177 27111 25211
rect 29837 25177 29871 25211
rect 29929 25177 29963 25211
rect 30849 25177 30883 25211
rect 31493 25177 31527 25211
rect 31585 25177 31619 25211
rect 33793 25177 33827 25211
rect 34345 25177 34379 25211
rect 1777 25109 1811 25143
rect 10241 25109 10275 25143
rect 16221 25109 16255 25143
rect 18521 25109 18555 25143
rect 20729 25109 20763 25143
rect 38209 25109 38243 25143
rect 9505 24837 9539 24871
rect 12173 24837 12207 24871
rect 17049 24837 17083 24871
rect 19993 24837 20027 24871
rect 20913 24837 20947 24871
rect 22661 24837 22695 24871
rect 24225 24837 24259 24871
rect 27353 24837 27387 24871
rect 30297 24837 30331 24871
rect 1777 24769 1811 24803
rect 10977 24769 11011 24803
rect 12081 24769 12115 24803
rect 12725 24769 12759 24803
rect 13369 24769 13403 24803
rect 14565 24769 14599 24803
rect 15209 24769 15243 24803
rect 16129 24769 16163 24803
rect 18429 24769 18463 24803
rect 19165 24769 19199 24803
rect 19257 24769 19291 24803
rect 25605 24769 25639 24803
rect 26249 24769 26283 24803
rect 26341 24769 26375 24803
rect 32965 24769 32999 24803
rect 33057 24769 33091 24803
rect 38025 24769 38059 24803
rect 9413 24701 9447 24735
rect 9689 24701 9723 24735
rect 11069 24701 11103 24735
rect 16957 24701 16991 24735
rect 17325 24701 17359 24735
rect 18521 24701 18555 24735
rect 19901 24701 19935 24735
rect 22569 24701 22603 24735
rect 22845 24701 22879 24735
rect 24133 24701 24167 24735
rect 25145 24701 25179 24735
rect 27169 24701 27203 24735
rect 29009 24701 29043 24735
rect 29469 24701 29503 24735
rect 30205 24701 30239 24735
rect 30849 24701 30883 24735
rect 12817 24633 12851 24667
rect 1593 24565 1627 24599
rect 13461 24565 13495 24599
rect 14657 24565 14691 24599
rect 15301 24565 15335 24599
rect 16221 24565 16255 24599
rect 25697 24565 25731 24599
rect 38209 24565 38243 24599
rect 24685 24361 24719 24395
rect 25973 24361 26007 24395
rect 26617 24293 26651 24327
rect 9413 24225 9447 24259
rect 10149 24225 10183 24259
rect 11161 24225 11195 24259
rect 12541 24225 12575 24259
rect 15945 24225 15979 24259
rect 17601 24225 17635 24259
rect 17969 24225 18003 24259
rect 21097 24225 21131 24259
rect 21373 24225 21407 24259
rect 28457 24225 28491 24259
rect 30021 24225 30055 24259
rect 31033 24225 31067 24259
rect 32137 24225 32171 24259
rect 32413 24225 32447 24259
rect 1777 24157 1811 24191
rect 8309 24157 8343 24191
rect 13553 24157 13587 24191
rect 14289 24167 14323 24201
rect 15209 24167 15243 24201
rect 19809 24157 19843 24191
rect 24593 24157 24627 24191
rect 25237 24157 25271 24191
rect 25881 24157 25915 24191
rect 26525 24157 26559 24191
rect 27445 24157 27479 24191
rect 38301 24157 38335 24191
rect 10241 24089 10275 24123
rect 11989 24089 12023 24123
rect 12081 24089 12115 24123
rect 13645 24089 13679 24123
rect 16037 24089 16071 24123
rect 16957 24089 16991 24123
rect 17693 24089 17727 24123
rect 21189 24089 21223 24123
rect 23029 24089 23063 24123
rect 23121 24089 23155 24123
rect 24041 24089 24075 24123
rect 28170 24089 28204 24123
rect 28266 24089 28300 24123
rect 30113 24089 30147 24123
rect 32229 24089 32263 24123
rect 1593 24021 1627 24055
rect 8401 24021 8435 24055
rect 14381 24021 14415 24055
rect 15301 24021 15335 24055
rect 19901 24021 19935 24055
rect 25329 24021 25363 24055
rect 27537 24021 27571 24055
rect 38117 24021 38151 24055
rect 1777 23817 1811 23851
rect 2421 23817 2455 23851
rect 10333 23817 10367 23851
rect 18245 23817 18279 23851
rect 30389 23817 30423 23851
rect 31677 23817 31711 23851
rect 33701 23817 33735 23851
rect 37841 23817 37875 23851
rect 11069 23749 11103 23783
rect 13829 23749 13863 23783
rect 15393 23749 15427 23783
rect 16313 23749 16347 23783
rect 18889 23749 18923 23783
rect 18981 23749 19015 23783
rect 20354 23749 20388 23783
rect 22098 23749 22132 23783
rect 22210 23749 22244 23783
rect 24317 23749 24351 23783
rect 26525 23749 26559 23783
rect 27353 23749 27387 23783
rect 28917 23749 28951 23783
rect 32597 23749 32631 23783
rect 1961 23681 1995 23715
rect 2605 23681 2639 23715
rect 10517 23681 10551 23715
rect 10977 23681 11011 23715
rect 11805 23681 11839 23715
rect 12541 23681 12575 23715
rect 16865 23681 16899 23715
rect 17509 23681 17543 23715
rect 18153 23681 18187 23715
rect 23581 23681 23615 23715
rect 24225 23681 24259 23715
rect 24869 23681 24903 23715
rect 25513 23681 25547 23715
rect 26433 23681 26467 23715
rect 30297 23681 30331 23715
rect 30941 23681 30975 23715
rect 31585 23681 31619 23715
rect 32505 23681 32539 23715
rect 33885 23681 33919 23715
rect 38025 23681 38059 23715
rect 13737 23613 13771 23647
rect 14565 23613 14599 23647
rect 15301 23613 15335 23647
rect 20269 23613 20303 23647
rect 20729 23613 20763 23647
rect 22385 23613 22419 23647
rect 27261 23613 27295 23647
rect 27537 23613 27571 23647
rect 28825 23613 28859 23647
rect 29101 23613 29135 23647
rect 12725 23545 12759 23579
rect 19441 23545 19475 23579
rect 11897 23477 11931 23511
rect 16957 23477 16991 23511
rect 17601 23477 17635 23511
rect 23673 23477 23707 23511
rect 24961 23477 24995 23511
rect 25605 23477 25639 23511
rect 31033 23477 31067 23511
rect 9137 23273 9171 23307
rect 10701 23273 10735 23307
rect 13645 23273 13679 23307
rect 23949 23273 23983 23307
rect 27813 23273 27847 23307
rect 28457 23273 28491 23307
rect 7297 23137 7331 23171
rect 14381 23137 14415 23171
rect 14657 23137 14691 23171
rect 15853 23137 15887 23171
rect 18429 23137 18463 23171
rect 22937 23137 22971 23171
rect 24685 23137 24719 23171
rect 29837 23137 29871 23171
rect 7205 23069 7239 23103
rect 7849 23069 7883 23103
rect 9321 23069 9355 23103
rect 10609 23069 10643 23103
rect 11253 23069 11287 23103
rect 13553 23069 13587 23103
rect 19441 23069 19475 23103
rect 21005 23069 21039 23103
rect 21649 23069 21683 23103
rect 21741 23069 21775 23103
rect 23857 23069 23891 23103
rect 26157 23069 26191 23103
rect 27077 23069 27111 23103
rect 27721 23069 27755 23103
rect 28365 23069 28399 23103
rect 29009 23069 29043 23103
rect 31309 23069 31343 23103
rect 35265 23069 35299 23103
rect 11989 23001 12023 23035
rect 12081 23001 12115 23035
rect 13001 23001 13035 23035
rect 14473 23001 14507 23035
rect 15945 23001 15979 23035
rect 16865 23001 16899 23035
rect 17417 23001 17451 23035
rect 17509 23001 17543 23035
rect 19533 23001 19567 23035
rect 22385 23001 22419 23035
rect 22477 23001 22511 23035
rect 24777 23001 24811 23035
rect 25697 23001 25731 23035
rect 29929 23001 29963 23035
rect 30849 23001 30883 23035
rect 32045 23001 32079 23035
rect 32137 23001 32171 23035
rect 33057 23001 33091 23035
rect 7941 22933 7975 22967
rect 11345 22933 11379 22967
rect 21097 22933 21131 22967
rect 26249 22933 26283 22967
rect 27169 22933 27203 22967
rect 29101 22933 29135 22967
rect 31401 22933 31435 22967
rect 35081 22933 35115 22967
rect 19625 22729 19659 22763
rect 20269 22729 20303 22763
rect 7757 22661 7791 22695
rect 10241 22661 10275 22695
rect 11161 22661 11195 22695
rect 13369 22661 13403 22695
rect 15117 22661 15151 22695
rect 15209 22661 15243 22695
rect 22477 22661 22511 22695
rect 24225 22661 24259 22695
rect 27353 22661 27387 22695
rect 28549 22661 28583 22695
rect 29469 22661 29503 22695
rect 30205 22661 30239 22695
rect 31125 22661 31159 22695
rect 1777 22593 1811 22627
rect 12081 22593 12115 22627
rect 12541 22593 12575 22627
rect 17233 22593 17267 22627
rect 18337 22593 18371 22627
rect 19533 22593 19567 22627
rect 20177 22593 20211 22627
rect 25605 22593 25639 22627
rect 26249 22593 26283 22627
rect 31585 22593 31619 22627
rect 32321 22593 32355 22627
rect 32965 22593 32999 22627
rect 34897 22593 34931 22627
rect 38025 22593 38059 22627
rect 7573 22525 7607 22559
rect 9413 22525 9447 22559
rect 10149 22525 10183 22559
rect 13277 22525 13311 22559
rect 14289 22525 14323 22559
rect 16129 22525 16163 22559
rect 22385 22525 22419 22559
rect 22661 22525 22695 22559
rect 24133 22525 24167 22559
rect 25145 22525 25179 22559
rect 27261 22525 27295 22559
rect 27537 22525 27571 22559
rect 28457 22525 28491 22559
rect 30113 22525 30147 22559
rect 33057 22457 33091 22491
rect 38209 22457 38243 22491
rect 1593 22389 1627 22423
rect 11897 22389 11931 22423
rect 12633 22389 12667 22423
rect 17325 22389 17359 22423
rect 18429 22389 18463 22423
rect 25697 22389 25731 22423
rect 26341 22389 26375 22423
rect 31677 22389 31711 22423
rect 32413 22389 32447 22423
rect 34989 22389 35023 22423
rect 8401 22185 8435 22219
rect 38117 22117 38151 22151
rect 7481 22049 7515 22083
rect 10149 22049 10183 22083
rect 12725 22049 12759 22083
rect 15117 22049 15151 22083
rect 15761 22049 15795 22083
rect 18797 22049 18831 22083
rect 20453 22049 20487 22083
rect 23581 22049 23615 22083
rect 25973 22049 26007 22083
rect 27905 22049 27939 22083
rect 30849 22049 30883 22083
rect 33793 22049 33827 22083
rect 1593 21981 1627 22015
rect 7389 21981 7423 22015
rect 8309 21981 8343 22015
rect 13553 21981 13587 22015
rect 14381 21981 14415 22015
rect 19717 21981 19751 22015
rect 22661 21981 22695 22015
rect 23489 21981 23523 22015
rect 32321 21981 32355 22015
rect 33057 21981 33091 22015
rect 33701 21981 33735 22015
rect 35173 21981 35207 22015
rect 38301 21981 38335 22015
rect 10241 21913 10275 21947
rect 11161 21913 11195 21947
rect 11713 21913 11747 21947
rect 11805 21913 11839 21947
rect 15209 21913 15243 21947
rect 16313 21913 16347 21947
rect 16405 21913 16439 21947
rect 16957 21913 16991 21947
rect 17785 21913 17819 21947
rect 17877 21913 17911 21947
rect 19809 21913 19843 21947
rect 20545 21913 20579 21947
rect 21097 21913 21131 21947
rect 25145 21913 25179 21947
rect 25237 21913 25271 21947
rect 26893 21913 26927 21947
rect 26985 21913 27019 21947
rect 28457 21913 28491 21947
rect 28549 21913 28583 21947
rect 29101 21913 29135 21947
rect 30941 21913 30975 21947
rect 31861 21913 31895 21947
rect 33149 21913 33183 21947
rect 1777 21845 1811 21879
rect 13645 21845 13679 21879
rect 14473 21845 14507 21879
rect 22753 21845 22787 21879
rect 29745 21845 29779 21879
rect 32413 21845 32447 21879
rect 34989 21845 35023 21879
rect 10425 21641 10459 21675
rect 11069 21641 11103 21675
rect 12449 21641 12483 21675
rect 15301 21641 15335 21675
rect 20361 21641 20395 21675
rect 22109 21641 22143 21675
rect 27813 21641 27847 21675
rect 33057 21641 33091 21675
rect 13093 21573 13127 21607
rect 13829 21573 13863 21607
rect 14381 21573 14415 21607
rect 16037 21573 16071 21607
rect 17233 21573 17267 21607
rect 19073 21573 19107 21607
rect 23673 21573 23707 21607
rect 25237 21573 25271 21607
rect 28542 21573 28576 21607
rect 29653 21573 29687 21607
rect 30757 21573 30791 21607
rect 30849 21573 30883 21607
rect 10333 21505 10367 21539
rect 10977 21505 11011 21539
rect 11713 21505 11747 21539
rect 12357 21505 12391 21539
rect 13001 21505 13035 21539
rect 15945 21505 15979 21539
rect 18337 21505 18371 21539
rect 18981 21505 19015 21539
rect 19625 21505 19659 21539
rect 20269 21505 20303 21539
rect 20913 21505 20947 21539
rect 22017 21505 22051 21539
rect 22661 21505 22695 21539
rect 27629 21505 27663 21539
rect 29561 21505 29595 21539
rect 32321 21505 32355 21539
rect 32965 21505 32999 21539
rect 33609 21505 33643 21539
rect 34253 21505 34287 21539
rect 13737 21437 13771 21471
rect 17141 21437 17175 21471
rect 23581 21437 23615 21471
rect 24133 21437 24167 21471
rect 25145 21437 25179 21471
rect 25973 21437 26007 21471
rect 28458 21437 28492 21471
rect 31033 21437 31067 21471
rect 33701 21437 33735 21471
rect 17693 21369 17727 21403
rect 29009 21369 29043 21403
rect 11805 21301 11839 21335
rect 18429 21301 18463 21335
rect 19717 21301 19751 21335
rect 21005 21301 21039 21335
rect 22753 21301 22787 21335
rect 32413 21301 32447 21335
rect 34345 21301 34379 21335
rect 13645 21097 13679 21131
rect 14565 21097 14599 21131
rect 23949 21097 23983 21131
rect 24685 21097 24719 21131
rect 38117 21097 38151 21131
rect 29837 21029 29871 21063
rect 31033 21029 31067 21063
rect 15853 20961 15887 20995
rect 17417 20961 17451 20995
rect 25513 20961 25547 20995
rect 25697 20961 25731 20995
rect 27997 20961 28031 20995
rect 28273 20961 28307 20995
rect 30481 20961 30515 20995
rect 31861 20961 31895 20995
rect 1593 20893 1627 20927
rect 12081 20893 12115 20927
rect 13553 20893 13587 20927
rect 14473 20893 14507 20927
rect 15117 20893 15151 20927
rect 21465 20893 21499 20927
rect 23857 20893 23891 20927
rect 24593 20893 24627 20927
rect 29745 20893 29779 20927
rect 32965 20893 32999 20927
rect 33609 20893 33643 20927
rect 38301 20893 38335 20927
rect 15945 20825 15979 20859
rect 16865 20825 16899 20859
rect 17509 20825 17543 20859
rect 18429 20825 18463 20859
rect 19901 20825 19935 20859
rect 19993 20825 20027 20859
rect 20913 20825 20947 20859
rect 22201 20825 22235 20859
rect 22293 20825 22327 20859
rect 23213 20825 23247 20859
rect 27353 20825 27387 20859
rect 28089 20825 28123 20859
rect 30573 20825 30607 20859
rect 31953 20825 31987 20859
rect 32505 20825 32539 20859
rect 33701 20825 33735 20859
rect 1777 20757 1811 20791
rect 12173 20757 12207 20791
rect 15209 20757 15243 20791
rect 21557 20757 21591 20791
rect 33057 20757 33091 20791
rect 6837 20553 6871 20587
rect 13737 20553 13771 20587
rect 16221 20553 16255 20587
rect 20361 20553 20395 20587
rect 14473 20485 14507 20519
rect 17049 20485 17083 20519
rect 18889 20485 18923 20519
rect 22201 20485 22235 20519
rect 24041 20485 24075 20519
rect 24133 20485 24167 20519
rect 27353 20485 27387 20519
rect 28917 20485 28951 20519
rect 30757 20485 30791 20519
rect 32413 20485 32447 20519
rect 32505 20485 32539 20519
rect 33609 20485 33643 20519
rect 1961 20417 1995 20451
rect 7021 20417 7055 20451
rect 12173 20417 12207 20451
rect 13001 20417 13035 20451
rect 13645 20417 13679 20451
rect 16129 20417 16163 20451
rect 20269 20417 20303 20451
rect 20913 20417 20947 20451
rect 25513 20417 25547 20451
rect 26157 20417 26191 20451
rect 33517 20417 33551 20451
rect 34161 20417 34195 20451
rect 34805 20417 34839 20451
rect 14381 20349 14415 20383
rect 15209 20349 15243 20383
rect 16957 20349 16991 20383
rect 17877 20349 17911 20383
rect 18797 20349 18831 20383
rect 19809 20349 19843 20383
rect 22109 20349 22143 20383
rect 23121 20349 23155 20383
rect 24317 20349 24351 20383
rect 27261 20349 27295 20383
rect 27629 20349 27663 20383
rect 28825 20349 28859 20383
rect 29101 20349 29135 20383
rect 30665 20349 30699 20383
rect 31309 20349 31343 20383
rect 34253 20349 34287 20383
rect 13093 20281 13127 20315
rect 32965 20281 32999 20315
rect 1777 20213 1811 20247
rect 12265 20213 12299 20247
rect 21005 20213 21039 20247
rect 25605 20213 25639 20247
rect 26249 20213 26283 20247
rect 34897 20213 34931 20247
rect 16129 20009 16163 20043
rect 17417 20009 17451 20043
rect 33057 20009 33091 20043
rect 34989 20009 35023 20043
rect 20085 19941 20119 19975
rect 38301 19941 38335 19975
rect 1869 19873 1903 19907
rect 12265 19873 12299 19907
rect 19533 19873 19567 19907
rect 21373 19873 21407 19907
rect 22937 19873 22971 19907
rect 23213 19873 23247 19907
rect 24685 19873 24719 19907
rect 24961 19873 24995 19907
rect 26985 19873 27019 19907
rect 27445 19873 27479 19907
rect 28733 19873 28767 19907
rect 29837 19873 29871 19907
rect 33701 19873 33735 19907
rect 1593 19805 1627 19839
rect 12909 19805 12943 19839
rect 15393 19805 15427 19839
rect 16037 19805 16071 19839
rect 16681 19805 16715 19839
rect 17325 19805 17359 19839
rect 20637 19805 20671 19839
rect 26157 19805 26191 19839
rect 28089 19805 28123 19839
rect 30481 19805 30515 19839
rect 31861 19805 31895 19839
rect 32321 19805 32355 19839
rect 32965 19805 32999 19839
rect 33609 19805 33643 19839
rect 34897 19805 34931 19839
rect 11621 19737 11655 19771
rect 11713 19737 11747 19771
rect 15485 19737 15519 19771
rect 18061 19737 18095 19771
rect 18153 19737 18187 19771
rect 18705 19737 18739 19771
rect 19625 19737 19659 19771
rect 21465 19737 21499 19771
rect 22385 19737 22419 19771
rect 23029 19737 23063 19771
rect 24754 19737 24788 19771
rect 27077 19737 27111 19771
rect 29929 19737 29963 19771
rect 31217 19737 31251 19771
rect 31309 19737 31343 19771
rect 38117 19737 38151 19771
rect 13001 19669 13035 19703
rect 16773 19669 16807 19703
rect 20729 19669 20763 19703
rect 26249 19669 26283 19703
rect 28181 19669 28215 19703
rect 32413 19669 32447 19703
rect 7573 19465 7607 19499
rect 8401 19465 8435 19499
rect 9137 19465 9171 19499
rect 13185 19465 13219 19499
rect 13829 19465 13863 19499
rect 14473 19465 14507 19499
rect 28825 19465 28859 19499
rect 35173 19465 35207 19499
rect 36277 19465 36311 19499
rect 38117 19465 38151 19499
rect 10149 19397 10183 19431
rect 10241 19397 10275 19431
rect 17417 19397 17451 19431
rect 18613 19397 18647 19431
rect 20177 19397 20211 19431
rect 21097 19397 21131 19431
rect 22109 19397 22143 19431
rect 22937 19397 22971 19431
rect 23666 19397 23700 19431
rect 25145 19397 25179 19431
rect 25237 19397 25271 19431
rect 27353 19397 27387 19431
rect 29745 19397 29779 19431
rect 31217 19397 31251 19431
rect 33425 19397 33459 19431
rect 33517 19397 33551 19431
rect 34621 19397 34655 19431
rect 1593 19329 1627 19363
rect 7481 19329 7515 19363
rect 8585 19329 8619 19363
rect 9045 19329 9079 19363
rect 13093 19329 13127 19363
rect 13737 19329 13771 19363
rect 14381 19329 14415 19363
rect 15117 19329 15151 19363
rect 15209 19329 15243 19363
rect 22017 19329 22051 19363
rect 22845 19329 22879 19363
rect 28733 19329 28767 19363
rect 32321 19329 32355 19363
rect 34529 19329 34563 19363
rect 36461 19329 36495 19363
rect 38301 19329 38335 19363
rect 11161 19261 11195 19295
rect 17325 19261 17359 19295
rect 18521 19261 18555 19295
rect 19533 19261 19567 19295
rect 20085 19261 20119 19295
rect 23581 19261 23615 19295
rect 24133 19261 24167 19295
rect 26157 19261 26191 19295
rect 27261 19261 27295 19295
rect 28273 19261 28307 19295
rect 29653 19261 29687 19295
rect 30021 19261 30055 19295
rect 33701 19261 33735 19295
rect 17877 19193 17911 19227
rect 31401 19193 31435 19227
rect 1777 19125 1811 19159
rect 32413 19125 32447 19159
rect 8401 18921 8435 18955
rect 12633 18921 12667 18955
rect 17049 18921 17083 18955
rect 18613 18921 18647 18955
rect 24685 18921 24719 18955
rect 34989 18921 35023 18955
rect 23489 18853 23523 18887
rect 11069 18785 11103 18819
rect 12081 18785 12115 18819
rect 19533 18785 19567 18819
rect 22937 18785 22971 18819
rect 29837 18785 29871 18819
rect 30481 18785 30515 18819
rect 32781 18785 32815 18819
rect 33149 18785 33183 18819
rect 6561 18717 6595 18751
rect 8309 18717 8343 18751
rect 12541 18717 12575 18751
rect 13185 18717 13219 18751
rect 15945 18717 15979 18751
rect 16957 18717 16991 18751
rect 18521 18717 18555 18751
rect 20637 18717 20671 18751
rect 21557 18717 21591 18751
rect 22201 18717 22235 18751
rect 24593 18717 24627 18751
rect 28825 18717 28859 18751
rect 34897 18717 34931 18751
rect 11161 18649 11195 18683
rect 19625 18649 19659 18683
rect 20177 18649 20211 18683
rect 23029 18649 23063 18683
rect 25789 18649 25823 18683
rect 25881 18649 25915 18683
rect 26801 18649 26835 18683
rect 27353 18649 27387 18683
rect 27445 18649 27479 18683
rect 28365 18649 28399 18683
rect 29929 18649 29963 18683
rect 31033 18649 31067 18683
rect 31125 18649 31159 18683
rect 31677 18649 31711 18683
rect 32873 18649 32907 18683
rect 6653 18581 6687 18615
rect 13277 18581 13311 18615
rect 16037 18581 16071 18615
rect 20729 18581 20763 18615
rect 21649 18581 21683 18615
rect 22293 18581 22327 18615
rect 28917 18581 28951 18615
rect 1593 18377 1627 18411
rect 13277 18377 13311 18411
rect 15669 18377 15703 18411
rect 33609 18377 33643 18411
rect 34897 18377 34931 18411
rect 6745 18309 6779 18343
rect 12173 18309 12207 18343
rect 12725 18309 12759 18343
rect 18061 18309 18095 18343
rect 20269 18309 20303 18343
rect 20361 18309 20395 18343
rect 23857 18309 23891 18343
rect 23949 18309 23983 18343
rect 26065 18309 26099 18343
rect 27353 18309 27387 18343
rect 28733 18309 28767 18343
rect 31033 18309 31067 18343
rect 32413 18309 32447 18343
rect 32505 18309 32539 18343
rect 34253 18309 34287 18343
rect 1777 18241 1811 18275
rect 9045 18241 9079 18275
rect 13185 18241 13219 18275
rect 15577 18241 15611 18275
rect 17233 18241 17267 18275
rect 19441 18241 19475 18275
rect 22293 18241 22327 18275
rect 22937 18241 22971 18275
rect 27905 18241 27939 18275
rect 28549 18241 28583 18275
rect 33517 18241 33551 18275
rect 34161 18241 34195 18275
rect 34805 18241 34839 18275
rect 35633 18241 35667 18275
rect 38117 18241 38151 18275
rect 6653 18173 6687 18207
rect 7665 18173 7699 18207
rect 8125 18173 8159 18207
rect 12081 18173 12115 18207
rect 17969 18173 18003 18207
rect 18337 18173 18371 18207
rect 24777 18173 24811 18207
rect 25973 18173 26007 18207
rect 27261 18173 27295 18207
rect 30205 18173 30239 18207
rect 30941 18173 30975 18207
rect 32689 18173 32723 18207
rect 20821 18105 20855 18139
rect 26525 18105 26559 18139
rect 31493 18105 31527 18139
rect 38301 18105 38335 18139
rect 9137 18037 9171 18071
rect 17325 18037 17359 18071
rect 19533 18037 19567 18071
rect 22385 18037 22419 18071
rect 23029 18037 23063 18071
rect 35449 18037 35483 18071
rect 6561 17833 6595 17867
rect 21097 17833 21131 17867
rect 32781 17833 32815 17867
rect 27353 17765 27387 17799
rect 9229 17697 9263 17731
rect 13185 17697 13219 17731
rect 16497 17697 16531 17731
rect 17509 17697 17543 17731
rect 24685 17697 24719 17731
rect 26801 17697 26835 17731
rect 28641 17697 28675 17731
rect 6469 17629 6503 17663
rect 7113 17629 7147 17663
rect 7757 17629 7791 17663
rect 8401 17629 8435 17663
rect 10793 17629 10827 17663
rect 11437 17629 11471 17663
rect 14289 17629 14323 17663
rect 15117 17629 15151 17663
rect 15761 17629 15795 17663
rect 18061 17629 18095 17663
rect 18705 17629 18739 17663
rect 21005 17629 21039 17663
rect 23305 17629 23339 17663
rect 27905 17629 27939 17663
rect 28549 17629 28583 17663
rect 32689 17629 32723 17663
rect 33333 17629 33367 17663
rect 33977 17629 34011 17663
rect 34897 17629 34931 17663
rect 34989 17629 35023 17663
rect 35725 17629 35759 17663
rect 7849 17561 7883 17595
rect 9321 17561 9355 17595
rect 9873 17561 9907 17595
rect 12173 17561 12207 17595
rect 12265 17561 12299 17595
rect 16589 17561 16623 17595
rect 19717 17561 19751 17595
rect 19809 17561 19843 17595
rect 20361 17561 20395 17595
rect 21833 17561 21867 17595
rect 21925 17561 21959 17595
rect 22845 17561 22879 17595
rect 24777 17561 24811 17595
rect 25697 17561 25731 17595
rect 26893 17561 26927 17595
rect 30021 17561 30055 17595
rect 30113 17561 30147 17595
rect 31033 17561 31067 17595
rect 31585 17561 31619 17595
rect 31677 17561 31711 17595
rect 32229 17561 32263 17595
rect 33425 17561 33459 17595
rect 7205 17493 7239 17527
rect 8493 17493 8527 17527
rect 10885 17493 10919 17527
rect 11529 17493 11563 17527
rect 14381 17493 14415 17527
rect 15209 17493 15243 17527
rect 15853 17493 15887 17527
rect 18153 17493 18187 17527
rect 18797 17493 18831 17527
rect 23397 17493 23431 17527
rect 27997 17493 28031 17527
rect 34069 17493 34103 17527
rect 35541 17493 35575 17527
rect 16957 17289 16991 17323
rect 31677 17289 31711 17323
rect 32413 17289 32447 17323
rect 33057 17289 33091 17323
rect 33701 17289 33735 17323
rect 7021 17221 7055 17255
rect 7573 17221 7607 17255
rect 8125 17221 8159 17255
rect 8217 17221 8251 17255
rect 9137 17221 9171 17255
rect 11897 17221 11931 17255
rect 15301 17221 15335 17255
rect 18337 17221 18371 17255
rect 20913 17221 20947 17255
rect 22293 17221 22327 17255
rect 22385 17221 22419 17255
rect 23949 17221 23983 17255
rect 24869 17221 24903 17255
rect 25513 17221 25547 17255
rect 28641 17221 28675 17255
rect 30205 17221 30239 17255
rect 1869 17153 1903 17187
rect 5825 17153 5859 17187
rect 9689 17153 9723 17187
rect 10333 17153 10367 17187
rect 10977 17153 11011 17187
rect 13461 17153 13495 17187
rect 14473 17153 14507 17187
rect 16865 17153 16899 17187
rect 17509 17153 17543 17187
rect 19717 17153 19751 17187
rect 27169 17153 27203 17187
rect 31585 17153 31619 17187
rect 32321 17153 32355 17187
rect 32965 17153 32999 17187
rect 33609 17153 33643 17187
rect 38301 17153 38335 17187
rect 1593 17085 1627 17119
rect 5917 17085 5951 17119
rect 6929 17085 6963 17119
rect 11805 17085 11839 17119
rect 12449 17085 12483 17119
rect 15209 17085 15243 17119
rect 15669 17085 15703 17119
rect 18245 17085 18279 17119
rect 18521 17085 18555 17119
rect 19993 17085 20027 17119
rect 20821 17085 20855 17119
rect 23305 17085 23339 17119
rect 23857 17085 23891 17119
rect 25421 17085 25455 17119
rect 26433 17085 26467 17119
rect 27353 17085 27387 17119
rect 28549 17085 28583 17119
rect 29377 17085 29411 17119
rect 30113 17085 30147 17119
rect 31033 17085 31067 17119
rect 21373 17017 21407 17051
rect 9781 16949 9815 16983
rect 10425 16949 10459 16983
rect 11069 16949 11103 16983
rect 13553 16949 13587 16983
rect 14565 16949 14599 16983
rect 17601 16949 17635 16983
rect 38117 16949 38151 16983
rect 23305 16745 23339 16779
rect 25973 16745 26007 16779
rect 7389 16609 7423 16643
rect 8217 16609 8251 16643
rect 15945 16609 15979 16643
rect 20085 16609 20119 16643
rect 30941 16609 30975 16643
rect 32505 16609 32539 16643
rect 1961 16541 1995 16575
rect 5365 16541 5399 16575
rect 6009 16541 6043 16575
rect 6653 16541 6687 16575
rect 10977 16541 11011 16575
rect 11621 16541 11655 16575
rect 12265 16541 12299 16575
rect 12909 16541 12943 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 14933 16541 14967 16575
rect 17049 16541 17083 16575
rect 18061 16541 18095 16575
rect 18705 16541 18739 16575
rect 24593 16541 24627 16575
rect 25237 16541 25271 16575
rect 25329 16541 25363 16575
rect 25881 16541 25915 16575
rect 28457 16541 28491 16575
rect 29745 16541 29779 16575
rect 33977 16541 34011 16575
rect 34897 16541 34931 16575
rect 6745 16473 6779 16507
rect 7481 16473 7515 16507
rect 9229 16473 9263 16507
rect 9321 16473 9355 16507
rect 10241 16473 10275 16507
rect 15025 16473 15059 16507
rect 15669 16473 15703 16507
rect 15761 16473 15795 16507
rect 20177 16473 20211 16507
rect 21097 16473 21131 16507
rect 21649 16473 21683 16507
rect 21741 16473 21775 16507
rect 22661 16473 22695 16507
rect 23213 16473 23247 16507
rect 24685 16473 24719 16507
rect 26985 16473 27019 16507
rect 27077 16473 27111 16507
rect 27997 16473 28031 16507
rect 28733 16473 28767 16507
rect 29837 16473 29871 16507
rect 31033 16473 31067 16507
rect 31953 16473 31987 16507
rect 32597 16473 32631 16507
rect 33517 16473 33551 16507
rect 34989 16473 35023 16507
rect 1777 16405 1811 16439
rect 5457 16405 5491 16439
rect 6101 16405 6135 16439
rect 11069 16405 11103 16439
rect 11713 16405 11747 16439
rect 12357 16405 12391 16439
rect 13001 16405 13035 16439
rect 13645 16405 13679 16439
rect 14381 16405 14415 16439
rect 17141 16405 17175 16439
rect 18153 16405 18187 16439
rect 18797 16405 18831 16439
rect 34069 16405 34103 16439
rect 24133 16201 24167 16235
rect 31033 16201 31067 16235
rect 31677 16201 31711 16235
rect 6837 16133 6871 16167
rect 8401 16133 8435 16167
rect 10241 16133 10275 16167
rect 11805 16133 11839 16167
rect 11897 16133 11931 16167
rect 12817 16133 12851 16167
rect 14381 16133 14415 16167
rect 17141 16133 17175 16167
rect 17233 16133 17267 16167
rect 18889 16133 18923 16167
rect 22477 16133 22511 16167
rect 22569 16133 22603 16167
rect 24777 16133 24811 16167
rect 27353 16133 27387 16167
rect 32505 16133 32539 16167
rect 1593 16065 1627 16099
rect 13461 16065 13495 16099
rect 16129 16063 16163 16097
rect 20269 16065 20303 16099
rect 21281 16065 21315 16099
rect 24041 16065 24075 16099
rect 24685 16065 24719 16099
rect 25329 16065 25363 16099
rect 25973 16065 26007 16099
rect 28733 16065 28767 16099
rect 29653 16065 29687 16099
rect 30297 16065 30331 16099
rect 30941 16065 30975 16099
rect 31585 16065 31619 16099
rect 38025 16065 38059 16099
rect 5825 15997 5859 16031
rect 6745 15997 6779 16031
rect 7021 15997 7055 16031
rect 8309 15997 8343 16031
rect 8677 15997 8711 16031
rect 10149 15997 10183 16031
rect 11161 15997 11195 16031
rect 14289 15997 14323 16031
rect 14565 15997 14599 16031
rect 17969 15997 18003 16031
rect 18797 15997 18831 16031
rect 19073 15997 19107 16031
rect 23489 15997 23523 16031
rect 26249 15997 26283 16031
rect 27261 15997 27295 16031
rect 28273 15997 28307 16031
rect 29009 15997 29043 16031
rect 32413 15997 32447 16031
rect 33425 15997 33459 16031
rect 30389 15929 30423 15963
rect 1777 15861 1811 15895
rect 13553 15861 13587 15895
rect 16221 15861 16255 15895
rect 20361 15861 20395 15895
rect 21373 15861 21407 15895
rect 25421 15861 25455 15895
rect 29745 15861 29779 15895
rect 38209 15861 38243 15895
rect 26893 15657 26927 15691
rect 29837 15657 29871 15691
rect 30481 15657 30515 15691
rect 31769 15657 31803 15691
rect 7297 15521 7331 15555
rect 8217 15521 8251 15555
rect 9689 15521 9723 15555
rect 9965 15521 9999 15555
rect 13001 15521 13035 15555
rect 18797 15521 18831 15555
rect 21097 15521 21131 15555
rect 22937 15521 22971 15555
rect 24869 15521 24903 15555
rect 33333 15521 33367 15555
rect 5181 15453 5215 15487
rect 11621 15453 11655 15487
rect 12265 15453 12299 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 14841 15453 14875 15487
rect 15485 15453 15519 15487
rect 16129 15453 16163 15487
rect 16773 15453 16807 15487
rect 17417 15453 17451 15487
rect 18061 15453 18095 15487
rect 18697 15453 18731 15487
rect 19625 15453 19659 15487
rect 20269 15453 20303 15487
rect 20913 15453 20947 15487
rect 21833 15453 21867 15487
rect 22109 15453 22143 15487
rect 22753 15453 22787 15487
rect 23673 15453 23707 15487
rect 24593 15453 24627 15487
rect 25513 15453 25547 15487
rect 26157 15453 26191 15487
rect 26801 15453 26835 15487
rect 27537 15453 27571 15487
rect 28641 15453 28675 15487
rect 29745 15453 29779 15487
rect 30389 15453 30423 15487
rect 31033 15453 31067 15487
rect 31677 15453 31711 15487
rect 38025 15453 38059 15487
rect 1685 15385 1719 15419
rect 1869 15385 1903 15419
rect 5273 15385 5307 15419
rect 5917 15385 5951 15419
rect 6009 15385 6043 15419
rect 6561 15385 6595 15419
rect 7389 15385 7423 15419
rect 9781 15385 9815 15419
rect 17509 15385 17543 15419
rect 28089 15385 28123 15419
rect 33425 15385 33459 15419
rect 34345 15385 34379 15419
rect 11713 15317 11747 15351
rect 12357 15317 12391 15351
rect 13645 15317 13679 15351
rect 14933 15317 14967 15351
rect 15577 15317 15611 15351
rect 16221 15317 16255 15351
rect 16865 15317 16899 15351
rect 18153 15317 18187 15351
rect 19717 15317 19751 15351
rect 20361 15317 20395 15351
rect 23765 15317 23799 15351
rect 25605 15317 25639 15351
rect 26249 15317 26283 15351
rect 28733 15317 28767 15351
rect 31125 15317 31159 15351
rect 38209 15317 38243 15351
rect 32413 15113 32447 15147
rect 6929 15045 6963 15079
rect 8309 15045 8343 15079
rect 10149 15045 10183 15079
rect 16221 15045 16255 15079
rect 18705 15045 18739 15079
rect 29837 15045 29871 15079
rect 30665 15045 30699 15079
rect 31217 15045 31251 15079
rect 6009 14977 6043 15011
rect 14841 14977 14875 15011
rect 15485 14977 15519 15011
rect 16129 14977 16163 15011
rect 17233 14977 17267 15011
rect 17877 14977 17911 15011
rect 20361 14977 20395 15011
rect 21005 14977 21039 15011
rect 22293 14977 22327 15011
rect 23673 14977 23707 15011
rect 24593 14977 24627 15011
rect 25237 14977 25271 15011
rect 25881 14977 25915 15011
rect 27169 14977 27203 15011
rect 27813 14977 27847 15011
rect 28457 14977 28491 15011
rect 29101 14977 29135 15011
rect 29745 14977 29779 15011
rect 32321 14977 32355 15011
rect 38025 14977 38059 15011
rect 6837 14909 6871 14943
rect 7481 14909 7515 14943
rect 8217 14909 8251 14943
rect 8493 14909 8527 14943
rect 10057 14909 10091 14943
rect 10701 14909 10735 14943
rect 12265 14909 12299 14943
rect 14289 14909 14323 14943
rect 18613 14909 18647 14943
rect 18889 14909 18923 14943
rect 20453 14909 20487 14943
rect 21281 14909 21315 14943
rect 23029 14909 23063 14943
rect 23857 14909 23891 14943
rect 25973 14909 26007 14943
rect 30573 14909 30607 14943
rect 15577 14841 15611 14875
rect 29193 14841 29227 14875
rect 5825 14773 5859 14807
rect 12528 14773 12562 14807
rect 14933 14773 14967 14807
rect 17325 14773 17359 14807
rect 17969 14773 18003 14807
rect 24685 14773 24719 14807
rect 25329 14773 25363 14807
rect 27261 14773 27295 14807
rect 27905 14773 27939 14807
rect 28549 14773 28583 14807
rect 37841 14773 37875 14807
rect 2237 14569 2271 14603
rect 17233 14569 17267 14603
rect 23857 14569 23891 14603
rect 28917 14569 28951 14603
rect 37381 14569 37415 14603
rect 13645 14501 13679 14535
rect 5549 14433 5583 14467
rect 7573 14433 7607 14467
rect 8493 14433 8527 14467
rect 9689 14433 9723 14467
rect 11069 14433 11103 14467
rect 23029 14433 23063 14467
rect 25513 14433 25547 14467
rect 1593 14365 1627 14399
rect 10977 14365 11011 14399
rect 11621 14365 11655 14399
rect 12265 14365 12299 14399
rect 12909 14365 12943 14399
rect 13001 14365 13035 14399
rect 13553 14365 13587 14399
rect 14565 14365 14599 14399
rect 15209 14365 15243 14399
rect 15853 14365 15887 14399
rect 16497 14365 16531 14399
rect 16589 14365 16623 14399
rect 17141 14365 17175 14399
rect 19441 14365 19475 14399
rect 21741 14365 21775 14399
rect 22845 14365 22879 14399
rect 23765 14365 23799 14399
rect 24593 14365 24627 14399
rect 27537 14365 27571 14399
rect 27997 14365 28031 14399
rect 28825 14365 28859 14399
rect 31217 14365 31251 14399
rect 37565 14365 37599 14399
rect 38025 14365 38059 14399
rect 5641 14297 5675 14331
rect 6561 14297 6595 14331
rect 7665 14297 7699 14331
rect 9321 14297 9355 14331
rect 9413 14297 9447 14331
rect 12357 14297 12391 14331
rect 17877 14297 17911 14331
rect 17969 14297 18003 14331
rect 18889 14297 18923 14331
rect 19717 14297 19751 14331
rect 22293 14297 22327 14331
rect 24685 14297 24719 14331
rect 25789 14297 25823 14331
rect 30113 14297 30147 14331
rect 30205 14297 30239 14331
rect 30757 14297 30791 14331
rect 1777 14229 1811 14263
rect 11713 14229 11747 14263
rect 14657 14229 14691 14263
rect 15301 14229 15335 14263
rect 15945 14229 15979 14263
rect 21189 14229 21223 14263
rect 28089 14229 28123 14263
rect 31309 14229 31343 14263
rect 38209 14229 38243 14263
rect 5917 14025 5951 14059
rect 6837 14025 6871 14059
rect 7481 14025 7515 14059
rect 8125 14025 8159 14059
rect 8769 14025 8803 14059
rect 11069 14025 11103 14059
rect 18613 14025 18647 14059
rect 21465 14025 21499 14059
rect 23857 14025 23891 14059
rect 30021 14025 30055 14059
rect 9505 13957 9539 13991
rect 13369 13957 13403 13991
rect 17141 13957 17175 13991
rect 5825 13889 5859 13923
rect 6745 13889 6779 13923
rect 7389 13889 7423 13923
rect 8033 13889 8067 13923
rect 8677 13889 8711 13923
rect 10977 13889 11011 13923
rect 12265 13889 12299 13923
rect 16129 13889 16163 13923
rect 16865 13889 16899 13923
rect 19073 13889 19107 13923
rect 24869 13889 24903 13923
rect 29929 13889 29963 13923
rect 30573 13889 30607 13923
rect 9413 13821 9447 13855
rect 9689 13821 9723 13855
rect 12357 13821 12391 13855
rect 13093 13821 13127 13855
rect 15117 13821 15151 13855
rect 19165 13821 19199 13855
rect 19717 13821 19751 13855
rect 19993 13821 20027 13855
rect 22109 13821 22143 13855
rect 26617 13821 26651 13855
rect 27169 13821 27203 13855
rect 27445 13821 27479 13855
rect 29193 13821 29227 13855
rect 30665 13821 30699 13855
rect 16221 13685 16255 13719
rect 22372 13685 22406 13719
rect 25132 13685 25166 13719
rect 9229 13481 9263 13515
rect 10057 13481 10091 13515
rect 10701 13481 10735 13515
rect 11976 13481 12010 13515
rect 15945 13481 15979 13515
rect 38117 13481 38151 13515
rect 1777 13413 1811 13447
rect 7573 13345 7607 13379
rect 11713 13345 11747 13379
rect 16497 13345 16531 13379
rect 18521 13345 18555 13379
rect 23397 13345 23431 13379
rect 24777 13345 24811 13379
rect 27997 13345 28031 13379
rect 1593 13277 1627 13311
rect 4353 13277 4387 13311
rect 6837 13277 6871 13311
rect 9137 13277 9171 13311
rect 9965 13277 9999 13311
rect 10609 13277 10643 13311
rect 13737 13277 13771 13311
rect 15209 13277 15243 13311
rect 15301 13277 15335 13311
rect 15853 13277 15887 13311
rect 19441 13277 19475 13311
rect 20085 13277 20119 13311
rect 20729 13277 20763 13311
rect 21373 13277 21407 13311
rect 23857 13277 23891 13311
rect 33333 13277 33367 13311
rect 38301 13277 38335 13311
rect 7665 13209 7699 13243
rect 8585 13209 8619 13243
rect 16773 13209 16807 13243
rect 21649 13209 21683 13243
rect 25053 13209 25087 13243
rect 26801 13209 26835 13243
rect 27261 13209 27295 13243
rect 4353 13141 4387 13175
rect 6929 13141 6963 13175
rect 19533 13141 19567 13175
rect 20177 13141 20211 13175
rect 20821 13141 20855 13175
rect 23949 13141 23983 13175
rect 33149 13141 33183 13175
rect 9505 12937 9539 12971
rect 25237 12937 25271 12971
rect 1869 12869 1903 12903
rect 7573 12869 7607 12903
rect 8493 12869 8527 12903
rect 11805 12869 11839 12903
rect 14473 12869 14507 12903
rect 15669 12869 15703 12903
rect 17785 12869 17819 12903
rect 1685 12801 1719 12835
rect 3985 12801 4019 12835
rect 5089 12801 5123 12835
rect 5825 12801 5859 12835
rect 6745 12801 6779 12835
rect 9413 12801 9447 12835
rect 10517 12801 10551 12835
rect 11713 12801 11747 12835
rect 12449 12801 12483 12835
rect 14933 12801 14967 12835
rect 17509 12801 17543 12835
rect 20545 12801 20579 12835
rect 24501 12801 24535 12835
rect 25145 12801 25179 12835
rect 30757 12801 30791 12835
rect 34897 12801 34931 12835
rect 38117 12801 38151 12835
rect 7481 12733 7515 12767
rect 12725 12733 12759 12767
rect 19533 12733 19567 12767
rect 21281 12733 21315 12767
rect 22017 12733 22051 12767
rect 22293 12733 22327 12767
rect 24041 12733 24075 12767
rect 5917 12665 5951 12699
rect 3801 12597 3835 12631
rect 4905 12597 4939 12631
rect 6837 12597 6871 12631
rect 10609 12597 10643 12631
rect 24593 12597 24627 12631
rect 30849 12597 30883 12631
rect 34713 12597 34747 12631
rect 38209 12597 38243 12631
rect 5089 12393 5123 12427
rect 10701 12393 10735 12427
rect 15748 12393 15782 12427
rect 28641 12393 28675 12427
rect 34161 12393 34195 12427
rect 34989 12393 35023 12427
rect 9229 12257 9263 12291
rect 9873 12257 9907 12291
rect 11713 12257 11747 12291
rect 13737 12257 13771 12291
rect 15485 12257 15519 12291
rect 18705 12257 18739 12291
rect 20177 12257 20211 12291
rect 25697 12257 25731 12291
rect 31861 12257 31895 12291
rect 5089 12189 5123 12223
rect 6929 12189 6963 12223
rect 7757 12189 7791 12223
rect 8401 12189 8435 12223
rect 10609 12189 10643 12223
rect 17969 12189 18003 12223
rect 23213 12189 23247 12223
rect 28549 12189 28583 12223
rect 34069 12189 34103 12223
rect 34897 12189 34931 12223
rect 38117 12189 38151 12223
rect 9321 12121 9355 12155
rect 11989 12121 12023 12155
rect 17509 12121 17543 12155
rect 20453 12121 20487 12155
rect 22201 12121 22235 12155
rect 25973 12121 26007 12155
rect 27721 12121 27755 12155
rect 30849 12121 30883 12155
rect 30941 12121 30975 12155
rect 7021 12053 7055 12087
rect 7849 12053 7883 12087
rect 8493 12053 8527 12087
rect 23305 12053 23339 12087
rect 38209 12053 38243 12087
rect 31585 11849 31619 11883
rect 32597 11849 32631 11883
rect 5457 11781 5491 11815
rect 8401 11781 8435 11815
rect 9958 11781 9992 11815
rect 10885 11781 10919 11815
rect 18613 11781 18647 11815
rect 20361 11781 20395 11815
rect 23765 11781 23799 11815
rect 36829 11781 36863 11815
rect 2513 11713 2547 11747
rect 4169 11713 4203 11747
rect 6009 11713 6043 11747
rect 6929 11713 6963 11747
rect 7573 11713 7607 11747
rect 11713 11713 11747 11747
rect 18337 11713 18371 11747
rect 23489 11713 23523 11747
rect 30205 11713 30239 11747
rect 30849 11713 30883 11747
rect 31493 11713 31527 11747
rect 32505 11713 32539 11747
rect 36093 11713 36127 11747
rect 36737 11713 36771 11747
rect 37473 11713 37507 11747
rect 38117 11713 38151 11747
rect 5365 11645 5399 11679
rect 8309 11645 8343 11679
rect 8585 11645 8619 11679
rect 9873 11645 9907 11679
rect 12357 11645 12391 11679
rect 12633 11645 12667 11679
rect 14565 11645 14599 11679
rect 14841 11645 14875 11679
rect 27169 11645 27203 11679
rect 27445 11645 27479 11679
rect 29193 11645 29227 11679
rect 7665 11577 7699 11611
rect 37565 11577 37599 11611
rect 2329 11509 2363 11543
rect 3985 11509 4019 11543
rect 7021 11509 7055 11543
rect 11805 11509 11839 11543
rect 14105 11509 14139 11543
rect 16313 11509 16347 11543
rect 25237 11509 25271 11543
rect 30297 11509 30331 11543
rect 30941 11509 30975 11543
rect 36185 11509 36219 11543
rect 38209 11509 38243 11543
rect 5181 11305 5215 11339
rect 6837 11305 6871 11339
rect 9229 11305 9263 11339
rect 11529 11305 11563 11339
rect 13737 11305 13771 11339
rect 24041 11305 24075 11339
rect 2329 11237 2363 11271
rect 3341 11237 3375 11271
rect 30481 11237 30515 11271
rect 37473 11237 37507 11271
rect 38301 11237 38335 11271
rect 5825 11169 5859 11203
rect 7481 11169 7515 11203
rect 7849 11169 7883 11203
rect 9781 11169 9815 11203
rect 11989 11169 12023 11203
rect 12265 11169 12299 11203
rect 15209 11169 15243 11203
rect 15485 11169 15519 11203
rect 16957 11169 16991 11203
rect 19441 11169 19475 11203
rect 19717 11169 19751 11203
rect 21465 11169 21499 11203
rect 22293 11169 22327 11203
rect 22569 11169 22603 11203
rect 26249 11169 26283 11203
rect 28273 11169 28307 11203
rect 32873 11169 32907 11203
rect 1593 11101 1627 11135
rect 2513 11101 2547 11135
rect 3249 11101 3283 11135
rect 4169 11101 4203 11135
rect 5365 11101 5399 11135
rect 6745 11101 6779 11135
rect 9137 11101 9171 11135
rect 14281 11101 14315 11135
rect 14381 11101 14415 11135
rect 29929 11101 29963 11135
rect 30389 11101 30423 11135
rect 31033 11101 31067 11135
rect 31677 11101 31711 11135
rect 36185 11101 36219 11135
rect 37381 11101 37415 11135
rect 7573 11033 7607 11067
rect 10057 11033 10091 11067
rect 26525 11033 26559 11067
rect 31769 11033 31803 11067
rect 32597 11033 32631 11067
rect 32689 11033 32723 11067
rect 36277 11033 36311 11067
rect 38117 11033 38151 11067
rect 1777 10965 1811 10999
rect 3985 10965 4019 10999
rect 29745 10965 29779 10999
rect 31125 10965 31159 10999
rect 2237 10761 2271 10795
rect 4629 10761 4663 10795
rect 5917 10761 5951 10795
rect 32597 10761 32631 10795
rect 7205 10693 7239 10727
rect 7757 10693 7791 10727
rect 8401 10693 8435 10727
rect 9321 10693 9355 10727
rect 9965 10693 9999 10727
rect 14473 10693 14507 10727
rect 24501 10693 24535 10727
rect 29469 10693 29503 10727
rect 29561 10693 29595 10727
rect 30481 10693 30515 10727
rect 38301 10693 38335 10727
rect 1777 10625 1811 10659
rect 2421 10625 2455 10659
rect 2881 10625 2915 10659
rect 3525 10625 3559 10659
rect 4537 10625 4571 10659
rect 5181 10625 5215 10659
rect 5825 10625 5859 10659
rect 11713 10625 11747 10659
rect 12449 10625 12483 10659
rect 15117 10625 15151 10659
rect 15577 10625 15611 10659
rect 17417 10625 17451 10659
rect 30941 10625 30975 10659
rect 31585 10625 31619 10659
rect 33241 10625 33275 10659
rect 35449 10625 35483 10659
rect 36093 10625 36127 10659
rect 36737 10625 36771 10659
rect 38117 10625 38151 10659
rect 7113 10557 7147 10591
rect 8309 10557 8343 10591
rect 9873 10557 9907 10591
rect 10149 10557 10183 10591
rect 12725 10557 12759 10591
rect 17693 10557 17727 10591
rect 19441 10557 19475 10591
rect 24225 10557 24259 10591
rect 26249 10557 26283 10591
rect 27169 10557 27203 10591
rect 27445 10557 27479 10591
rect 35541 10557 35575 10591
rect 31033 10489 31067 10523
rect 36829 10489 36863 10523
rect 1593 10421 1627 10455
rect 2973 10421 3007 10455
rect 3617 10421 3651 10455
rect 5273 10421 5307 10455
rect 11805 10421 11839 10455
rect 14933 10421 14967 10455
rect 15669 10421 15703 10455
rect 28917 10421 28951 10455
rect 31677 10421 31711 10455
rect 33333 10421 33367 10455
rect 36185 10421 36219 10455
rect 1593 10217 1627 10251
rect 6285 10217 6319 10251
rect 6929 10217 6963 10251
rect 32321 10217 32355 10251
rect 32965 10217 32999 10251
rect 35633 10217 35667 10251
rect 2237 10149 2271 10183
rect 4353 10149 4387 10183
rect 18889 10149 18923 10183
rect 38117 10149 38151 10183
rect 7573 10081 7607 10115
rect 8493 10081 8527 10115
rect 9781 10081 9815 10115
rect 14289 10081 14323 10115
rect 16313 10081 16347 10115
rect 17417 10081 17451 10115
rect 21097 10081 21131 10115
rect 22845 10081 22879 10115
rect 25513 10081 25547 10115
rect 27537 10081 27571 10115
rect 29929 10081 29963 10115
rect 30113 10081 30147 10115
rect 33609 10081 33643 10115
rect 1777 10013 1811 10047
rect 2421 10013 2455 10047
rect 3433 10013 3467 10047
rect 4261 10013 4295 10047
rect 4905 10013 4939 10047
rect 5733 10013 5767 10047
rect 6193 10013 6227 10047
rect 6837 10013 6871 10047
rect 9505 10013 9539 10047
rect 11713 10013 11747 10047
rect 13737 10013 13771 10047
rect 17141 10013 17175 10047
rect 20361 10013 20395 10047
rect 20821 10013 20855 10047
rect 28733 10013 28767 10047
rect 32229 10013 32263 10047
rect 32873 10013 32907 10047
rect 33517 10013 33551 10047
rect 34161 10013 34195 10047
rect 34897 10013 34931 10047
rect 35541 10013 35575 10047
rect 36921 10013 36955 10047
rect 37381 10013 37415 10047
rect 38301 10013 38335 10047
rect 7665 9945 7699 9979
rect 11989 9945 12023 9979
rect 14565 9945 14599 9979
rect 25789 9945 25823 9979
rect 27997 9945 28031 9979
rect 31769 9945 31803 9979
rect 34989 9945 35023 9979
rect 37473 9945 37507 9979
rect 3249 9877 3283 9911
rect 4997 9877 5031 9911
rect 5549 9877 5583 9911
rect 11253 9877 11287 9911
rect 20177 9877 20211 9911
rect 34253 9877 34287 9911
rect 36737 9877 36771 9911
rect 17509 9673 17543 9707
rect 26617 9673 26651 9707
rect 6837 9605 6871 9639
rect 7389 9605 7423 9639
rect 8033 9605 8067 9639
rect 11989 9605 12023 9639
rect 13737 9605 13771 9639
rect 14841 9605 14875 9639
rect 19257 9605 19291 9639
rect 21005 9605 21039 9639
rect 22293 9605 22327 9639
rect 27445 9605 27479 9639
rect 30297 9605 30331 9639
rect 1777 9537 1811 9571
rect 2605 9537 2639 9571
rect 3249 9537 3283 9571
rect 3893 9537 3927 9571
rect 4537 9537 4571 9571
rect 5181 9537 5215 9571
rect 5825 9537 5859 9571
rect 14565 9537 14599 9571
rect 16865 9537 16899 9571
rect 17693 9537 17727 9571
rect 18153 9537 18187 9571
rect 18981 9537 19015 9571
rect 22017 9537 22051 9571
rect 27169 9537 27203 9571
rect 29377 9537 29411 9571
rect 32321 9537 32355 9571
rect 32965 9537 32999 9571
rect 33609 9537 33643 9571
rect 34253 9537 34287 9571
rect 34897 9537 34931 9571
rect 35817 9537 35851 9571
rect 36461 9537 36495 9571
rect 37473 9537 37507 9571
rect 37565 9537 37599 9571
rect 38301 9537 38335 9571
rect 3985 9469 4019 9503
rect 6745 9469 6779 9503
rect 7941 9469 7975 9503
rect 8585 9469 8619 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 11713 9469 11747 9503
rect 16313 9469 16347 9503
rect 23765 9469 23799 9503
rect 24869 9469 24903 9503
rect 25145 9469 25179 9503
rect 30205 9469 30239 9503
rect 30481 9469 30515 9503
rect 1593 9401 1627 9435
rect 32413 9401 32447 9435
rect 33701 9401 33735 9435
rect 35633 9401 35667 9435
rect 2697 9333 2731 9367
rect 3341 9333 3375 9367
rect 4629 9333 4663 9367
rect 5273 9333 5307 9367
rect 5917 9333 5951 9367
rect 11161 9333 11195 9367
rect 16957 9333 16991 9367
rect 18245 9333 18279 9367
rect 28917 9333 28951 9367
rect 29469 9333 29503 9367
rect 33057 9333 33091 9367
rect 34345 9333 34379 9367
rect 34989 9333 35023 9367
rect 36277 9333 36311 9367
rect 38117 9333 38151 9367
rect 13553 9129 13587 9163
rect 28549 9129 28583 9163
rect 35817 9129 35851 9163
rect 37013 9129 37047 9163
rect 36369 9061 36403 9095
rect 4353 8993 4387 9027
rect 5089 8993 5123 9027
rect 6377 8993 6411 9027
rect 7573 8993 7607 9027
rect 8585 8993 8619 9027
rect 10977 8993 11011 9027
rect 14657 8993 14691 9027
rect 16405 8993 16439 9027
rect 20821 8993 20855 9027
rect 21097 8993 21131 9027
rect 22845 8993 22879 9027
rect 23949 8993 23983 9027
rect 25973 8993 26007 9027
rect 27997 8993 28031 9027
rect 29929 8993 29963 9027
rect 30757 8993 30791 9027
rect 31861 8993 31895 9027
rect 1961 8925 1995 8959
rect 2605 8925 2639 8959
rect 3249 8925 3283 8959
rect 4997 8925 5031 8959
rect 5641 8925 5675 8959
rect 7021 8925 7055 8959
rect 13461 8925 13495 8959
rect 16865 8925 16899 8959
rect 18889 8925 18923 8959
rect 20177 8925 20211 8959
rect 23857 8925 23891 8959
rect 25329 8925 25363 8959
rect 28457 8925 28491 8959
rect 32597 8925 32631 8959
rect 33241 8925 33275 8959
rect 33333 8925 33367 8959
rect 33885 8925 33919 8959
rect 34897 8925 34931 8959
rect 35725 8925 35759 8959
rect 36553 8925 36587 8959
rect 37197 8925 37231 8959
rect 38025 8925 38059 8959
rect 2697 8857 2731 8891
rect 6469 8857 6503 8891
rect 7665 8857 7699 8891
rect 9505 8857 9539 8891
rect 9597 8857 9631 8891
rect 10517 8857 10551 8891
rect 11253 8857 11287 8891
rect 13001 8857 13035 8891
rect 14933 8857 14967 8891
rect 17141 8857 17175 8891
rect 19441 8857 19475 8891
rect 24593 8857 24627 8891
rect 26249 8857 26283 8891
rect 30021 8857 30055 8891
rect 31493 8857 31527 8891
rect 31585 8857 31619 8891
rect 33977 8857 34011 8891
rect 2053 8789 2087 8823
rect 3341 8789 3375 8823
rect 5733 8789 5767 8823
rect 32689 8789 32723 8823
rect 34989 8789 35023 8823
rect 38209 8789 38243 8823
rect 32413 8585 32447 8619
rect 34989 8585 35023 8619
rect 5450 8517 5484 8551
rect 6830 8517 6864 8551
rect 8033 8517 8067 8551
rect 8953 8517 8987 8551
rect 9689 8517 9723 8551
rect 12633 8517 12667 8551
rect 14841 8517 14875 8551
rect 17141 8517 17175 8551
rect 23765 8517 23799 8551
rect 27445 8517 27479 8551
rect 29561 8517 29595 8551
rect 30481 8517 30515 8551
rect 33057 8517 33091 8551
rect 35633 8517 35667 8551
rect 1777 8449 1811 8483
rect 2421 8449 2455 8483
rect 3249 8449 3283 8483
rect 3709 8449 3743 8483
rect 4353 8449 4387 8483
rect 9413 8449 9447 8483
rect 11713 8449 11747 8483
rect 12357 8449 12391 8483
rect 19073 8449 19107 8483
rect 22017 8449 22051 8483
rect 24225 8449 24259 8483
rect 26617 8449 26651 8483
rect 29469 8449 29503 8483
rect 32321 8449 32355 8483
rect 32965 8449 32999 8483
rect 33609 8449 33643 8483
rect 34253 8449 34287 8483
rect 34897 8449 34931 8483
rect 35541 8449 35575 8483
rect 36185 8449 36219 8483
rect 38025 8449 38059 8483
rect 4445 8381 4479 8415
rect 5365 8381 5399 8415
rect 6745 8381 6779 8415
rect 7021 8381 7055 8415
rect 7941 8381 7975 8415
rect 11161 8381 11195 8415
rect 14565 8381 14599 8415
rect 16865 8381 16899 8415
rect 18613 8381 18647 8415
rect 21097 8381 21131 8415
rect 24501 8381 24535 8415
rect 27169 8381 27203 8415
rect 28917 8381 28951 8415
rect 30389 8381 30423 8415
rect 30665 8381 30699 8415
rect 1869 8313 1903 8347
rect 3065 8313 3099 8347
rect 5917 8313 5951 8347
rect 14105 8313 14139 8347
rect 16313 8313 16347 8347
rect 25973 8313 26007 8347
rect 26433 8313 26467 8347
rect 33701 8313 33735 8347
rect 34345 8313 34379 8347
rect 36277 8313 36311 8347
rect 38209 8313 38243 8347
rect 2513 8245 2547 8279
rect 3801 8245 3835 8279
rect 11805 8245 11839 8279
rect 19330 8245 19364 8279
rect 4721 8041 4755 8075
rect 5365 8041 5399 8075
rect 28733 8041 28767 8075
rect 34989 8041 35023 8075
rect 35633 8041 35667 8075
rect 4077 7973 4111 8007
rect 11253 7973 11287 8007
rect 24685 7973 24719 8007
rect 36921 7973 36955 8007
rect 7573 7905 7607 7939
rect 9781 7905 9815 7939
rect 13737 7905 13771 7939
rect 15209 7905 15243 7939
rect 17141 7905 17175 7939
rect 17417 7905 17451 7939
rect 19441 7905 19475 7939
rect 21465 7905 21499 7939
rect 22017 7905 22051 7939
rect 22293 7905 22327 7939
rect 23765 7905 23799 7939
rect 26249 7905 26283 7939
rect 32413 7905 32447 7939
rect 1593 7837 1627 7871
rect 2605 7837 2639 7871
rect 3249 7837 3283 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 5273 7837 5307 7871
rect 9505 7837 9539 7871
rect 11713 7837 11747 7871
rect 14289 7837 14323 7871
rect 14933 7837 14967 7871
rect 24593 7837 24627 7871
rect 25605 7837 25639 7871
rect 28917 7837 28951 7871
rect 30481 7837 30515 7871
rect 32873 7837 32907 7871
rect 33517 7837 33551 7871
rect 34161 7837 34195 7871
rect 34897 7837 34931 7871
rect 35541 7837 35575 7871
rect 36185 7837 36219 7871
rect 36829 7837 36863 7871
rect 38025 7837 38059 7871
rect 6009 7769 6043 7803
rect 6101 7769 6135 7803
rect 7021 7769 7055 7803
rect 7665 7769 7699 7803
rect 8585 7769 8619 7803
rect 11989 7769 12023 7803
rect 19717 7769 19751 7803
rect 26525 7769 26559 7803
rect 28273 7769 28307 7803
rect 29745 7769 29779 7803
rect 31401 7769 31435 7803
rect 31493 7769 31527 7803
rect 33609 7769 33643 7803
rect 1777 7701 1811 7735
rect 2697 7701 2731 7735
rect 3341 7701 3375 7735
rect 14381 7701 14415 7735
rect 16681 7701 16715 7735
rect 18889 7701 18923 7735
rect 25697 7701 25731 7735
rect 32965 7701 32999 7735
rect 34253 7701 34287 7735
rect 36277 7701 36311 7735
rect 38209 7701 38243 7735
rect 3985 7497 4019 7531
rect 4629 7497 4663 7531
rect 11805 7497 11839 7531
rect 17417 7497 17451 7531
rect 20913 7497 20947 7531
rect 23765 7497 23799 7531
rect 25973 7497 26007 7531
rect 31677 7497 31711 7531
rect 34161 7497 34195 7531
rect 37565 7497 37599 7531
rect 2145 7429 2179 7463
rect 6837 7429 6871 7463
rect 7941 7429 7975 7463
rect 8033 7429 8067 7463
rect 8953 7429 8987 7463
rect 12633 7429 12667 7463
rect 14381 7429 14415 7463
rect 15577 7429 15611 7463
rect 19809 7429 19843 7463
rect 22293 7429 22327 7463
rect 27445 7429 27479 7463
rect 29653 7429 29687 7463
rect 32413 7429 32447 7463
rect 32505 7429 32539 7463
rect 36185 7429 36219 7463
rect 2053 7361 2087 7395
rect 2789 7361 2823 7395
rect 3249 7361 3283 7395
rect 3893 7361 3927 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 11713 7361 11747 7395
rect 14841 7361 14875 7395
rect 16957 7361 16991 7395
rect 20269 7361 20303 7395
rect 21097 7361 21131 7395
rect 22017 7361 22051 7395
rect 26617 7361 26651 7395
rect 27158 7361 27192 7395
rect 29377 7361 29411 7395
rect 31585 7361 31619 7395
rect 33057 7361 33091 7395
rect 33517 7361 33551 7395
rect 34805 7361 34839 7395
rect 36093 7361 36127 7395
rect 36921 7361 36955 7395
rect 37473 7361 37507 7395
rect 38301 7361 38335 7395
rect 5273 7293 5307 7327
rect 6745 7293 6779 7327
rect 7021 7293 7055 7327
rect 9413 7293 9447 7327
rect 9689 7293 9723 7327
rect 12357 7293 12391 7327
rect 17785 7293 17819 7327
rect 18061 7293 18095 7327
rect 24225 7293 24259 7327
rect 24501 7293 24535 7327
rect 35449 7293 35483 7327
rect 5917 7225 5951 7259
rect 11161 7225 11195 7259
rect 17049 7225 17083 7259
rect 26433 7225 26467 7259
rect 34897 7225 34931 7259
rect 2605 7157 2639 7191
rect 3341 7157 3375 7191
rect 20361 7157 20395 7191
rect 28917 7157 28951 7191
rect 31125 7157 31159 7191
rect 33609 7157 33643 7191
rect 36737 7157 36771 7191
rect 38117 7157 38151 7191
rect 4353 6953 4387 6987
rect 7100 6953 7134 6987
rect 16478 6953 16512 6987
rect 20992 6953 21026 6987
rect 26512 6953 26546 6987
rect 28733 6953 28767 6987
rect 30008 6953 30042 6987
rect 2697 6817 2731 6851
rect 9229 6817 9263 6851
rect 11069 6817 11103 6851
rect 15025 6817 15059 6851
rect 16221 6817 16255 6851
rect 23305 6817 23339 6851
rect 26249 6817 26283 6851
rect 28273 6817 28307 6851
rect 29745 6817 29779 6851
rect 32045 6817 32079 6851
rect 32413 6817 32447 6851
rect 34897 6817 34931 6851
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 3249 6749 3283 6783
rect 4261 6749 4295 6783
rect 5089 6749 5123 6783
rect 5549 6749 5583 6783
rect 6193 6749 6227 6783
rect 6837 6749 6871 6783
rect 13093 6749 13127 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 18889 6749 18923 6783
rect 19441 6749 19475 6783
rect 20729 6749 20763 6783
rect 22753 6749 22787 6783
rect 23213 6749 23247 6783
rect 23857 6749 23891 6783
rect 24593 6749 24627 6783
rect 25237 6749 25271 6783
rect 28917 6749 28951 6783
rect 33517 6749 33551 6783
rect 33609 6749 33643 6783
rect 34161 6749 34195 6783
rect 35541 6749 35575 6783
rect 36185 6749 36219 6783
rect 36829 6749 36863 6783
rect 38025 6749 38059 6783
rect 3341 6681 3375 6715
rect 9597 6681 9631 6715
rect 9689 6681 9723 6715
rect 10609 6681 10643 6715
rect 11345 6681 11379 6715
rect 14289 6681 14323 6715
rect 18245 6681 18279 6715
rect 32137 6681 32171 6715
rect 2053 6613 2087 6647
rect 4905 6613 4939 6647
rect 5641 6613 5675 6647
rect 6285 6613 6319 6647
rect 8585 6613 8619 6647
rect 18705 6613 18739 6647
rect 19625 6613 19659 6647
rect 23949 6613 23983 6647
rect 24685 6613 24719 6647
rect 25329 6613 25363 6647
rect 31493 6613 31527 6647
rect 34253 6613 34287 6647
rect 35633 6613 35667 6647
rect 36277 6613 36311 6647
rect 36921 6613 36955 6647
rect 38209 6613 38243 6647
rect 3709 6409 3743 6443
rect 11161 6409 11195 6443
rect 23765 6409 23799 6443
rect 28917 6409 28951 6443
rect 36185 6409 36219 6443
rect 36829 6409 36863 6443
rect 5089 6341 5123 6375
rect 6009 6341 6043 6375
rect 7481 6341 7515 6375
rect 9689 6341 9723 6375
rect 12541 6341 12575 6375
rect 15393 6341 15427 6375
rect 17141 6341 17175 6375
rect 32321 6341 32355 6375
rect 34046 6341 34080 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 2973 6273 3007 6307
rect 3617 6273 3651 6307
rect 4261 6273 4295 6307
rect 6561 6273 6595 6307
rect 7205 6273 7239 6307
rect 9413 6273 9447 6307
rect 12265 6273 12299 6307
rect 14749 6273 14783 6307
rect 21005 6273 21039 6307
rect 26433 6273 26467 6307
rect 27169 6273 27203 6307
rect 29377 6273 29411 6307
rect 31769 6273 31803 6307
rect 33517 6273 33551 6307
rect 36093 6273 36127 6307
rect 36737 6273 36771 6307
rect 38117 6273 38151 6307
rect 4353 6205 4387 6239
rect 4997 6205 5031 6239
rect 14289 6205 14323 6239
rect 16221 6205 16255 6239
rect 17049 6205 17083 6239
rect 17325 6205 17359 6239
rect 18521 6205 18555 6239
rect 18797 6205 18831 6239
rect 20545 6205 20579 6239
rect 22017 6205 22051 6239
rect 22293 6205 22327 6239
rect 24225 6205 24259 6239
rect 24501 6205 24535 6239
rect 27445 6205 27479 6239
rect 29653 6205 29687 6239
rect 32229 6205 32263 6239
rect 32505 6205 32539 6239
rect 33977 6205 34011 6239
rect 34253 6205 34287 6239
rect 35449 6205 35483 6239
rect 1777 6137 1811 6171
rect 2421 6137 2455 6171
rect 6653 6137 6687 6171
rect 3065 6069 3099 6103
rect 8953 6069 8987 6103
rect 14841 6069 14875 6103
rect 21097 6069 21131 6103
rect 25973 6069 26007 6103
rect 26525 6069 26559 6103
rect 31125 6069 31159 6103
rect 31585 6069 31619 6103
rect 38209 6069 38243 6103
rect 7100 5865 7134 5899
rect 35633 5865 35667 5899
rect 1869 5797 1903 5831
rect 3341 5797 3375 5831
rect 8585 5797 8619 5831
rect 11253 5797 11287 5831
rect 16405 5797 16439 5831
rect 28641 5797 28675 5831
rect 34161 5797 34195 5831
rect 34989 5797 35023 5831
rect 36277 5797 36311 5831
rect 9505 5729 9539 5763
rect 9781 5729 9815 5763
rect 11713 5729 11747 5763
rect 11989 5729 12023 5763
rect 14657 5729 14691 5763
rect 16865 5729 16899 5763
rect 20453 5729 20487 5763
rect 23673 5729 23707 5763
rect 25145 5729 25179 5763
rect 26157 5729 26191 5763
rect 29745 5729 29779 5763
rect 32045 5729 32079 5763
rect 2329 5661 2363 5695
rect 3249 5661 3283 5695
rect 4261 5661 4295 5695
rect 6837 5661 6871 5695
rect 19717 5661 19751 5695
rect 22937 5661 22971 5695
rect 24869 5661 24903 5695
rect 28825 5661 28859 5695
rect 34897 5661 34931 5695
rect 35541 5661 35575 5695
rect 36185 5661 36219 5695
rect 37289 5661 37323 5695
rect 38025 5661 38059 5695
rect 1685 5593 1719 5627
rect 5365 5593 5399 5627
rect 5457 5593 5491 5627
rect 6377 5593 6411 5627
rect 13737 5593 13771 5627
rect 14933 5593 14967 5627
rect 17141 5593 17175 5627
rect 18889 5593 18923 5627
rect 20729 5593 20763 5627
rect 22477 5593 22511 5627
rect 26433 5593 26467 5627
rect 28181 5593 28215 5627
rect 30021 5593 30055 5627
rect 32137 5593 32171 5627
rect 33057 5593 33091 5627
rect 33609 5593 33643 5627
rect 33701 5593 33735 5627
rect 2513 5525 2547 5559
rect 4353 5525 4387 5559
rect 19901 5525 19935 5559
rect 31493 5525 31527 5559
rect 37473 5525 37507 5559
rect 38209 5525 38243 5559
rect 7021 5321 7055 5355
rect 19165 5321 19199 5355
rect 3525 5253 3559 5287
rect 4997 5253 5031 5287
rect 5089 5253 5123 5287
rect 6929 5253 6963 5287
rect 9965 5253 9999 5287
rect 10057 5253 10091 5287
rect 14841 5253 14875 5287
rect 18797 5253 18831 5287
rect 24593 5253 24627 5287
rect 27445 5253 27479 5287
rect 32321 5253 32355 5287
rect 33517 5253 33551 5287
rect 33977 5253 34011 5287
rect 34069 5253 34103 5287
rect 1593 5185 1627 5219
rect 2329 5185 2363 5219
rect 7573 5185 7607 5219
rect 11713 5185 11747 5219
rect 19441 5185 19475 5219
rect 21465 5185 21499 5219
rect 29193 5185 29227 5219
rect 35449 5185 35483 5219
rect 36645 5185 36679 5219
rect 3433 5117 3467 5151
rect 4445 5117 4479 5151
rect 5273 5117 5307 5151
rect 7757 5101 7791 5135
rect 9413 5117 9447 5151
rect 10977 5117 11011 5151
rect 11989 5117 12023 5151
rect 13737 5117 13771 5151
rect 14565 5117 14599 5151
rect 16773 5117 16807 5151
rect 19717 5117 19751 5151
rect 22017 5117 22051 5151
rect 22293 5117 22327 5151
rect 24317 5117 24351 5151
rect 26341 5117 26375 5151
rect 27169 5117 27203 5151
rect 29653 5117 29687 5151
rect 29929 5117 29963 5151
rect 32229 5117 32263 5151
rect 32505 5117 32539 5151
rect 34897 5117 34931 5151
rect 37473 5117 37507 5151
rect 37749 5117 37783 5151
rect 16313 5049 16347 5083
rect 23765 5049 23799 5083
rect 35541 5049 35575 5083
rect 1777 4981 1811 5015
rect 2513 4981 2547 5015
rect 17036 4981 17070 5015
rect 31401 4981 31435 5015
rect 36829 4981 36863 5015
rect 1777 4777 1811 4811
rect 2513 4777 2547 4811
rect 4077 4777 4111 4811
rect 8585 4777 8619 4811
rect 16313 4777 16347 4811
rect 6377 4709 6411 4743
rect 29101 4709 29135 4743
rect 4629 4641 4663 4675
rect 9505 4641 9539 4675
rect 16865 4641 16899 4675
rect 21189 4641 21223 4675
rect 25329 4641 25363 4675
rect 27997 4641 28031 4675
rect 29745 4641 29779 4675
rect 31953 4641 31987 4675
rect 35173 4641 35207 4675
rect 37473 4641 37507 4675
rect 3065 4573 3099 4607
rect 3985 4573 4019 4607
rect 6837 4573 6871 4607
rect 11253 4573 11287 4607
rect 14565 4573 14599 4607
rect 19441 4573 19475 4607
rect 20913 4573 20947 4607
rect 23397 4573 23431 4607
rect 24593 4573 24627 4607
rect 25973 4573 26007 4607
rect 34161 4573 34195 4607
rect 34253 4573 34287 4607
rect 34897 4573 34931 4607
rect 36737 4573 36771 4607
rect 37749 4573 37783 4607
rect 1685 4505 1719 4539
rect 2421 4505 2455 4539
rect 4905 4505 4939 4539
rect 7113 4505 7147 4539
rect 9229 4505 9263 4539
rect 9321 4505 9355 4539
rect 11529 4505 11563 4539
rect 13277 4505 13311 4539
rect 14841 4505 14875 4539
rect 17141 4505 17175 4539
rect 18889 4505 18923 4539
rect 20177 4505 20211 4539
rect 22937 4505 22971 4539
rect 26249 4505 26283 4539
rect 28549 4505 28583 4539
rect 28641 4505 28675 4539
rect 30021 4505 30055 4539
rect 32229 4505 32263 4539
rect 3249 4437 3283 4471
rect 23581 4437 23615 4471
rect 31493 4437 31527 4471
rect 33701 4437 33735 4471
rect 36921 4437 36955 4471
rect 33885 4233 33919 4267
rect 2881 4165 2915 4199
rect 4537 4165 4571 4199
rect 7021 4165 7055 4199
rect 11713 4165 11747 4199
rect 15117 4165 15151 4199
rect 16129 4165 16163 4199
rect 17417 4165 17451 4199
rect 22201 4165 22235 4199
rect 34621 4165 34655 4199
rect 34713 4165 34747 4199
rect 1593 4097 1627 4131
rect 8953 4097 8987 4131
rect 20821 4097 20855 4131
rect 23857 4097 23891 4131
rect 26341 4097 26375 4131
rect 29653 4097 29687 4131
rect 32137 4097 32171 4131
rect 34161 4097 34195 4131
rect 36185 4097 36219 4131
rect 37749 4097 37783 4131
rect 2789 4029 2823 4063
rect 3801 4029 3835 4063
rect 4261 4029 4295 4063
rect 6745 4029 6779 4063
rect 9137 4029 9171 4063
rect 10793 4029 10827 4063
rect 12449 4029 12483 4063
rect 13093 4029 13127 4063
rect 13369 4029 13403 4063
rect 16313 4029 16347 4063
rect 18061 4029 18095 4063
rect 18337 4029 18371 4063
rect 20085 4029 20119 4063
rect 20545 4029 20579 4063
rect 22109 4029 22143 4063
rect 23121 4029 23155 4063
rect 24133 4029 24167 4063
rect 25881 4029 25915 4063
rect 27169 4029 27203 4063
rect 29193 4029 29227 4063
rect 29929 4029 29963 4063
rect 31401 4029 31435 4063
rect 32413 4029 32447 4063
rect 35633 4029 35667 4063
rect 37473 4029 37507 4063
rect 6009 3961 6043 3995
rect 26433 3961 26467 3995
rect 1777 3893 1811 3927
rect 8493 3893 8527 3927
rect 17509 3893 17543 3927
rect 27432 3893 27466 3927
rect 36369 3893 36403 3927
rect 6377 3689 6411 3723
rect 38209 3689 38243 3723
rect 3341 3621 3375 3655
rect 2789 3553 2823 3587
rect 4629 3553 4663 3587
rect 7113 3553 7147 3587
rect 9229 3553 9263 3587
rect 10057 3553 10091 3587
rect 13093 3553 13127 3587
rect 14289 3553 14323 3587
rect 17141 3553 17175 3587
rect 20269 3553 20303 3587
rect 22017 3553 22051 3587
rect 22569 3553 22603 3587
rect 22937 3553 22971 3587
rect 25789 3553 25823 3587
rect 30757 3553 30791 3587
rect 30941 3553 30975 3587
rect 32597 3553 32631 3587
rect 33149 3553 33183 3587
rect 35265 3553 35299 3587
rect 36553 3553 36587 3587
rect 37565 3553 37599 3587
rect 1961 3485 1995 3519
rect 3985 3485 4019 3519
rect 6837 3485 6871 3519
rect 11069 3485 11103 3519
rect 13553 3485 13587 3519
rect 16865 3485 16899 3519
rect 19993 3485 20027 3519
rect 24593 3485 24627 3519
rect 27813 3485 27847 3519
rect 28273 3485 28307 3519
rect 30021 3485 30055 3519
rect 38117 3485 38151 3519
rect 2881 3417 2915 3451
rect 4905 3417 4939 3451
rect 9321 3417 9355 3451
rect 11345 3417 11379 3451
rect 14565 3417 14599 3451
rect 16313 3417 16347 3451
rect 18889 3417 18923 3451
rect 22661 3417 22695 3451
rect 26065 3417 26099 3451
rect 29101 3417 29135 3451
rect 33241 3417 33275 3451
rect 34161 3417 34195 3451
rect 34989 3417 35023 3451
rect 35081 3417 35115 3451
rect 36645 3417 36679 3451
rect 2145 3349 2179 3383
rect 4077 3349 4111 3383
rect 8585 3349 8619 3383
rect 13645 3349 13679 3383
rect 24777 3349 24811 3383
rect 30205 3349 30239 3383
rect 2237 3145 2271 3179
rect 26525 3145 26559 3179
rect 2145 3077 2179 3111
rect 4537 3077 4571 3111
rect 7376 3077 7410 3111
rect 19533 3077 19567 3111
rect 21281 3077 21315 3111
rect 24501 3077 24535 3111
rect 27445 3077 27479 3111
rect 34621 3077 34655 3111
rect 34713 3077 34747 3111
rect 35633 3077 35667 3111
rect 2789 3009 2823 3043
rect 3525 3009 3559 3043
rect 4261 3009 4295 3043
rect 11805 3009 11839 3043
rect 14289 3009 14323 3043
rect 19257 3009 19291 3043
rect 22017 3009 22051 3043
rect 24225 3009 24259 3043
rect 26433 3009 26467 3043
rect 36369 3009 36403 3043
rect 37749 3009 37783 3043
rect 6009 2941 6043 2975
rect 7113 2941 7147 2975
rect 9321 2941 9355 2975
rect 9597 2941 9631 2975
rect 13829 2941 13863 2975
rect 14565 2941 14599 2975
rect 16313 2941 16347 2975
rect 16865 2941 16899 2975
rect 17141 2941 17175 2975
rect 22293 2941 22327 2975
rect 25973 2941 26007 2975
rect 27169 2941 27203 2975
rect 29193 2941 29227 2975
rect 29653 2941 29687 2975
rect 29929 2941 29963 2975
rect 31401 2941 31435 2975
rect 32321 2941 32355 2975
rect 32597 2941 32631 2975
rect 36093 2941 36127 2975
rect 37473 2941 37507 2975
rect 2973 2805 3007 2839
rect 3709 2805 3743 2839
rect 8861 2805 8895 2839
rect 11069 2805 11103 2839
rect 12062 2805 12096 2839
rect 18613 2805 18647 2839
rect 23765 2805 23799 2839
rect 34069 2805 34103 2839
rect 1869 2601 1903 2635
rect 28917 2601 28951 2635
rect 2329 2533 2363 2567
rect 2605 2533 2639 2567
rect 4353 2533 4387 2567
rect 11161 2533 11195 2567
rect 15945 2533 15979 2567
rect 34069 2533 34103 2567
rect 6009 2465 6043 2499
rect 6837 2465 6871 2499
rect 7113 2465 7147 2499
rect 8585 2465 8619 2499
rect 9413 2465 9447 2499
rect 11713 2465 11747 2499
rect 14197 2465 14231 2499
rect 16865 2465 16899 2499
rect 19441 2465 19475 2499
rect 22017 2465 22051 2499
rect 22293 2465 22327 2499
rect 24593 2465 24627 2499
rect 27169 2465 27203 2499
rect 29745 2465 29779 2499
rect 32321 2465 32355 2499
rect 34897 2465 34931 2499
rect 35173 2465 35207 2499
rect 37473 2465 37507 2499
rect 37749 2465 37783 2499
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 3157 2397 3191 2431
rect 4169 2397 4203 2431
rect 4997 2329 5031 2363
rect 5089 2329 5123 2363
rect 9689 2329 9723 2363
rect 11989 2329 12023 2363
rect 13737 2329 13771 2363
rect 14473 2329 14507 2363
rect 17141 2329 17175 2363
rect 18889 2329 18923 2363
rect 19717 2329 19751 2363
rect 21465 2329 21499 2363
rect 24869 2329 24903 2363
rect 27445 2329 27479 2363
rect 30021 2329 30055 2363
rect 32597 2329 32631 2363
rect 3341 2261 3375 2295
rect 16313 2261 16347 2295
rect 23765 2261 23799 2295
rect 26341 2261 26375 2295
rect 31493 2261 31527 2295
rect 36645 2261 36679 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 14 37272 20 37324
rect 72 37312 78 37324
rect 2958 37312 2964 37324
rect 72 37284 2964 37312
rect 72 37272 78 37284
rect 2958 37272 2964 37284
rect 3016 37272 3022 37324
rect 10318 37312 10324 37324
rect 10279 37284 10324 37312
rect 10318 37272 10324 37284
rect 10376 37272 10382 37324
rect 15470 37312 15476 37324
rect 15431 37284 15476 37312
rect 15470 37272 15476 37284
rect 15528 37272 15534 37324
rect 16850 37272 16856 37324
rect 16908 37312 16914 37324
rect 17129 37315 17187 37321
rect 17129 37312 17141 37315
rect 16908 37284 17141 37312
rect 16908 37272 16914 37284
rect 17129 37281 17141 37284
rect 17175 37281 17187 37315
rect 17129 37275 17187 37281
rect 18141 37315 18199 37321
rect 18141 37281 18153 37315
rect 18187 37312 18199 37315
rect 19426 37312 19432 37324
rect 18187 37284 19432 37312
rect 18187 37281 18199 37284
rect 18141 37275 18199 37281
rect 19426 37272 19432 37284
rect 19484 37272 19490 37324
rect 23661 37315 23719 37321
rect 23661 37281 23673 37315
rect 23707 37312 23719 37315
rect 23842 37312 23848 37324
rect 23707 37284 23848 37312
rect 23707 37281 23719 37284
rect 23661 37275 23719 37281
rect 23842 37272 23848 37284
rect 23900 37272 23906 37324
rect 26329 37315 26387 37321
rect 26329 37281 26341 37315
rect 26375 37312 26387 37315
rect 26510 37312 26516 37324
rect 26375 37284 26516 37312
rect 26375 37281 26387 37284
rect 26329 37275 26387 37281
rect 26510 37272 26516 37284
rect 26568 37272 26574 37324
rect 31570 37272 31576 37324
rect 31628 37312 31634 37324
rect 32309 37315 32367 37321
rect 32309 37312 32321 37315
rect 31628 37284 32321 37312
rect 31628 37272 31634 37284
rect 32309 37281 32321 37284
rect 32355 37281 32367 37315
rect 32309 37275 32367 37281
rect 37461 37315 37519 37321
rect 37461 37281 37473 37315
rect 37507 37312 37519 37315
rect 38010 37312 38016 37324
rect 37507 37284 38016 37312
rect 37507 37281 37519 37284
rect 37461 37275 37519 37281
rect 38010 37272 38016 37284
rect 38068 37272 38074 37324
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37213 1915 37247
rect 1857 37207 1915 37213
rect 2869 37247 2927 37253
rect 2869 37213 2881 37247
rect 2915 37244 2927 37247
rect 3050 37244 3056 37256
rect 2915 37216 3056 37244
rect 2915 37213 2927 37216
rect 2869 37207 2927 37213
rect 1872 37176 1900 37207
rect 3050 37204 3056 37216
rect 3108 37204 3114 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4157 37247 4215 37253
rect 4157 37244 4169 37247
rect 3292 37216 4169 37244
rect 3292 37204 3298 37216
rect 4157 37213 4169 37216
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4617 37247 4675 37253
rect 4617 37213 4629 37247
rect 4663 37244 4675 37247
rect 5074 37244 5080 37256
rect 4663 37216 5080 37244
rect 4663 37213 4675 37216
rect 4617 37207 4675 37213
rect 5074 37204 5080 37216
rect 5132 37204 5138 37256
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5537 37247 5595 37253
rect 5537 37244 5549 37247
rect 5224 37216 5549 37244
rect 5224 37204 5230 37216
rect 5537 37213 5549 37216
rect 5583 37213 5595 37247
rect 6546 37244 6552 37256
rect 6507 37216 6552 37244
rect 5537 37207 5595 37213
rect 6546 37204 6552 37216
rect 6604 37204 6610 37256
rect 7834 37244 7840 37256
rect 7795 37216 7840 37244
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9732 37216 9873 37244
rect 9732 37204 9738 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 10597 37247 10655 37253
rect 10597 37213 10609 37247
rect 10643 37244 10655 37247
rect 10643 37216 10732 37244
rect 10643 37213 10655 37216
rect 10597 37207 10655 37213
rect 10704 37188 10732 37216
rect 12158 37204 12164 37256
rect 12216 37244 12222 37256
rect 12345 37247 12403 37253
rect 12345 37244 12357 37247
rect 12216 37216 12357 37244
rect 12216 37204 12222 37216
rect 12345 37213 12357 37216
rect 12391 37213 12403 37247
rect 12345 37207 12403 37213
rect 12986 37204 12992 37256
rect 13044 37244 13050 37256
rect 14277 37247 14335 37253
rect 14277 37244 14289 37247
rect 13044 37216 14289 37244
rect 13044 37204 13050 37216
rect 14277 37213 14289 37216
rect 14323 37213 14335 37247
rect 15746 37244 15752 37256
rect 15707 37216 15752 37244
rect 14277 37207 14335 37213
rect 15746 37204 15752 37216
rect 15804 37204 15810 37256
rect 16114 37204 16120 37256
rect 16172 37244 16178 37256
rect 16945 37247 17003 37253
rect 16945 37244 16957 37247
rect 16172 37216 16957 37244
rect 16172 37204 16178 37216
rect 16945 37213 16957 37216
rect 16991 37213 17003 37247
rect 16945 37207 17003 37213
rect 17957 37247 18015 37253
rect 17957 37213 17969 37247
rect 18003 37244 18015 37247
rect 18046 37244 18052 37256
rect 18003 37216 18052 37244
rect 18003 37213 18015 37216
rect 17957 37207 18015 37213
rect 18046 37204 18052 37216
rect 18104 37204 18110 37256
rect 18598 37244 18604 37256
rect 18559 37216 18604 37244
rect 18598 37204 18604 37216
rect 18656 37204 18662 37256
rect 19978 37244 19984 37256
rect 19939 37216 19984 37244
rect 19978 37204 19984 37216
rect 20036 37204 20042 37256
rect 20717 37247 20775 37253
rect 20717 37213 20729 37247
rect 20763 37244 20775 37247
rect 21174 37244 21180 37256
rect 20763 37216 21180 37244
rect 20763 37213 20775 37216
rect 20717 37207 20775 37213
rect 21174 37204 21180 37216
rect 21232 37204 21238 37256
rect 21266 37204 21272 37256
rect 21324 37244 21330 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 21324 37216 22201 37244
rect 21324 37204 21330 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22649 37247 22707 37253
rect 22649 37244 22661 37247
rect 22520 37216 22661 37244
rect 22520 37204 22526 37216
rect 22649 37213 22661 37216
rect 22695 37213 22707 37247
rect 22649 37207 22707 37213
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23477 37247 23535 37253
rect 23477 37244 23489 37247
rect 23256 37216 23489 37244
rect 23256 37204 23262 37216
rect 23477 37213 23489 37216
rect 23523 37213 23535 37247
rect 23477 37207 23535 37213
rect 24026 37204 24032 37256
rect 24084 37244 24090 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 24084 37216 24593 37244
rect 24084 37204 24090 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 25317 37247 25375 37253
rect 25317 37213 25329 37247
rect 25363 37213 25375 37247
rect 25317 37207 25375 37213
rect 10502 37176 10508 37188
rect 1872 37148 10508 37176
rect 10502 37136 10508 37148
rect 10560 37136 10566 37188
rect 10686 37136 10692 37188
rect 10744 37176 10750 37188
rect 13354 37176 13360 37188
rect 10744 37148 13360 37176
rect 10744 37136 10750 37148
rect 13354 37136 13360 37148
rect 13412 37136 13418 37188
rect 24394 37176 24400 37188
rect 22020 37148 24400 37176
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 3053 37111 3111 37117
rect 3053 37108 3065 37111
rect 2832 37080 3065 37108
rect 2832 37068 2838 37080
rect 3053 37077 3065 37080
rect 3099 37077 3111 37111
rect 3970 37108 3976 37120
rect 3931 37080 3976 37108
rect 3053 37071 3111 37077
rect 3970 37068 3976 37080
rect 4028 37068 4034 37120
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4801 37111 4859 37117
rect 4801 37108 4813 37111
rect 4672 37080 4813 37108
rect 4672 37068 4678 37080
rect 4801 37077 4813 37080
rect 4847 37077 4859 37111
rect 5350 37108 5356 37120
rect 5311 37080 5356 37108
rect 4801 37071 4859 37077
rect 5350 37068 5356 37080
rect 5408 37068 5414 37120
rect 5810 37068 5816 37120
rect 5868 37108 5874 37120
rect 6733 37111 6791 37117
rect 6733 37108 6745 37111
rect 5868 37080 6745 37108
rect 5868 37068 5874 37080
rect 6733 37077 6745 37080
rect 6779 37077 6791 37111
rect 6733 37071 6791 37077
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 8021 37071 8079 37077
rect 9677 37111 9735 37117
rect 9677 37077 9689 37111
rect 9723 37108 9735 37111
rect 10962 37108 10968 37120
rect 9723 37080 10968 37108
rect 9723 37077 9735 37080
rect 9677 37071 9735 37077
rect 10962 37068 10968 37080
rect 11020 37068 11026 37120
rect 12434 37068 12440 37120
rect 12492 37108 12498 37120
rect 12529 37111 12587 37117
rect 12529 37108 12541 37111
rect 12492 37080 12541 37108
rect 12492 37068 12498 37080
rect 12529 37077 12541 37080
rect 12575 37077 12587 37111
rect 12529 37071 12587 37077
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13596 37080 14473 37108
rect 13596 37068 13602 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 14461 37071 14519 37077
rect 18690 37068 18696 37120
rect 18748 37108 18754 37120
rect 18785 37111 18843 37117
rect 18785 37108 18797 37111
rect 18748 37080 18797 37108
rect 18748 37068 18754 37080
rect 18785 37077 18797 37080
rect 18831 37077 18843 37111
rect 18785 37071 18843 37077
rect 20070 37068 20076 37120
rect 20128 37108 20134 37120
rect 20165 37111 20223 37117
rect 20165 37108 20177 37111
rect 20128 37080 20177 37108
rect 20128 37068 20134 37080
rect 20165 37077 20177 37080
rect 20211 37077 20223 37111
rect 20165 37071 20223 37077
rect 20714 37068 20720 37120
rect 20772 37108 20778 37120
rect 22020 37117 22048 37148
rect 24394 37136 24400 37148
rect 24452 37136 24458 37188
rect 25332 37176 25360 37207
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26145 37247 26203 37253
rect 26145 37244 26157 37247
rect 25832 37216 26157 37244
rect 25832 37204 25838 37216
rect 26145 37213 26157 37216
rect 26191 37213 26203 37247
rect 26145 37207 26203 37213
rect 27157 37247 27215 37253
rect 27157 37213 27169 37247
rect 27203 37244 27215 37247
rect 27522 37244 27528 37256
rect 27203 37216 27528 37244
rect 27203 37213 27215 37216
rect 27157 37207 27215 37213
rect 27522 37204 27528 37216
rect 27580 37204 27586 37256
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 28077 37247 28135 37253
rect 28077 37244 28089 37247
rect 27764 37216 28089 37244
rect 27764 37204 27770 37216
rect 28077 37213 28089 37216
rect 28123 37213 28135 37247
rect 28077 37207 28135 37213
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29181 37247 29239 37253
rect 29181 37244 29193 37247
rect 29052 37216 29193 37244
rect 29052 37204 29058 37216
rect 29181 37213 29193 37216
rect 29227 37213 29239 37247
rect 29730 37244 29736 37256
rect 29691 37216 29736 37244
rect 29181 37207 29239 37213
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 30432 37216 30665 37244
rect 30432 37204 30438 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 30653 37207 30711 37213
rect 30742 37204 30748 37256
rect 30800 37244 30806 37256
rect 32585 37247 32643 37253
rect 32585 37244 32597 37247
rect 30800 37216 32597 37244
rect 30800 37204 30806 37216
rect 32585 37213 32597 37216
rect 32631 37213 32643 37247
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 32585 37207 32643 37213
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34848 37216 34897 37244
rect 34848 37204 34854 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 34974 37204 34980 37256
rect 35032 37244 35038 37256
rect 35713 37247 35771 37253
rect 35713 37244 35725 37247
rect 35032 37216 35725 37244
rect 35032 37204 35038 37216
rect 35713 37213 35725 37216
rect 35759 37213 35771 37247
rect 35713 37207 35771 37213
rect 36262 37204 36268 37256
rect 36320 37244 36326 37256
rect 36357 37247 36415 37253
rect 36357 37244 36369 37247
rect 36320 37216 36369 37244
rect 36320 37204 36326 37216
rect 36357 37213 36369 37216
rect 36403 37213 36415 37247
rect 36357 37207 36415 37213
rect 37737 37247 37795 37253
rect 37737 37213 37749 37247
rect 37783 37213 37795 37247
rect 37737 37207 37795 37213
rect 24504 37148 25360 37176
rect 20901 37111 20959 37117
rect 20901 37108 20913 37111
rect 20772 37080 20913 37108
rect 20772 37068 20778 37080
rect 20901 37077 20913 37080
rect 20947 37077 20959 37111
rect 20901 37071 20959 37077
rect 22005 37111 22063 37117
rect 22005 37077 22017 37111
rect 22051 37077 22063 37111
rect 22005 37071 22063 37077
rect 22554 37068 22560 37120
rect 22612 37108 22618 37120
rect 22833 37111 22891 37117
rect 22833 37108 22845 37111
rect 22612 37080 22845 37108
rect 22612 37068 22618 37080
rect 22833 37077 22845 37080
rect 22879 37077 22891 37111
rect 22833 37071 22891 37077
rect 22922 37068 22928 37120
rect 22980 37108 22986 37120
rect 24504 37108 24532 37148
rect 26050 37136 26056 37188
rect 26108 37176 26114 37188
rect 26108 37148 27936 37176
rect 26108 37136 26114 37148
rect 22980 37080 24532 37108
rect 22980 37068 22986 37080
rect 24578 37068 24584 37120
rect 24636 37108 24642 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24636 37080 24777 37108
rect 24636 37068 24642 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25501 37111 25559 37117
rect 25501 37108 25513 37111
rect 25188 37080 25513 37108
rect 25188 37068 25194 37080
rect 25501 37077 25513 37080
rect 25547 37077 25559 37111
rect 25501 37071 25559 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27908 37117 27936 37148
rect 28902 37136 28908 37188
rect 28960 37176 28966 37188
rect 35897 37179 35955 37185
rect 35897 37176 35909 37179
rect 28960 37148 35909 37176
rect 28960 37136 28966 37148
rect 35897 37145 35909 37148
rect 35943 37145 35955 37179
rect 37752 37176 37780 37207
rect 35897 37139 35955 37145
rect 36004 37148 37780 37176
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 27893 37111 27951 37117
rect 27893 37077 27905 37111
rect 27939 37077 27951 37111
rect 28994 37108 29000 37120
rect 28955 37080 29000 37108
rect 27893 37071 27951 37077
rect 28994 37068 29000 37080
rect 29052 37068 29058 37120
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29696 37080 29929 37108
rect 29696 37068 29702 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 30466 37108 30472 37120
rect 30427 37080 30472 37108
rect 29917 37071 29975 37077
rect 30466 37068 30472 37080
rect 30524 37068 30530 37120
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35069 37071 35127 37077
rect 35434 37068 35440 37120
rect 35492 37108 35498 37120
rect 36004 37108 36032 37148
rect 35492 37080 36032 37108
rect 35492 37068 35498 37080
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36541 37111 36599 37117
rect 36541 37108 36553 37111
rect 36136 37080 36553 37108
rect 36136 37068 36142 37080
rect 36541 37077 36553 37080
rect 36587 37077 36599 37111
rect 36541 37071 36599 37077
rect 37090 37068 37096 37120
rect 37148 37108 37154 37120
rect 39298 37108 39304 37120
rect 37148 37080 39304 37108
rect 37148 37068 37154 37080
rect 39298 37068 39304 37080
rect 39356 37068 39362 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1302 36864 1308 36916
rect 1360 36904 1366 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 1360 36876 1777 36904
rect 1360 36864 1366 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 2501 36907 2559 36913
rect 2501 36873 2513 36907
rect 2547 36904 2559 36907
rect 2866 36904 2872 36916
rect 2547 36876 2872 36904
rect 2547 36873 2559 36876
rect 2501 36867 2559 36873
rect 2866 36864 2872 36876
rect 2924 36864 2930 36916
rect 3050 36864 3056 36916
rect 3108 36864 3114 36916
rect 3142 36864 3148 36916
rect 3200 36904 3206 36916
rect 3237 36907 3295 36913
rect 3237 36904 3249 36907
rect 3200 36876 3249 36904
rect 3200 36864 3206 36876
rect 3237 36873 3249 36876
rect 3283 36873 3295 36907
rect 3237 36867 3295 36873
rect 6825 36907 6883 36913
rect 6825 36873 6837 36907
rect 6871 36873 6883 36907
rect 10686 36904 10692 36916
rect 6825 36867 6883 36873
rect 7760 36876 10692 36904
rect 3068 36836 3096 36864
rect 5442 36836 5448 36848
rect 3068 36808 5448 36836
rect 5442 36796 5448 36808
rect 5500 36796 5506 36848
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36737 1639 36771
rect 2314 36768 2320 36780
rect 2275 36740 2320 36768
rect 1581 36731 1639 36737
rect 1596 36700 1624 36731
rect 2314 36728 2320 36740
rect 2372 36728 2378 36780
rect 3053 36771 3111 36777
rect 3053 36737 3065 36771
rect 3099 36768 3111 36771
rect 6840 36768 6868 36867
rect 3099 36740 6868 36768
rect 7009 36771 7067 36777
rect 3099 36737 3111 36740
rect 3053 36731 3111 36737
rect 7009 36737 7021 36771
rect 7055 36737 7067 36771
rect 7760 36768 7788 36876
rect 10686 36864 10692 36876
rect 10744 36864 10750 36916
rect 11606 36864 11612 36916
rect 11664 36904 11670 36916
rect 11885 36907 11943 36913
rect 11885 36904 11897 36907
rect 11664 36876 11897 36904
rect 11664 36864 11670 36876
rect 11885 36873 11897 36876
rect 11931 36873 11943 36907
rect 11885 36867 11943 36873
rect 19521 36907 19579 36913
rect 19521 36873 19533 36907
rect 19567 36904 19579 36907
rect 19978 36904 19984 36916
rect 19567 36876 19984 36904
rect 19567 36873 19579 36876
rect 19521 36867 19579 36873
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 20257 36907 20315 36913
rect 20257 36873 20269 36907
rect 20303 36873 20315 36907
rect 22462 36904 22468 36916
rect 22423 36876 22468 36904
rect 20257 36867 20315 36873
rect 7834 36796 7840 36848
rect 7892 36836 7898 36848
rect 20272 36836 20300 36867
rect 22462 36864 22468 36876
rect 22520 36864 22526 36916
rect 24026 36904 24032 36916
rect 23987 36876 24032 36904
rect 24026 36864 24032 36876
rect 24084 36864 24090 36916
rect 32214 36864 32220 36916
rect 32272 36904 32278 36916
rect 32493 36907 32551 36913
rect 32493 36904 32505 36907
rect 32272 36876 32505 36904
rect 32272 36864 32278 36876
rect 32493 36873 32505 36876
rect 32539 36873 32551 36907
rect 32493 36867 32551 36873
rect 36081 36907 36139 36913
rect 36081 36873 36093 36907
rect 36127 36904 36139 36907
rect 36170 36904 36176 36916
rect 36127 36876 36176 36904
rect 36127 36873 36139 36876
rect 36081 36867 36139 36873
rect 36170 36864 36176 36876
rect 36228 36864 36234 36916
rect 36722 36864 36728 36916
rect 36780 36864 36786 36916
rect 28902 36836 28908 36848
rect 7892 36808 20300 36836
rect 20456 36808 28908 36836
rect 7892 36796 7898 36808
rect 8113 36771 8171 36777
rect 8113 36768 8125 36771
rect 7760 36740 8125 36768
rect 7009 36731 7067 36737
rect 8113 36737 8125 36740
rect 8159 36737 8171 36771
rect 8113 36731 8171 36737
rect 2406 36700 2412 36712
rect 1596 36672 2412 36700
rect 2406 36660 2412 36672
rect 2464 36660 2470 36712
rect 3970 36660 3976 36712
rect 4028 36700 4034 36712
rect 6914 36700 6920 36712
rect 4028 36672 6920 36700
rect 4028 36660 4034 36672
rect 6914 36660 6920 36672
rect 6972 36660 6978 36712
rect 7024 36700 7052 36731
rect 9030 36728 9036 36780
rect 9088 36768 9094 36780
rect 9309 36771 9367 36777
rect 9309 36768 9321 36771
rect 9088 36740 9321 36768
rect 9088 36728 9094 36740
rect 9309 36737 9321 36740
rect 9355 36737 9367 36771
rect 9309 36731 9367 36737
rect 10318 36728 10324 36780
rect 10376 36768 10382 36780
rect 11701 36771 11759 36777
rect 11701 36768 11713 36771
rect 10376 36740 11713 36768
rect 10376 36728 10382 36740
rect 11701 36737 11713 36740
rect 11747 36737 11759 36771
rect 11701 36731 11759 36737
rect 14182 36728 14188 36780
rect 14240 36768 14246 36780
rect 14277 36771 14335 36777
rect 14277 36768 14289 36771
rect 14240 36740 14289 36768
rect 14240 36728 14246 36740
rect 14277 36737 14289 36740
rect 14323 36737 14335 36771
rect 14277 36731 14335 36737
rect 16758 36728 16764 36780
rect 16816 36768 16822 36780
rect 17037 36771 17095 36777
rect 17037 36768 17049 36771
rect 16816 36740 17049 36768
rect 16816 36728 16822 36740
rect 17037 36737 17049 36740
rect 17083 36737 17095 36771
rect 18874 36768 18880 36780
rect 18835 36740 18880 36768
rect 17037 36731 17095 36737
rect 18874 36728 18880 36740
rect 18932 36728 18938 36780
rect 20456 36777 20484 36808
rect 28902 36796 28908 36808
rect 28960 36796 28966 36848
rect 30282 36796 30288 36848
rect 30340 36836 30346 36848
rect 36740 36836 36768 36864
rect 37553 36839 37611 36845
rect 37553 36836 37565 36839
rect 30340 36808 35112 36836
rect 36740 36808 37565 36836
rect 30340 36796 30346 36808
rect 18969 36771 19027 36777
rect 18969 36737 18981 36771
rect 19015 36768 19027 36771
rect 19705 36771 19763 36777
rect 19705 36768 19717 36771
rect 19015 36740 19717 36768
rect 19015 36737 19027 36740
rect 18969 36731 19027 36737
rect 19705 36737 19717 36740
rect 19751 36737 19763 36771
rect 19705 36731 19763 36737
rect 20441 36771 20499 36777
rect 20441 36737 20453 36771
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 22649 36771 22707 36777
rect 22649 36737 22661 36771
rect 22695 36737 22707 36771
rect 23566 36768 23572 36780
rect 23527 36740 23572 36768
rect 22649 36731 22707 36737
rect 12894 36700 12900 36712
rect 7024 36672 12900 36700
rect 12894 36660 12900 36672
rect 12952 36700 12958 36712
rect 14553 36703 14611 36709
rect 14553 36700 14565 36703
rect 12952 36672 14565 36700
rect 12952 36660 12958 36672
rect 14553 36669 14565 36672
rect 14599 36669 14611 36703
rect 22664 36700 22692 36731
rect 23566 36728 23572 36740
rect 23624 36728 23630 36780
rect 24210 36768 24216 36780
rect 24171 36740 24216 36768
rect 24210 36728 24216 36740
rect 24268 36728 24274 36780
rect 35084 36777 35112 36808
rect 37553 36805 37565 36808
rect 37599 36805 37611 36839
rect 37553 36799 37611 36805
rect 32309 36771 32367 36777
rect 32309 36737 32321 36771
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 35069 36771 35127 36777
rect 35069 36737 35081 36771
rect 35115 36737 35127 36771
rect 35069 36731 35127 36737
rect 23014 36700 23020 36712
rect 22664 36672 23020 36700
rect 14553 36663 14611 36669
rect 23014 36660 23020 36672
rect 23072 36700 23078 36712
rect 30742 36700 30748 36712
rect 23072 36672 30748 36700
rect 23072 36660 23078 36672
rect 30742 36660 30748 36672
rect 30800 36660 30806 36712
rect 5074 36592 5080 36644
rect 5132 36632 5138 36644
rect 7929 36635 7987 36641
rect 7929 36632 7941 36635
rect 5132 36604 7941 36632
rect 5132 36592 5138 36604
rect 7929 36601 7941 36604
rect 7975 36601 7987 36635
rect 7929 36595 7987 36601
rect 23385 36635 23443 36641
rect 23385 36601 23397 36635
rect 23431 36632 23443 36635
rect 32324 36632 32352 36731
rect 35526 36728 35532 36780
rect 35584 36768 35590 36780
rect 35897 36771 35955 36777
rect 35897 36768 35909 36771
rect 35584 36740 35909 36768
rect 35584 36728 35590 36740
rect 35897 36737 35909 36740
rect 35943 36737 35955 36771
rect 35897 36731 35955 36737
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36768 36783 36771
rect 36814 36768 36820 36780
rect 36771 36740 36820 36768
rect 36771 36737 36783 36740
rect 36725 36731 36783 36737
rect 36814 36728 36820 36740
rect 36872 36728 36878 36780
rect 23431 36604 32352 36632
rect 35161 36635 35219 36641
rect 23431 36601 23443 36604
rect 23385 36595 23443 36601
rect 35161 36601 35173 36635
rect 35207 36632 35219 36635
rect 37366 36632 37372 36644
rect 35207 36604 37372 36632
rect 35207 36601 35219 36604
rect 35161 36595 35219 36601
rect 37366 36592 37372 36604
rect 37424 36592 37430 36644
rect 5350 36524 5356 36576
rect 5408 36564 5414 36576
rect 9030 36564 9036 36576
rect 5408 36536 9036 36564
rect 5408 36524 5414 36536
rect 9030 36524 9036 36536
rect 9088 36524 9094 36576
rect 9125 36567 9183 36573
rect 9125 36533 9137 36567
rect 9171 36564 9183 36567
rect 9398 36564 9404 36576
rect 9171 36536 9404 36564
rect 9171 36533 9183 36536
rect 9125 36527 9183 36533
rect 9398 36524 9404 36536
rect 9456 36524 9462 36576
rect 16853 36567 16911 36573
rect 16853 36533 16865 36567
rect 16899 36564 16911 36567
rect 17034 36564 17040 36576
rect 16899 36536 17040 36564
rect 16899 36533 16911 36536
rect 16853 36527 16911 36533
rect 17034 36524 17040 36536
rect 17092 36524 17098 36576
rect 35526 36564 35532 36576
rect 35487 36536 35532 36564
rect 35526 36524 35532 36536
rect 35584 36524 35590 36576
rect 36814 36564 36820 36576
rect 36775 36536 36820 36564
rect 36814 36524 36820 36536
rect 36872 36524 36878 36576
rect 37642 36564 37648 36576
rect 37603 36536 37648 36564
rect 37642 36524 37648 36536
rect 37700 36524 37706 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 658 36320 664 36372
rect 716 36360 722 36372
rect 2501 36363 2559 36369
rect 2501 36360 2513 36363
rect 716 36332 2513 36360
rect 716 36320 722 36332
rect 2501 36329 2513 36332
rect 2547 36329 2559 36363
rect 2501 36323 2559 36329
rect 15746 36320 15752 36372
rect 15804 36360 15810 36372
rect 23566 36360 23572 36372
rect 15804 36332 23572 36360
rect 15804 36320 15810 36332
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 36725 36363 36783 36369
rect 36725 36329 36737 36363
rect 36771 36360 36783 36363
rect 38654 36360 38660 36372
rect 36771 36332 38660 36360
rect 36771 36329 36783 36332
rect 36725 36323 36783 36329
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 23474 36252 23480 36304
rect 23532 36292 23538 36304
rect 36814 36292 36820 36304
rect 23532 36264 36820 36292
rect 23532 36252 23538 36264
rect 36814 36252 36820 36264
rect 36872 36252 36878 36304
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 2317 36159 2375 36165
rect 2317 36125 2329 36159
rect 2363 36156 2375 36159
rect 2682 36156 2688 36168
rect 2363 36128 2688 36156
rect 2363 36125 2375 36128
rect 2317 36119 2375 36125
rect 2682 36116 2688 36128
rect 2740 36116 2746 36168
rect 2958 36116 2964 36168
rect 3016 36156 3022 36168
rect 3237 36159 3295 36165
rect 3237 36156 3249 36159
rect 3016 36128 3249 36156
rect 3016 36116 3022 36128
rect 3237 36125 3249 36128
rect 3283 36125 3295 36159
rect 3237 36119 3295 36125
rect 7098 36116 7104 36168
rect 7156 36156 7162 36168
rect 7377 36159 7435 36165
rect 7377 36156 7389 36159
rect 7156 36128 7389 36156
rect 7156 36116 7162 36128
rect 7377 36125 7389 36128
rect 7423 36125 7435 36159
rect 36538 36156 36544 36168
rect 36499 36128 36544 36156
rect 7377 36119 7435 36125
rect 36538 36116 36544 36128
rect 36596 36116 36602 36168
rect 37182 36116 37188 36168
rect 37240 36156 37246 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37240 36128 38025 36156
rect 37240 36116 37246 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 1857 36091 1915 36097
rect 1857 36057 1869 36091
rect 1903 36088 1915 36091
rect 2222 36088 2228 36100
rect 1903 36060 2228 36088
rect 1903 36057 1915 36060
rect 1857 36051 1915 36057
rect 2222 36048 2228 36060
rect 2280 36048 2286 36100
rect 5442 36048 5448 36100
rect 5500 36088 5506 36100
rect 16114 36088 16120 36100
rect 5500 36060 16120 36088
rect 5500 36048 5506 36060
rect 16114 36048 16120 36060
rect 16172 36048 16178 36100
rect 37090 36048 37096 36100
rect 37148 36088 37154 36100
rect 37369 36091 37427 36097
rect 37369 36088 37381 36091
rect 37148 36060 37381 36088
rect 37148 36048 37154 36060
rect 37369 36057 37381 36060
rect 37415 36057 37427 36091
rect 37550 36088 37556 36100
rect 37511 36060 37556 36088
rect 37369 36051 37427 36057
rect 37550 36048 37556 36060
rect 37608 36048 37614 36100
rect 3053 36023 3111 36029
rect 3053 35989 3065 36023
rect 3099 36020 3111 36023
rect 5810 36020 5816 36032
rect 3099 35992 5816 36020
rect 3099 35989 3111 35992
rect 3053 35983 3111 35989
rect 5810 35980 5816 35992
rect 5868 35980 5874 36032
rect 6454 35980 6460 36032
rect 6512 36020 6518 36032
rect 7193 36023 7251 36029
rect 7193 36020 7205 36023
rect 6512 35992 7205 36020
rect 6512 35980 6518 35992
rect 7193 35989 7205 35992
rect 7239 35989 7251 36023
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 7193 35983 7251 35989
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 2314 35816 2320 35828
rect 2275 35788 2320 35816
rect 2314 35776 2320 35788
rect 2372 35776 2378 35828
rect 23385 35819 23443 35825
rect 23385 35785 23397 35819
rect 23431 35816 23443 35819
rect 24210 35816 24216 35828
rect 23431 35788 24216 35816
rect 23431 35785 23443 35788
rect 23385 35779 23443 35785
rect 24210 35776 24216 35788
rect 24268 35776 24274 35828
rect 38197 35819 38255 35825
rect 38197 35785 38209 35819
rect 38243 35816 38255 35819
rect 38286 35816 38292 35828
rect 38243 35788 38292 35816
rect 38243 35785 38255 35788
rect 38197 35779 38255 35785
rect 38286 35776 38292 35788
rect 38344 35776 38350 35828
rect 1596 35720 6914 35748
rect 1596 35689 1624 35720
rect 1581 35683 1639 35689
rect 1581 35649 1593 35683
rect 1627 35649 1639 35683
rect 1581 35643 1639 35649
rect 1854 35640 1860 35692
rect 1912 35680 1918 35692
rect 2501 35683 2559 35689
rect 2501 35680 2513 35683
rect 1912 35652 2513 35680
rect 1912 35640 1918 35652
rect 2501 35649 2513 35652
rect 2547 35649 2559 35683
rect 2501 35643 2559 35649
rect 6886 35544 6914 35720
rect 20346 35708 20352 35760
rect 20404 35748 20410 35760
rect 20404 35720 23336 35748
rect 20404 35708 20410 35720
rect 23308 35689 23336 35720
rect 22189 35683 22247 35689
rect 22189 35649 22201 35683
rect 22235 35649 22247 35683
rect 22189 35643 22247 35649
rect 23293 35683 23351 35689
rect 23293 35649 23305 35683
rect 23339 35649 23351 35683
rect 23293 35643 23351 35649
rect 22204 35612 22232 35643
rect 36722 35640 36728 35692
rect 36780 35680 36786 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 36780 35652 38025 35680
rect 36780 35640 36786 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 23474 35612 23480 35624
rect 22204 35584 23480 35612
rect 23474 35572 23480 35584
rect 23532 35572 23538 35624
rect 22005 35547 22063 35553
rect 22005 35544 22017 35547
rect 6886 35516 22017 35544
rect 22005 35513 22017 35516
rect 22051 35513 22063 35547
rect 22005 35507 22063 35513
rect 1762 35476 1768 35488
rect 1723 35448 1768 35476
rect 1762 35436 1768 35448
rect 1820 35436 1826 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 37182 35272 37188 35284
rect 37143 35244 37188 35272
rect 37182 35232 37188 35244
rect 37240 35232 37246 35284
rect 37366 35068 37372 35080
rect 37327 35040 37372 35068
rect 37366 35028 37372 35040
rect 37424 35028 37430 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 37660 35040 38025 35068
rect 37458 34892 37464 34944
rect 37516 34932 37522 34944
rect 37660 34941 37688 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 37645 34935 37703 34941
rect 37645 34932 37657 34935
rect 37516 34904 37657 34932
rect 37516 34892 37522 34904
rect 37645 34901 37657 34904
rect 37691 34901 37703 34935
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 37645 34895 37703 34901
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 2590 34728 2596 34740
rect 1627 34700 2596 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 2590 34688 2596 34700
rect 2648 34688 2654 34740
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 31754 34552 31760 34604
rect 31812 34592 31818 34604
rect 37737 34595 37795 34601
rect 37737 34592 37749 34595
rect 31812 34564 37749 34592
rect 31812 34552 31818 34564
rect 37737 34561 37749 34564
rect 37783 34561 37795 34595
rect 37737 34555 37795 34561
rect 37182 34484 37188 34536
rect 37240 34524 37246 34536
rect 37461 34527 37519 34533
rect 37461 34524 37473 34527
rect 37240 34496 37473 34524
rect 37240 34484 37246 34496
rect 37461 34493 37473 34496
rect 37507 34493 37519 34527
rect 37461 34487 37519 34493
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 17126 33804 17132 33856
rect 17184 33844 17190 33856
rect 33594 33844 33600 33856
rect 17184 33816 33600 33844
rect 17184 33804 17190 33816
rect 33594 33804 33600 33816
rect 33652 33804 33658 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 35805 33643 35863 33649
rect 35805 33609 35817 33643
rect 35851 33640 35863 33643
rect 36722 33640 36728 33652
rect 35851 33612 36728 33640
rect 35851 33609 35863 33612
rect 35805 33603 35863 33609
rect 36722 33600 36728 33612
rect 36780 33600 36786 33652
rect 1581 33507 1639 33513
rect 1581 33473 1593 33507
rect 1627 33504 1639 33507
rect 4614 33504 4620 33516
rect 1627 33476 4620 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 4614 33464 4620 33476
rect 4672 33464 4678 33516
rect 5810 33504 5816 33516
rect 5771 33476 5816 33504
rect 5810 33464 5816 33476
rect 5868 33464 5874 33516
rect 27341 33507 27399 33513
rect 27341 33504 27353 33507
rect 26206 33476 27353 33504
rect 2038 33396 2044 33448
rect 2096 33436 2102 33448
rect 26206 33436 26234 33476
rect 27341 33473 27353 33476
rect 27387 33504 27399 33507
rect 27617 33507 27675 33513
rect 27617 33504 27629 33507
rect 27387 33476 27629 33504
rect 27387 33473 27399 33476
rect 27341 33467 27399 33473
rect 27617 33473 27629 33476
rect 27663 33473 27675 33507
rect 27617 33467 27675 33473
rect 34606 33464 34612 33516
rect 34664 33504 34670 33516
rect 35989 33507 36047 33513
rect 35989 33504 36001 33507
rect 34664 33476 36001 33504
rect 34664 33464 34670 33476
rect 35989 33473 36001 33476
rect 36035 33473 36047 33507
rect 35989 33467 36047 33473
rect 38013 33507 38071 33513
rect 38013 33473 38025 33507
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 2096 33408 26234 33436
rect 2096 33396 2102 33408
rect 1762 33368 1768 33380
rect 1723 33340 1768 33368
rect 1762 33328 1768 33340
rect 1820 33328 1826 33380
rect 27157 33371 27215 33377
rect 27157 33337 27169 33371
rect 27203 33368 27215 33371
rect 38028 33368 38056 33467
rect 38194 33368 38200 33380
rect 27203 33340 38056 33368
rect 38155 33340 38200 33368
rect 27203 33337 27215 33340
rect 27157 33331 27215 33337
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 5905 33303 5963 33309
rect 5905 33269 5917 33303
rect 5951 33300 5963 33303
rect 8938 33300 8944 33312
rect 5951 33272 8944 33300
rect 5951 33269 5963 33272
rect 5905 33263 5963 33269
rect 8938 33260 8944 33272
rect 8996 33260 9002 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 26050 32892 26056 32904
rect 26011 32864 26056 32892
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 19334 32716 19340 32768
rect 19392 32756 19398 32768
rect 19429 32759 19487 32765
rect 19429 32756 19441 32759
rect 19392 32728 19441 32756
rect 19392 32716 19398 32728
rect 19429 32725 19441 32728
rect 19475 32725 19487 32759
rect 19429 32719 19487 32725
rect 25222 32716 25228 32768
rect 25280 32756 25286 32768
rect 26145 32759 26203 32765
rect 26145 32756 26157 32759
rect 25280 32728 26157 32756
rect 25280 32716 25286 32728
rect 26145 32725 26157 32728
rect 26191 32725 26203 32759
rect 26145 32719 26203 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 2682 32512 2688 32564
rect 2740 32552 2746 32564
rect 33318 32552 33324 32564
rect 2740 32524 33324 32552
rect 2740 32512 2746 32524
rect 33318 32512 33324 32524
rect 33376 32512 33382 32564
rect 19334 32484 19340 32496
rect 19295 32456 19340 32484
rect 19334 32444 19340 32456
rect 19392 32444 19398 32496
rect 19429 32487 19487 32493
rect 19429 32453 19441 32487
rect 19475 32484 19487 32487
rect 19978 32484 19984 32496
rect 19475 32456 19984 32484
rect 19475 32453 19487 32456
rect 19429 32447 19487 32453
rect 19978 32444 19984 32456
rect 20036 32444 20042 32496
rect 20346 32484 20352 32496
rect 20307 32456 20352 32484
rect 20346 32444 20352 32456
rect 20404 32444 20410 32496
rect 28994 32376 29000 32428
rect 29052 32416 29058 32428
rect 30653 32419 30711 32425
rect 30653 32416 30665 32419
rect 29052 32388 30665 32416
rect 29052 32376 29058 32388
rect 30653 32385 30665 32388
rect 30699 32385 30711 32419
rect 30653 32379 30711 32385
rect 33134 32376 33140 32428
rect 33192 32416 33198 32428
rect 37737 32419 37795 32425
rect 37737 32416 37749 32419
rect 33192 32388 37749 32416
rect 33192 32376 33198 32388
rect 37737 32385 37749 32388
rect 37783 32385 37795 32419
rect 37737 32379 37795 32385
rect 1578 32348 1584 32360
rect 1539 32320 1584 32348
rect 1578 32308 1584 32320
rect 1636 32308 1642 32360
rect 1854 32348 1860 32360
rect 1815 32320 1860 32348
rect 1854 32308 1860 32320
rect 1912 32308 1918 32360
rect 37458 32348 37464 32360
rect 37419 32320 37464 32348
rect 37458 32308 37464 32320
rect 37516 32308 37522 32360
rect 30742 32212 30748 32224
rect 30703 32184 30748 32212
rect 30742 32172 30748 32184
rect 30800 32172 30806 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 9122 31900 9128 31952
rect 9180 31940 9186 31952
rect 9217 31943 9275 31949
rect 9217 31940 9229 31943
rect 9180 31912 9229 31940
rect 9180 31900 9186 31912
rect 9217 31909 9229 31912
rect 9263 31909 9275 31943
rect 9217 31903 9275 31909
rect 12621 31943 12679 31949
rect 12621 31909 12633 31943
rect 12667 31940 12679 31943
rect 14458 31940 14464 31952
rect 12667 31912 14464 31940
rect 12667 31909 12679 31912
rect 12621 31903 12679 31909
rect 14458 31900 14464 31912
rect 14516 31900 14522 31952
rect 38194 31940 38200 31952
rect 38155 31912 38200 31940
rect 38194 31900 38200 31912
rect 38252 31900 38258 31952
rect 6454 31872 6460 31884
rect 5736 31844 6460 31872
rect 1581 31807 1639 31813
rect 1581 31773 1593 31807
rect 1627 31804 1639 31807
rect 1670 31804 1676 31816
rect 1627 31776 1676 31804
rect 1627 31773 1639 31776
rect 1581 31767 1639 31773
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 5736 31813 5764 31844
rect 6454 31832 6460 31844
rect 6512 31832 6518 31884
rect 10962 31832 10968 31884
rect 11020 31872 11026 31884
rect 11020 31844 13216 31872
rect 11020 31832 11026 31844
rect 5721 31807 5779 31813
rect 5721 31773 5733 31807
rect 5767 31773 5779 31807
rect 5721 31767 5779 31773
rect 5813 31807 5871 31813
rect 5813 31773 5825 31807
rect 5859 31804 5871 31807
rect 6086 31804 6092 31816
rect 5859 31776 6092 31804
rect 5859 31773 5871 31776
rect 5813 31767 5871 31773
rect 6086 31764 6092 31776
rect 6144 31764 6150 31816
rect 9030 31764 9036 31816
rect 9088 31804 9094 31816
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 9088 31776 9137 31804
rect 9088 31764 9094 31776
rect 9125 31773 9137 31776
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 9398 31764 9404 31816
rect 9456 31804 9462 31816
rect 13188 31813 13216 31844
rect 12529 31807 12587 31813
rect 12529 31804 12541 31807
rect 9456 31776 12541 31804
rect 9456 31764 9462 31776
rect 12529 31773 12541 31776
rect 12575 31773 12587 31807
rect 12529 31767 12587 31773
rect 13173 31807 13231 31813
rect 13173 31773 13185 31807
rect 13219 31773 13231 31807
rect 13173 31767 13231 31773
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31804 13323 31807
rect 14734 31804 14740 31816
rect 13311 31776 14740 31804
rect 13311 31773 13323 31776
rect 13265 31767 13323 31773
rect 14734 31764 14740 31776
rect 14792 31764 14798 31816
rect 38010 31804 38016 31816
rect 37971 31776 38016 31804
rect 38010 31764 38016 31776
rect 38068 31764 38074 31816
rect 1762 31668 1768 31680
rect 1723 31640 1768 31668
rect 1762 31628 1768 31640
rect 1820 31628 1826 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 38010 31424 38016 31476
rect 38068 31464 38074 31476
rect 38105 31467 38163 31473
rect 38105 31464 38117 31467
rect 38068 31436 38117 31464
rect 38068 31424 38074 31436
rect 38105 31433 38117 31436
rect 38151 31433 38163 31467
rect 38105 31427 38163 31433
rect 17126 31396 17132 31408
rect 17087 31368 17132 31396
rect 17126 31356 17132 31368
rect 17184 31356 17190 31408
rect 6914 31288 6920 31340
rect 6972 31328 6978 31340
rect 7561 31331 7619 31337
rect 7561 31328 7573 31331
rect 6972 31300 7573 31328
rect 6972 31288 6978 31300
rect 7561 31297 7573 31300
rect 7607 31297 7619 31331
rect 7561 31291 7619 31297
rect 13814 31288 13820 31340
rect 13872 31328 13878 31340
rect 14645 31331 14703 31337
rect 14645 31328 14657 31331
rect 13872 31300 14657 31328
rect 13872 31288 13878 31300
rect 14645 31297 14657 31300
rect 14691 31297 14703 31331
rect 14645 31291 14703 31297
rect 16574 31288 16580 31340
rect 16632 31328 16638 31340
rect 16945 31331 17003 31337
rect 16945 31328 16957 31331
rect 16632 31300 16957 31328
rect 16632 31288 16638 31300
rect 16945 31297 16957 31300
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 25501 31331 25559 31337
rect 25501 31297 25513 31331
rect 25547 31328 25559 31331
rect 30466 31328 30472 31340
rect 25547 31300 30472 31328
rect 25547 31297 25559 31300
rect 25501 31291 25559 31297
rect 30466 31288 30472 31300
rect 30524 31288 30530 31340
rect 35434 31288 35440 31340
rect 35492 31328 35498 31340
rect 37461 31331 37519 31337
rect 37461 31328 37473 31331
rect 35492 31300 37473 31328
rect 35492 31288 35498 31300
rect 37461 31297 37473 31300
rect 37507 31297 37519 31331
rect 37461 31291 37519 31297
rect 37553 31331 37611 31337
rect 37553 31297 37565 31331
rect 37599 31328 37611 31331
rect 38289 31331 38347 31337
rect 38289 31328 38301 31331
rect 37599 31300 38301 31328
rect 37599 31297 37611 31300
rect 37553 31291 37611 31297
rect 38289 31297 38301 31300
rect 38335 31297 38347 31331
rect 38289 31291 38347 31297
rect 14458 31260 14464 31272
rect 14419 31232 14464 31260
rect 14458 31220 14464 31232
rect 14516 31220 14522 31272
rect 14826 31220 14832 31272
rect 14884 31260 14890 31272
rect 15565 31263 15623 31269
rect 15565 31260 15577 31263
rect 14884 31232 15577 31260
rect 14884 31220 14890 31232
rect 15565 31229 15577 31232
rect 15611 31229 15623 31263
rect 15565 31223 15623 31229
rect 7374 31084 7380 31136
rect 7432 31124 7438 31136
rect 7653 31127 7711 31133
rect 7653 31124 7665 31127
rect 7432 31096 7665 31124
rect 7432 31084 7438 31096
rect 7653 31093 7665 31096
rect 7699 31093 7711 31127
rect 14918 31124 14924 31136
rect 14879 31096 14924 31124
rect 7653 31087 7711 31093
rect 14918 31084 14924 31096
rect 14976 31084 14982 31136
rect 22094 31084 22100 31136
rect 22152 31124 22158 31136
rect 25593 31127 25651 31133
rect 25593 31124 25605 31127
rect 22152 31096 25605 31124
rect 22152 31084 22158 31096
rect 25593 31093 25605 31096
rect 25639 31093 25651 31127
rect 25593 31087 25651 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 4249 30923 4307 30929
rect 4249 30889 4261 30923
rect 4295 30920 4307 30923
rect 4614 30920 4620 30932
rect 4295 30892 4620 30920
rect 4295 30889 4307 30892
rect 4249 30883 4307 30889
rect 4614 30880 4620 30892
rect 4672 30880 4678 30932
rect 12986 30920 12992 30932
rect 12947 30892 12992 30920
rect 12986 30880 12992 30892
rect 13044 30880 13050 30932
rect 21174 30880 21180 30932
rect 21232 30920 21238 30932
rect 22649 30923 22707 30929
rect 22649 30920 22661 30923
rect 21232 30892 22661 30920
rect 21232 30880 21238 30892
rect 22649 30889 22661 30892
rect 22695 30889 22707 30923
rect 22649 30883 22707 30889
rect 14918 30812 14924 30864
rect 14976 30852 14982 30864
rect 15197 30855 15255 30861
rect 15197 30852 15209 30855
rect 14976 30824 15209 30852
rect 14976 30812 14982 30824
rect 15197 30821 15209 30824
rect 15243 30821 15255 30855
rect 15197 30815 15255 30821
rect 8938 30744 8944 30796
rect 8996 30784 9002 30796
rect 10965 30787 11023 30793
rect 10965 30784 10977 30787
rect 8996 30756 10977 30784
rect 8996 30744 9002 30756
rect 10965 30753 10977 30756
rect 11011 30753 11023 30787
rect 10965 30747 11023 30753
rect 11977 30787 12035 30793
rect 11977 30753 11989 30787
rect 12023 30784 12035 30787
rect 12802 30784 12808 30796
rect 12023 30756 12808 30784
rect 12023 30753 12035 30756
rect 11977 30747 12035 30753
rect 12802 30744 12808 30756
rect 12860 30744 12866 30796
rect 14826 30784 14832 30796
rect 14787 30756 14832 30784
rect 14826 30744 14832 30756
rect 14884 30744 14890 30796
rect 1762 30716 1768 30728
rect 1723 30688 1768 30716
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 4433 30719 4491 30725
rect 4433 30685 4445 30719
rect 4479 30716 4491 30719
rect 10686 30716 10692 30728
rect 4479 30688 10692 30716
rect 4479 30685 4491 30688
rect 4433 30679 4491 30685
rect 10686 30676 10692 30688
rect 10744 30676 10750 30728
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 12406 30688 13185 30716
rect 11054 30608 11060 30660
rect 11112 30648 11118 30660
rect 11112 30620 11157 30648
rect 11112 30608 11118 30620
rect 11606 30608 11612 30660
rect 11664 30648 11670 30660
rect 12406 30648 12434 30688
rect 13173 30685 13185 30688
rect 13219 30685 13231 30719
rect 13173 30679 13231 30685
rect 15013 30719 15071 30725
rect 15013 30685 15025 30719
rect 15059 30716 15071 30719
rect 15378 30716 15384 30728
rect 15059 30688 15384 30716
rect 15059 30685 15071 30688
rect 15013 30679 15071 30685
rect 15378 30676 15384 30688
rect 15436 30676 15442 30728
rect 22833 30719 22891 30725
rect 22833 30685 22845 30719
rect 22879 30685 22891 30719
rect 22833 30679 22891 30685
rect 11664 30620 12434 30648
rect 22848 30648 22876 30679
rect 24394 30676 24400 30728
rect 24452 30716 24458 30728
rect 24581 30719 24639 30725
rect 24581 30716 24593 30719
rect 24452 30688 24593 30716
rect 24452 30676 24458 30688
rect 24581 30685 24593 30688
rect 24627 30685 24639 30719
rect 24581 30679 24639 30685
rect 25590 30648 25596 30660
rect 22848 30620 25596 30648
rect 11664 30608 11670 30620
rect 25590 30608 25596 30620
rect 25648 30608 25654 30660
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 6730 30580 6736 30592
rect 1627 30552 6736 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 24673 30583 24731 30589
rect 24673 30549 24685 30583
rect 24719 30580 24731 30583
rect 29086 30580 29092 30592
rect 24719 30552 29092 30580
rect 24719 30549 24731 30552
rect 24673 30543 24731 30549
rect 29086 30540 29092 30552
rect 29144 30540 29150 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 11054 30336 11060 30388
rect 11112 30376 11118 30388
rect 12161 30379 12219 30385
rect 12161 30376 12173 30379
rect 11112 30348 12173 30376
rect 11112 30336 11118 30348
rect 12161 30345 12173 30348
rect 12207 30345 12219 30379
rect 12161 30339 12219 30345
rect 21818 30336 21824 30388
rect 21876 30376 21882 30388
rect 21876 30348 24256 30376
rect 21876 30336 21882 30348
rect 13173 30311 13231 30317
rect 13173 30277 13185 30311
rect 13219 30308 13231 30311
rect 13814 30308 13820 30320
rect 13219 30280 13820 30308
rect 13219 30277 13231 30280
rect 13173 30271 13231 30277
rect 13814 30268 13820 30280
rect 13872 30268 13878 30320
rect 14458 30308 14464 30320
rect 14419 30280 14464 30308
rect 14458 30268 14464 30280
rect 14516 30268 14522 30320
rect 14553 30311 14611 30317
rect 14553 30277 14565 30311
rect 14599 30308 14611 30311
rect 16022 30308 16028 30320
rect 14599 30280 16028 30308
rect 14599 30277 14611 30280
rect 14553 30271 14611 30277
rect 16022 30268 16028 30280
rect 16080 30268 16086 30320
rect 16209 30311 16267 30317
rect 16209 30277 16221 30311
rect 16255 30308 16267 30311
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 16255 30280 17049 30308
rect 16255 30277 16267 30280
rect 16209 30271 16267 30277
rect 17037 30277 17049 30280
rect 17083 30277 17095 30311
rect 17037 30271 17095 30277
rect 17589 30311 17647 30317
rect 17589 30277 17601 30311
rect 17635 30308 17647 30311
rect 18874 30308 18880 30320
rect 17635 30280 18880 30308
rect 17635 30277 17647 30280
rect 17589 30271 17647 30277
rect 12069 30243 12127 30249
rect 12069 30209 12081 30243
rect 12115 30209 12127 30243
rect 12069 30203 12127 30209
rect 12084 30172 12112 30203
rect 12158 30200 12164 30252
rect 12216 30240 12222 30252
rect 13081 30243 13139 30249
rect 13081 30240 13093 30243
rect 12216 30212 13093 30240
rect 12216 30200 12222 30212
rect 13081 30209 13093 30212
rect 13127 30240 13139 30243
rect 13725 30243 13783 30249
rect 13725 30240 13737 30243
rect 13127 30212 13737 30240
rect 13127 30209 13139 30212
rect 13081 30203 13139 30209
rect 13725 30209 13737 30212
rect 13771 30209 13783 30243
rect 16114 30240 16120 30252
rect 13725 30203 13783 30209
rect 15396 30212 15700 30240
rect 16075 30212 16120 30240
rect 15102 30172 15108 30184
rect 12084 30144 15108 30172
rect 15102 30132 15108 30144
rect 15160 30132 15166 30184
rect 14918 30064 14924 30116
rect 14976 30104 14982 30116
rect 15396 30104 15424 30212
rect 15473 30175 15531 30181
rect 15473 30141 15485 30175
rect 15519 30141 15531 30175
rect 15672 30172 15700 30212
rect 16114 30200 16120 30212
rect 16172 30200 16178 30252
rect 16945 30175 17003 30181
rect 16945 30172 16957 30175
rect 15672 30144 16957 30172
rect 15473 30135 15531 30141
rect 16945 30141 16957 30144
rect 16991 30141 17003 30175
rect 16945 30135 17003 30141
rect 14976 30076 15424 30104
rect 14976 30064 14982 30076
rect 13817 30039 13875 30045
rect 13817 30005 13829 30039
rect 13863 30036 13875 30039
rect 15010 30036 15016 30048
rect 13863 30008 15016 30036
rect 13863 30005 13875 30008
rect 13817 29999 13875 30005
rect 15010 29996 15016 30008
rect 15068 29996 15074 30048
rect 15488 30036 15516 30135
rect 16298 30064 16304 30116
rect 16356 30104 16362 30116
rect 17604 30104 17632 30271
rect 18874 30268 18880 30280
rect 18932 30268 18938 30320
rect 21910 30268 21916 30320
rect 21968 30308 21974 30320
rect 22189 30311 22247 30317
rect 22189 30308 22201 30311
rect 21968 30280 22201 30308
rect 21968 30268 21974 30280
rect 22189 30277 22201 30280
rect 22235 30277 22247 30311
rect 22189 30271 22247 30277
rect 24228 30308 24256 30348
rect 26694 30308 26700 30320
rect 24228 30280 26700 30308
rect 23474 30200 23480 30252
rect 23532 30240 23538 30252
rect 24228 30249 24256 30280
rect 26694 30268 26700 30280
rect 26752 30268 26758 30320
rect 26786 30268 26792 30320
rect 26844 30308 26850 30320
rect 29181 30311 29239 30317
rect 29181 30308 29193 30311
rect 26844 30280 29193 30308
rect 26844 30268 26850 30280
rect 29181 30277 29193 30280
rect 29227 30277 29239 30311
rect 29181 30271 29239 30277
rect 23569 30243 23627 30249
rect 23569 30240 23581 30243
rect 23532 30212 23581 30240
rect 23532 30200 23538 30212
rect 23569 30209 23581 30212
rect 23615 30209 23627 30243
rect 23569 30203 23627 30209
rect 24213 30243 24271 30249
rect 24213 30209 24225 30243
rect 24259 30209 24271 30243
rect 24213 30203 24271 30209
rect 25133 30243 25191 30249
rect 25133 30209 25145 30243
rect 25179 30240 25191 30243
rect 26329 30243 26387 30249
rect 26329 30240 26341 30243
rect 25179 30212 26341 30240
rect 25179 30209 25191 30212
rect 25133 30203 25191 30209
rect 26329 30209 26341 30212
rect 26375 30209 26387 30243
rect 38102 30240 38108 30252
rect 38063 30212 38108 30240
rect 26329 30203 26387 30209
rect 22094 30132 22100 30184
rect 22152 30172 22158 30184
rect 23106 30172 23112 30184
rect 22152 30144 22197 30172
rect 23019 30144 23112 30172
rect 22152 30132 22158 30144
rect 23106 30132 23112 30144
rect 23164 30172 23170 30184
rect 25498 30172 25504 30184
rect 23164 30144 25504 30172
rect 23164 30132 23170 30144
rect 25498 30132 25504 30144
rect 25556 30132 25562 30184
rect 16356 30076 17632 30104
rect 26344 30104 26372 30203
rect 38102 30200 38108 30212
rect 38160 30200 38166 30252
rect 29086 30172 29092 30184
rect 29047 30144 29092 30172
rect 29086 30132 29092 30144
rect 29144 30132 29150 30184
rect 35342 30172 35348 30184
rect 29196 30144 35348 30172
rect 29196 30104 29224 30144
rect 35342 30132 35348 30144
rect 35400 30132 35406 30184
rect 26344 30076 29224 30104
rect 29641 30107 29699 30113
rect 16356 30064 16362 30076
rect 29641 30073 29653 30107
rect 29687 30104 29699 30107
rect 31110 30104 31116 30116
rect 29687 30076 31116 30104
rect 29687 30073 29699 30076
rect 29641 30067 29699 30073
rect 31110 30064 31116 30076
rect 31168 30064 31174 30116
rect 38286 30104 38292 30116
rect 38247 30076 38292 30104
rect 38286 30064 38292 30076
rect 38344 30064 38350 30116
rect 17310 30036 17316 30048
rect 15488 30008 17316 30036
rect 17310 29996 17316 30008
rect 17368 29996 17374 30048
rect 23658 30036 23664 30048
rect 23619 30008 23664 30036
rect 23658 29996 23664 30008
rect 23716 29996 23722 30048
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 24305 30039 24363 30045
rect 24305 30036 24317 30039
rect 23808 30008 24317 30036
rect 23808 29996 23814 30008
rect 24305 30005 24317 30008
rect 24351 30005 24363 30039
rect 24305 29999 24363 30005
rect 24854 29996 24860 30048
rect 24912 30036 24918 30048
rect 25225 30039 25283 30045
rect 25225 30036 25237 30039
rect 24912 30008 25237 30036
rect 24912 29996 24918 30008
rect 25225 30005 25237 30008
rect 25271 30005 25283 30039
rect 25225 29999 25283 30005
rect 26421 30039 26479 30045
rect 26421 30005 26433 30039
rect 26467 30036 26479 30039
rect 26878 30036 26884 30048
rect 26467 30008 26884 30036
rect 26467 30005 26479 30008
rect 26421 29999 26479 30005
rect 26878 29996 26884 30008
rect 26936 29996 26942 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 10686 29832 10692 29844
rect 10647 29804 10692 29832
rect 10686 29792 10692 29804
rect 10744 29792 10750 29844
rect 15378 29832 15384 29844
rect 10796 29804 14872 29832
rect 15339 29804 15384 29832
rect 9490 29724 9496 29776
rect 9548 29764 9554 29776
rect 10796 29764 10824 29804
rect 9548 29736 10824 29764
rect 9548 29724 9554 29736
rect 11146 29724 11152 29776
rect 11204 29764 11210 29776
rect 11204 29736 14688 29764
rect 11204 29724 11210 29736
rect 2590 29656 2596 29708
rect 2648 29696 2654 29708
rect 2648 29668 6684 29696
rect 2648 29656 2654 29668
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 6362 29628 6368 29640
rect 1627 29600 6368 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 6362 29588 6368 29600
rect 6420 29588 6426 29640
rect 6656 29637 6684 29668
rect 6641 29631 6699 29637
rect 6641 29597 6653 29631
rect 6687 29597 6699 29631
rect 9122 29628 9128 29640
rect 9083 29600 9128 29628
rect 6641 29591 6699 29597
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 9306 29628 9312 29640
rect 9267 29600 9312 29628
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29628 10655 29631
rect 10962 29628 10968 29640
rect 10643 29600 10968 29628
rect 10643 29597 10655 29600
rect 10597 29591 10655 29597
rect 10962 29588 10968 29600
rect 11020 29588 11026 29640
rect 13354 29628 13360 29640
rect 13315 29600 13360 29628
rect 13354 29588 13360 29600
rect 13412 29588 13418 29640
rect 14660 29637 14688 29736
rect 14645 29631 14703 29637
rect 14645 29597 14657 29631
rect 14691 29597 14703 29631
rect 14844 29628 14872 29804
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 16022 29832 16028 29844
rect 15983 29804 16028 29832
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 18598 29792 18604 29844
rect 18656 29832 18662 29844
rect 18693 29835 18751 29841
rect 18693 29832 18705 29835
rect 18656 29804 18705 29832
rect 18656 29792 18662 29804
rect 18693 29801 18705 29804
rect 18739 29801 18751 29835
rect 21910 29832 21916 29844
rect 21871 29804 21916 29832
rect 18693 29795 18751 29801
rect 21910 29792 21916 29804
rect 21968 29792 21974 29844
rect 26786 29832 26792 29844
rect 26747 29804 26792 29832
rect 26786 29792 26792 29804
rect 26844 29792 26850 29844
rect 18049 29767 18107 29773
rect 18049 29733 18061 29767
rect 18095 29764 18107 29767
rect 18095 29736 24164 29764
rect 18095 29733 18107 29736
rect 18049 29727 18107 29733
rect 15102 29656 15108 29708
rect 15160 29696 15166 29708
rect 23198 29696 23204 29708
rect 15160 29668 23204 29696
rect 15160 29656 15166 29668
rect 15948 29637 15976 29668
rect 23198 29656 23204 29668
rect 23256 29656 23262 29708
rect 15289 29631 15347 29637
rect 15289 29628 15301 29631
rect 14844 29600 15301 29628
rect 14645 29591 14703 29597
rect 15289 29597 15301 29600
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29597 15991 29631
rect 17034 29628 17040 29640
rect 16995 29600 17040 29628
rect 15933 29591 15991 29597
rect 6733 29563 6791 29569
rect 6733 29529 6745 29563
rect 6779 29560 6791 29563
rect 13630 29560 13636 29572
rect 6779 29532 13636 29560
rect 6779 29529 6791 29532
rect 6733 29523 6791 29529
rect 13630 29520 13636 29532
rect 13688 29520 13694 29572
rect 15304 29560 15332 29591
rect 17034 29588 17040 29600
rect 17092 29588 17098 29640
rect 18230 29628 18236 29640
rect 18191 29600 18236 29628
rect 18230 29588 18236 29600
rect 18288 29588 18294 29640
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29628 18935 29631
rect 21450 29628 21456 29640
rect 18923 29600 21456 29628
rect 18923 29597 18935 29600
rect 18877 29591 18935 29597
rect 21450 29588 21456 29600
rect 21508 29588 21514 29640
rect 21821 29631 21879 29637
rect 21821 29597 21833 29631
rect 21867 29628 21879 29631
rect 22738 29628 22744 29640
rect 21867 29600 22744 29628
rect 21867 29597 21879 29600
rect 21821 29591 21879 29597
rect 22738 29588 22744 29600
rect 22796 29588 22802 29640
rect 23014 29628 23020 29640
rect 22975 29600 23020 29628
rect 23014 29588 23020 29600
rect 23072 29588 23078 29640
rect 23566 29588 23572 29640
rect 23624 29628 23630 29640
rect 23661 29631 23719 29637
rect 23661 29628 23673 29631
rect 23624 29600 23673 29628
rect 23624 29588 23630 29600
rect 23661 29597 23673 29600
rect 23707 29597 23719 29631
rect 23661 29591 23719 29597
rect 16758 29560 16764 29572
rect 15304 29532 16764 29560
rect 16758 29520 16764 29532
rect 16816 29520 16822 29572
rect 1762 29492 1768 29504
rect 1723 29464 1768 29492
rect 1762 29452 1768 29464
rect 1820 29452 1826 29504
rect 9766 29492 9772 29504
rect 9727 29464 9772 29492
rect 9766 29452 9772 29464
rect 9824 29452 9830 29504
rect 13449 29495 13507 29501
rect 13449 29461 13461 29495
rect 13495 29492 13507 29495
rect 13998 29492 14004 29504
rect 13495 29464 14004 29492
rect 13495 29461 13507 29464
rect 13449 29455 13507 29461
rect 13998 29452 14004 29464
rect 14056 29452 14062 29504
rect 14737 29495 14795 29501
rect 14737 29461 14749 29495
rect 14783 29492 14795 29495
rect 15102 29492 15108 29504
rect 14783 29464 15108 29492
rect 14783 29461 14795 29464
rect 14737 29455 14795 29461
rect 15102 29452 15108 29464
rect 15160 29452 15166 29504
rect 17129 29495 17187 29501
rect 17129 29461 17141 29495
rect 17175 29492 17187 29495
rect 18690 29492 18696 29504
rect 17175 29464 18696 29492
rect 17175 29461 17187 29464
rect 17129 29455 17187 29461
rect 18690 29452 18696 29464
rect 18748 29452 18754 29504
rect 23109 29495 23167 29501
rect 23109 29461 23121 29495
rect 23155 29492 23167 29495
rect 23382 29492 23388 29504
rect 23155 29464 23388 29492
rect 23155 29461 23167 29464
rect 23109 29455 23167 29461
rect 23382 29452 23388 29464
rect 23440 29452 23446 29504
rect 23753 29495 23811 29501
rect 23753 29461 23765 29495
rect 23799 29492 23811 29495
rect 24026 29492 24032 29504
rect 23799 29464 24032 29492
rect 23799 29461 23811 29464
rect 23753 29455 23811 29461
rect 24026 29452 24032 29464
rect 24084 29452 24090 29504
rect 24136 29492 24164 29736
rect 25222 29696 25228 29708
rect 25183 29668 25228 29696
rect 25222 29656 25228 29668
rect 25280 29656 25286 29708
rect 26694 29628 26700 29640
rect 26655 29600 26700 29628
rect 26694 29588 26700 29600
rect 26752 29588 26758 29640
rect 38010 29628 38016 29640
rect 37971 29600 38016 29628
rect 38010 29588 38016 29600
rect 38068 29588 38074 29640
rect 25314 29520 25320 29572
rect 25372 29560 25378 29572
rect 25372 29532 25417 29560
rect 25372 29520 25378 29532
rect 25498 29520 25504 29572
rect 25556 29560 25562 29572
rect 26237 29563 26295 29569
rect 26237 29560 26249 29563
rect 25556 29532 26249 29560
rect 25556 29520 25562 29532
rect 26237 29529 26249 29532
rect 26283 29529 26295 29563
rect 26237 29523 26295 29529
rect 29730 29492 29736 29504
rect 24136 29464 29736 29492
rect 29730 29452 29736 29464
rect 29788 29452 29794 29504
rect 38194 29492 38200 29504
rect 38155 29464 38200 29492
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 9306 29288 9312 29300
rect 9267 29260 9312 29288
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 14642 29248 14648 29300
rect 14700 29288 14706 29300
rect 14700 29260 15240 29288
rect 14700 29248 14706 29260
rect 13081 29223 13139 29229
rect 13081 29189 13093 29223
rect 13127 29220 13139 29223
rect 13817 29223 13875 29229
rect 13817 29220 13829 29223
rect 13127 29192 13829 29220
rect 13127 29189 13139 29192
rect 13081 29183 13139 29189
rect 13817 29189 13829 29192
rect 13863 29189 13875 29223
rect 15212 29220 15240 29260
rect 20622 29248 20628 29300
rect 20680 29288 20686 29300
rect 22005 29291 22063 29297
rect 22005 29288 22017 29291
rect 20680 29260 22017 29288
rect 20680 29248 20686 29260
rect 22005 29257 22017 29260
rect 22051 29257 22063 29291
rect 25314 29288 25320 29300
rect 25275 29260 25320 29288
rect 22005 29251 22063 29257
rect 25314 29248 25320 29260
rect 25372 29248 25378 29300
rect 21818 29220 21824 29232
rect 13817 29183 13875 29189
rect 14384 29192 15148 29220
rect 15212 29192 21824 29220
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29152 1639 29155
rect 6638 29152 6644 29164
rect 1627 29124 6644 29152
rect 1627 29121 1639 29124
rect 1581 29115 1639 29121
rect 6638 29112 6644 29124
rect 6696 29112 6702 29164
rect 9217 29155 9275 29161
rect 9217 29121 9229 29155
rect 9263 29152 9275 29155
rect 11146 29152 11152 29164
rect 9263 29124 11152 29152
rect 9263 29121 9275 29124
rect 9217 29115 9275 29121
rect 11146 29112 11152 29124
rect 11204 29112 11210 29164
rect 11330 29112 11336 29164
rect 11388 29152 11394 29164
rect 11701 29155 11759 29161
rect 11701 29152 11713 29155
rect 11388 29124 11713 29152
rect 11388 29112 11394 29124
rect 11701 29121 11713 29124
rect 11747 29121 11759 29155
rect 12989 29155 13047 29161
rect 12989 29152 13001 29155
rect 11701 29115 11759 29121
rect 11808 29124 13001 29152
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 11808 29084 11836 29124
rect 12989 29121 13001 29124
rect 13035 29121 13047 29155
rect 12989 29115 13047 29121
rect 9732 29056 11836 29084
rect 12345 29087 12403 29093
rect 9732 29044 9738 29056
rect 12345 29053 12357 29087
rect 12391 29084 12403 29087
rect 13725 29087 13783 29093
rect 13725 29084 13737 29087
rect 12391 29056 13737 29084
rect 12391 29053 12403 29056
rect 12345 29047 12403 29053
rect 13725 29053 13737 29056
rect 13771 29053 13783 29087
rect 14384 29084 14412 29192
rect 15010 29152 15016 29164
rect 14971 29124 15016 29152
rect 15010 29112 15016 29124
rect 15068 29112 15074 29164
rect 14826 29084 14832 29096
rect 13725 29047 13783 29053
rect 14200 29056 14412 29084
rect 14787 29056 14832 29084
rect 1762 29016 1768 29028
rect 1723 28988 1768 29016
rect 1762 28976 1768 28988
rect 1820 28976 1826 29028
rect 12250 28976 12256 29028
rect 12308 29016 12314 29028
rect 14200 29016 14228 29056
rect 14826 29044 14832 29056
rect 14884 29044 14890 29096
rect 15120 29084 15148 29192
rect 21818 29180 21824 29192
rect 21876 29180 21882 29232
rect 23474 29220 23480 29232
rect 22204 29192 23480 29220
rect 15838 29112 15844 29164
rect 15896 29152 15902 29164
rect 16025 29155 16083 29161
rect 16025 29152 16037 29155
rect 15896 29124 16037 29152
rect 15896 29112 15902 29124
rect 16025 29121 16037 29124
rect 16071 29121 16083 29155
rect 20898 29152 20904 29164
rect 20859 29124 20904 29152
rect 16025 29115 16083 29121
rect 20898 29112 20904 29124
rect 20956 29152 20962 29164
rect 22204 29161 22232 29192
rect 23474 29180 23480 29192
rect 23532 29180 23538 29232
rect 23750 29220 23756 29232
rect 23711 29192 23756 29220
rect 23750 29180 23756 29192
rect 23808 29180 23814 29232
rect 23934 29180 23940 29232
rect 23992 29220 23998 29232
rect 27982 29220 27988 29232
rect 23992 29192 27988 29220
rect 23992 29180 23998 29192
rect 22189 29155 22247 29161
rect 20956 29124 22140 29152
rect 20956 29112 20962 29124
rect 20622 29084 20628 29096
rect 15120 29056 20628 29084
rect 20622 29044 20628 29056
rect 20680 29044 20686 29096
rect 22112 29084 22140 29124
rect 22189 29121 22201 29155
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22925 29155 22983 29161
rect 22925 29121 22937 29155
rect 22971 29121 22983 29155
rect 25222 29152 25228 29164
rect 25183 29124 25228 29152
rect 22925 29115 22983 29121
rect 22940 29084 22968 29115
rect 25222 29112 25228 29124
rect 25280 29112 25286 29164
rect 26252 29161 26280 29192
rect 27982 29180 27988 29192
rect 28040 29180 28046 29232
rect 30742 29180 30748 29232
rect 30800 29220 30806 29232
rect 30929 29223 30987 29229
rect 30929 29220 30941 29223
rect 30800 29192 30941 29220
rect 30800 29180 30806 29192
rect 30929 29189 30941 29192
rect 30975 29189 30987 29223
rect 30929 29183 30987 29189
rect 31018 29180 31024 29232
rect 31076 29220 31082 29232
rect 31076 29192 31121 29220
rect 31076 29180 31082 29192
rect 26237 29155 26295 29161
rect 26237 29121 26249 29155
rect 26283 29121 26295 29155
rect 26237 29115 26295 29121
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29152 27215 29155
rect 28902 29152 28908 29164
rect 27203 29124 28908 29152
rect 27203 29121 27215 29124
rect 27157 29115 27215 29121
rect 28902 29112 28908 29124
rect 28960 29112 28966 29164
rect 23658 29084 23664 29096
rect 22112 29056 22968 29084
rect 23619 29056 23664 29084
rect 23658 29044 23664 29056
rect 23716 29044 23722 29096
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 23937 29087 23995 29093
rect 23937 29084 23949 29087
rect 23808 29056 23949 29084
rect 23808 29044 23814 29056
rect 23937 29053 23949 29056
rect 23983 29053 23995 29087
rect 23937 29047 23995 29053
rect 24136 29056 31754 29084
rect 12308 28988 14228 29016
rect 14277 29019 14335 29025
rect 12308 28976 12314 28988
rect 14277 28985 14289 29019
rect 14323 29016 14335 29019
rect 15286 29016 15292 29028
rect 14323 28988 15292 29016
rect 14323 28985 14335 28988
rect 14277 28979 14335 28985
rect 15286 28976 15292 28988
rect 15344 28976 15350 29028
rect 16209 29019 16267 29025
rect 15396 28988 15792 29016
rect 11514 28908 11520 28960
rect 11572 28948 11578 28960
rect 11793 28951 11851 28957
rect 11793 28948 11805 28951
rect 11572 28920 11805 28948
rect 11572 28908 11578 28920
rect 11793 28917 11805 28920
rect 11839 28917 11851 28951
rect 11793 28911 11851 28917
rect 11882 28908 11888 28960
rect 11940 28948 11946 28960
rect 15396 28948 15424 28988
rect 11940 28920 15424 28948
rect 15473 28951 15531 28957
rect 11940 28908 11946 28920
rect 15473 28917 15485 28951
rect 15519 28948 15531 28951
rect 15654 28948 15660 28960
rect 15519 28920 15660 28948
rect 15519 28917 15531 28920
rect 15473 28911 15531 28917
rect 15654 28908 15660 28920
rect 15712 28908 15718 28960
rect 15764 28948 15792 28988
rect 16209 28985 16221 29019
rect 16255 29016 16267 29019
rect 16255 28994 21956 29016
rect 16255 28988 22048 28994
rect 16255 28985 16267 28988
rect 16209 28979 16267 28985
rect 21928 28966 22048 28988
rect 16114 28948 16120 28960
rect 15764 28920 16120 28948
rect 16114 28908 16120 28920
rect 16172 28908 16178 28960
rect 16390 28908 16396 28960
rect 16448 28948 16454 28960
rect 20898 28948 20904 28960
rect 16448 28920 20904 28948
rect 16448 28908 16454 28920
rect 20898 28908 20904 28920
rect 20956 28908 20962 28960
rect 20993 28951 21051 28957
rect 20993 28917 21005 28951
rect 21039 28948 21051 28951
rect 21266 28948 21272 28960
rect 21039 28920 21272 28948
rect 21039 28917 21051 28920
rect 20993 28911 21051 28917
rect 21266 28908 21272 28920
rect 21324 28908 21330 28960
rect 22020 28948 22048 28966
rect 22112 28988 22784 29016
rect 22112 28948 22140 28988
rect 22020 28920 22140 28948
rect 22756 28948 22784 28988
rect 22830 28976 22836 29028
rect 22888 29016 22894 29028
rect 23017 29019 23075 29025
rect 23017 29016 23029 29019
rect 22888 28988 23029 29016
rect 22888 28976 22894 28988
rect 23017 28985 23029 28988
rect 23063 28985 23075 29019
rect 24136 29016 24164 29056
rect 27246 29016 27252 29028
rect 23017 28979 23075 28985
rect 23124 28988 24164 29016
rect 27207 28988 27252 29016
rect 23124 28948 23152 28988
rect 27246 28976 27252 28988
rect 27304 28976 27310 29028
rect 31110 28976 31116 29028
rect 31168 29016 31174 29028
rect 31481 29019 31539 29025
rect 31481 29016 31493 29019
rect 31168 28988 31493 29016
rect 31168 28976 31174 28988
rect 31481 28985 31493 28988
rect 31527 28985 31539 29019
rect 31726 29016 31754 29056
rect 37182 29044 37188 29096
rect 37240 29084 37246 29096
rect 37461 29087 37519 29093
rect 37461 29084 37473 29087
rect 37240 29056 37473 29084
rect 37240 29044 37246 29056
rect 37461 29053 37473 29056
rect 37507 29053 37519 29087
rect 37734 29084 37740 29096
rect 37695 29056 37740 29084
rect 37461 29047 37519 29053
rect 37734 29044 37740 29056
rect 37792 29044 37798 29096
rect 35526 29016 35532 29028
rect 31726 28988 35532 29016
rect 31481 28979 31539 28985
rect 35526 28976 35532 28988
rect 35584 28976 35590 29028
rect 22756 28920 23152 28948
rect 23474 28908 23480 28960
rect 23532 28948 23538 28960
rect 26142 28948 26148 28960
rect 23532 28920 26148 28948
rect 23532 28908 23538 28920
rect 26142 28908 26148 28920
rect 26200 28908 26206 28960
rect 26326 28948 26332 28960
rect 26287 28920 26332 28948
rect 26326 28908 26332 28920
rect 26384 28908 26390 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 6362 28744 6368 28756
rect 6323 28716 6368 28744
rect 6362 28704 6368 28716
rect 6420 28704 6426 28756
rect 9766 28704 9772 28756
rect 9824 28744 9830 28756
rect 10597 28747 10655 28753
rect 10597 28744 10609 28747
rect 9824 28716 10609 28744
rect 9824 28704 9830 28716
rect 10597 28713 10609 28716
rect 10643 28713 10655 28747
rect 10597 28707 10655 28713
rect 10870 28704 10876 28756
rect 10928 28744 10934 28756
rect 10928 28716 16160 28744
rect 10928 28704 10934 28716
rect 16022 28676 16028 28688
rect 13556 28648 16028 28676
rect 9122 28568 9128 28620
rect 9180 28608 9186 28620
rect 11425 28611 11483 28617
rect 11425 28608 11437 28611
rect 9180 28580 11437 28608
rect 9180 28568 9186 28580
rect 11425 28577 11437 28580
rect 11471 28577 11483 28611
rect 11425 28571 11483 28577
rect 5721 28543 5779 28549
rect 5721 28509 5733 28543
rect 5767 28509 5779 28543
rect 5721 28503 5779 28509
rect 5813 28543 5871 28549
rect 5813 28509 5825 28543
rect 5859 28540 5871 28543
rect 6549 28543 6607 28549
rect 6549 28540 6561 28543
rect 5859 28512 6561 28540
rect 5859 28509 5871 28512
rect 5813 28503 5871 28509
rect 6549 28509 6561 28512
rect 6595 28509 6607 28543
rect 6549 28503 6607 28509
rect 5736 28472 5764 28503
rect 6730 28500 6736 28552
rect 6788 28540 6794 28552
rect 7285 28543 7343 28549
rect 7285 28540 7297 28543
rect 6788 28512 7297 28540
rect 6788 28500 6794 28512
rect 7285 28509 7297 28512
rect 7331 28509 7343 28543
rect 7285 28503 7343 28509
rect 10229 28543 10287 28549
rect 10229 28509 10241 28543
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28540 10471 28543
rect 11054 28540 11060 28552
rect 10459 28512 11060 28540
rect 10459 28509 10471 28512
rect 10413 28503 10471 28509
rect 10244 28472 10272 28503
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 12894 28540 12900 28552
rect 12855 28512 12900 28540
rect 12894 28500 12900 28512
rect 12952 28500 12958 28552
rect 13556 28549 13584 28648
rect 16022 28636 16028 28648
rect 16080 28636 16086 28688
rect 14826 28568 14832 28620
rect 14884 28608 14890 28620
rect 14884 28580 15792 28608
rect 14884 28568 14890 28580
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28509 13599 28543
rect 13541 28503 13599 28509
rect 14277 28543 14335 28549
rect 14277 28509 14289 28543
rect 14323 28540 14335 28543
rect 14550 28540 14556 28552
rect 14323 28512 14556 28540
rect 14323 28509 14335 28512
rect 14277 28503 14335 28509
rect 14550 28500 14556 28512
rect 14608 28500 14614 28552
rect 11422 28472 11428 28484
rect 5736 28444 9076 28472
rect 10244 28444 11428 28472
rect 7377 28407 7435 28413
rect 7377 28373 7389 28407
rect 7423 28404 7435 28407
rect 7466 28404 7472 28416
rect 7423 28376 7472 28404
rect 7423 28373 7435 28376
rect 7377 28367 7435 28373
rect 7466 28364 7472 28376
rect 7524 28364 7530 28416
rect 9048 28404 9076 28444
rect 11422 28432 11428 28444
rect 11480 28432 11486 28484
rect 11514 28432 11520 28484
rect 11572 28472 11578 28484
rect 11572 28444 11617 28472
rect 11572 28432 11578 28444
rect 12434 28432 12440 28484
rect 12492 28472 12498 28484
rect 13633 28475 13691 28481
rect 12492 28444 12537 28472
rect 12492 28432 12498 28444
rect 13633 28441 13645 28475
rect 13679 28472 13691 28475
rect 14458 28472 14464 28484
rect 13679 28444 14464 28472
rect 13679 28441 13691 28444
rect 13633 28435 13691 28441
rect 14458 28432 14464 28444
rect 14516 28432 14522 28484
rect 14734 28432 14740 28484
rect 14792 28472 14798 28484
rect 15010 28472 15016 28484
rect 14792 28444 15016 28472
rect 14792 28432 14798 28444
rect 15010 28432 15016 28444
rect 15068 28432 15074 28484
rect 15102 28432 15108 28484
rect 15160 28472 15166 28484
rect 15160 28444 15205 28472
rect 15160 28432 15166 28444
rect 15286 28432 15292 28484
rect 15344 28472 15350 28484
rect 15657 28475 15715 28481
rect 15657 28472 15669 28475
rect 15344 28444 15669 28472
rect 15344 28432 15350 28444
rect 15657 28441 15669 28444
rect 15703 28441 15715 28475
rect 15764 28472 15792 28580
rect 16132 28549 16160 28716
rect 17310 28704 17316 28756
rect 17368 28744 17374 28756
rect 17368 28716 21404 28744
rect 17368 28704 17374 28716
rect 16206 28568 16212 28620
rect 16264 28608 16270 28620
rect 19352 28608 19380 28716
rect 19426 28636 19432 28688
rect 19484 28676 19490 28688
rect 20254 28676 20260 28688
rect 19484 28648 20260 28676
rect 19484 28636 19490 28648
rect 20254 28636 20260 28648
rect 20312 28636 20318 28688
rect 21376 28620 21404 28716
rect 22002 28704 22008 28756
rect 22060 28744 22066 28756
rect 22060 28716 31754 28744
rect 22060 28704 22066 28716
rect 30653 28679 30711 28685
rect 30653 28645 30665 28679
rect 30699 28676 30711 28679
rect 31018 28676 31024 28688
rect 30699 28648 31024 28676
rect 30699 28645 30711 28648
rect 30653 28639 30711 28645
rect 31018 28636 31024 28648
rect 31076 28636 31082 28688
rect 31726 28676 31754 28716
rect 33134 28676 33140 28688
rect 31726 28648 33140 28676
rect 33134 28636 33140 28648
rect 33192 28636 33198 28688
rect 19521 28611 19579 28617
rect 19521 28608 19533 28611
rect 16264 28580 19288 28608
rect 19352 28580 19533 28608
rect 16264 28568 16270 28580
rect 16117 28543 16175 28549
rect 16117 28509 16129 28543
rect 16163 28509 16175 28543
rect 16758 28540 16764 28552
rect 16719 28512 16764 28540
rect 16117 28503 16175 28509
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 19260 28540 19288 28580
rect 19521 28577 19533 28580
rect 19567 28577 19579 28611
rect 20070 28608 20076 28620
rect 20031 28580 20076 28608
rect 19521 28571 19579 28577
rect 20070 28568 20076 28580
rect 20128 28608 20134 28620
rect 20346 28608 20352 28620
rect 20128 28580 20352 28608
rect 20128 28568 20134 28580
rect 20346 28568 20352 28580
rect 20404 28568 20410 28620
rect 21358 28568 21364 28620
rect 21416 28608 21422 28620
rect 21453 28611 21511 28617
rect 21453 28608 21465 28611
rect 21416 28580 21465 28608
rect 21416 28568 21422 28580
rect 21453 28577 21465 28580
rect 21499 28577 21511 28611
rect 21453 28571 21511 28577
rect 22756 28580 25268 28608
rect 22756 28552 22784 28580
rect 19334 28540 19340 28552
rect 19260 28512 19340 28540
rect 19334 28500 19340 28512
rect 19392 28500 19398 28552
rect 22649 28543 22707 28549
rect 22649 28509 22661 28543
rect 22695 28540 22707 28543
rect 22738 28540 22744 28552
rect 22695 28512 22744 28540
rect 22695 28509 22707 28512
rect 22649 28503 22707 28509
rect 22738 28500 22744 28512
rect 22796 28500 22802 28552
rect 23293 28543 23351 28549
rect 23293 28509 23305 28543
rect 23339 28540 23351 28543
rect 24210 28540 24216 28552
rect 23339 28512 24216 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 24210 28500 24216 28512
rect 24268 28500 24274 28552
rect 24581 28543 24639 28549
rect 24581 28509 24593 28543
rect 24627 28540 24639 28543
rect 25130 28540 25136 28552
rect 24627 28512 25136 28540
rect 24627 28509 24639 28512
rect 24581 28503 24639 28509
rect 25130 28500 25136 28512
rect 25188 28500 25194 28552
rect 25240 28549 25268 28580
rect 26142 28568 26148 28620
rect 26200 28608 26206 28620
rect 37734 28608 37740 28620
rect 26200 28580 37740 28608
rect 26200 28568 26206 28580
rect 28276 28549 28304 28580
rect 37734 28568 37740 28580
rect 37792 28568 37798 28620
rect 25225 28543 25283 28549
rect 25225 28509 25237 28543
rect 25271 28509 25283 28543
rect 25225 28503 25283 28509
rect 28261 28543 28319 28549
rect 28261 28509 28273 28543
rect 28307 28509 28319 28543
rect 28261 28503 28319 28509
rect 28997 28543 29055 28549
rect 28997 28509 29009 28543
rect 29043 28540 29055 28543
rect 30561 28543 30619 28549
rect 30561 28540 30573 28543
rect 29043 28512 30573 28540
rect 29043 28509 29055 28512
rect 28997 28503 29055 28509
rect 30561 28509 30573 28512
rect 30607 28540 30619 28543
rect 32122 28540 32128 28552
rect 30607 28512 32128 28540
rect 30607 28509 30619 28512
rect 30561 28503 30619 28509
rect 32122 28500 32128 28512
rect 32180 28500 32186 28552
rect 17770 28472 17776 28484
rect 15764 28444 17776 28472
rect 15657 28435 15715 28441
rect 12894 28404 12900 28416
rect 9048 28376 12900 28404
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 12989 28407 13047 28413
rect 12989 28373 13001 28407
rect 13035 28404 13047 28407
rect 14182 28404 14188 28416
rect 13035 28376 14188 28404
rect 13035 28373 13047 28376
rect 12989 28367 13047 28373
rect 14182 28364 14188 28376
rect 14240 28364 14246 28416
rect 14366 28404 14372 28416
rect 14327 28376 14372 28404
rect 14366 28364 14372 28376
rect 14424 28364 14430 28416
rect 15672 28404 15700 28435
rect 17770 28432 17776 28444
rect 17828 28432 17834 28484
rect 19613 28475 19671 28481
rect 19613 28441 19625 28475
rect 19659 28441 19671 28475
rect 19613 28435 19671 28441
rect 21177 28475 21235 28481
rect 21177 28441 21189 28475
rect 21223 28441 21235 28475
rect 21177 28435 21235 28441
rect 15746 28404 15752 28416
rect 15672 28376 15752 28404
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 16022 28364 16028 28416
rect 16080 28404 16086 28416
rect 16209 28407 16267 28413
rect 16209 28404 16221 28407
rect 16080 28376 16221 28404
rect 16080 28364 16086 28376
rect 16209 28373 16221 28376
rect 16255 28373 16267 28407
rect 16850 28404 16856 28416
rect 16811 28376 16856 28404
rect 16209 28367 16267 28373
rect 16850 28364 16856 28376
rect 16908 28364 16914 28416
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 19628 28404 19656 28435
rect 19484 28376 19656 28404
rect 21192 28404 21220 28435
rect 21266 28432 21272 28484
rect 21324 28472 21330 28484
rect 21324 28444 21369 28472
rect 21324 28432 21330 28444
rect 24026 28432 24032 28484
rect 24084 28472 24090 28484
rect 25038 28472 25044 28484
rect 24084 28444 25044 28472
rect 24084 28432 24090 28444
rect 25038 28432 25044 28444
rect 25096 28472 25102 28484
rect 25961 28475 26019 28481
rect 25961 28472 25973 28475
rect 25096 28444 25973 28472
rect 25096 28432 25102 28444
rect 25961 28441 25973 28444
rect 26007 28441 26019 28475
rect 25961 28435 26019 28441
rect 26053 28475 26111 28481
rect 26053 28441 26065 28475
rect 26099 28472 26111 28475
rect 26326 28472 26332 28484
rect 26099 28444 26332 28472
rect 26099 28441 26111 28444
rect 26053 28435 26111 28441
rect 26326 28432 26332 28444
rect 26384 28432 26390 28484
rect 26970 28472 26976 28484
rect 26931 28444 26976 28472
rect 26970 28432 26976 28444
rect 27028 28432 27034 28484
rect 28353 28475 28411 28481
rect 28353 28441 28365 28475
rect 28399 28472 28411 28475
rect 29178 28472 29184 28484
rect 28399 28444 29184 28472
rect 28399 28441 28411 28444
rect 28353 28435 28411 28441
rect 29178 28432 29184 28444
rect 29236 28432 29242 28484
rect 21818 28404 21824 28416
rect 21192 28376 21824 28404
rect 19484 28364 19490 28376
rect 21818 28364 21824 28376
rect 21876 28364 21882 28416
rect 22741 28407 22799 28413
rect 22741 28373 22753 28407
rect 22787 28404 22799 28407
rect 23106 28404 23112 28416
rect 22787 28376 23112 28404
rect 22787 28373 22799 28376
rect 22741 28367 22799 28373
rect 23106 28364 23112 28376
rect 23164 28364 23170 28416
rect 23290 28364 23296 28416
rect 23348 28404 23354 28416
rect 23385 28407 23443 28413
rect 23385 28404 23397 28407
rect 23348 28376 23397 28404
rect 23348 28364 23354 28376
rect 23385 28373 23397 28376
rect 23431 28373 23443 28407
rect 23385 28367 23443 28373
rect 24673 28407 24731 28413
rect 24673 28373 24685 28407
rect 24719 28404 24731 28407
rect 24762 28404 24768 28416
rect 24719 28376 24768 28404
rect 24719 28373 24731 28376
rect 24673 28367 24731 28373
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 24854 28364 24860 28416
rect 24912 28404 24918 28416
rect 25317 28407 25375 28413
rect 25317 28404 25329 28407
rect 24912 28376 25329 28404
rect 24912 28364 24918 28376
rect 25317 28373 25329 28376
rect 25363 28373 25375 28407
rect 25317 28367 25375 28373
rect 28626 28364 28632 28416
rect 28684 28404 28690 28416
rect 29089 28407 29147 28413
rect 29089 28404 29101 28407
rect 28684 28376 29101 28404
rect 28684 28364 28690 28376
rect 29089 28373 29101 28376
rect 29135 28373 29147 28407
rect 29089 28367 29147 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 6638 28200 6644 28212
rect 6599 28172 6644 28200
rect 6638 28160 6644 28172
rect 6696 28160 6702 28212
rect 8389 28203 8447 28209
rect 8389 28169 8401 28203
rect 8435 28200 8447 28203
rect 14826 28200 14832 28212
rect 8435 28172 14832 28200
rect 8435 28169 8447 28172
rect 8389 28163 8447 28169
rect 14826 28160 14832 28172
rect 14884 28160 14890 28212
rect 16850 28200 16856 28212
rect 15396 28172 16856 28200
rect 1854 28092 1860 28144
rect 1912 28132 1918 28144
rect 1912 28104 8984 28132
rect 1912 28092 1918 28104
rect 6825 28067 6883 28073
rect 6825 28033 6837 28067
rect 6871 28033 6883 28067
rect 6825 28027 6883 28033
rect 7285 28067 7343 28073
rect 7285 28033 7297 28067
rect 7331 28064 7343 28067
rect 8294 28064 8300 28076
rect 7331 28036 8156 28064
rect 8255 28036 8300 28064
rect 7331 28033 7343 28036
rect 7285 28027 7343 28033
rect 6840 27996 6868 28027
rect 7377 27999 7435 28005
rect 7377 27996 7389 27999
rect 6840 27968 7389 27996
rect 7377 27965 7389 27968
rect 7423 27965 7435 27999
rect 8128 27996 8156 28036
rect 8294 28024 8300 28036
rect 8352 28024 8358 28076
rect 8956 28073 8984 28104
rect 9858 28092 9864 28144
rect 9916 28132 9922 28144
rect 13814 28132 13820 28144
rect 9916 28104 13820 28132
rect 9916 28092 9922 28104
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 8941 28067 8999 28073
rect 8941 28033 8953 28067
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 9033 28067 9091 28073
rect 9033 28033 9045 28067
rect 9079 28064 9091 28067
rect 10505 28067 10563 28073
rect 10505 28064 10517 28067
rect 9079 28036 10517 28064
rect 9079 28033 9091 28036
rect 9033 28027 9091 28033
rect 10505 28033 10517 28036
rect 10551 28064 10563 28067
rect 11422 28064 11428 28076
rect 10551 28036 11428 28064
rect 10551 28033 10563 28036
rect 10505 28027 10563 28033
rect 11422 28024 11428 28036
rect 11480 28024 11486 28076
rect 11698 28024 11704 28076
rect 11756 28064 11762 28076
rect 12066 28064 12072 28076
rect 11756 28036 12072 28064
rect 11756 28024 11762 28036
rect 12066 28024 12072 28036
rect 12124 28024 12130 28076
rect 13906 28024 13912 28076
rect 13964 28064 13970 28076
rect 14645 28067 14703 28073
rect 13964 28036 14596 28064
rect 13964 28024 13970 28036
rect 9582 27996 9588 28008
rect 8128 27968 9588 27996
rect 7377 27959 7435 27965
rect 9582 27956 9588 27968
rect 9640 27956 9646 28008
rect 10686 27996 10692 28008
rect 10647 27968 10692 27996
rect 10686 27956 10692 27968
rect 10744 27956 10750 28008
rect 12710 27996 12716 28008
rect 12671 27968 12716 27996
rect 12710 27956 12716 27968
rect 12768 27956 12774 28008
rect 13170 27956 13176 28008
rect 13228 27996 13234 28008
rect 13357 27999 13415 28005
rect 13357 27996 13369 27999
rect 13228 27968 13369 27996
rect 13228 27956 13234 27968
rect 13357 27965 13369 27968
rect 13403 27965 13415 27999
rect 13538 27996 13544 28008
rect 13499 27968 13544 27996
rect 13357 27959 13415 27965
rect 13538 27956 13544 27968
rect 13596 27956 13602 28008
rect 14461 27999 14519 28005
rect 14461 27965 14473 27999
rect 14507 27965 14519 27999
rect 14568 27996 14596 28036
rect 14645 28033 14657 28067
rect 14691 28064 14703 28067
rect 15396 28064 15424 28172
rect 16850 28160 16856 28172
rect 16908 28160 16914 28212
rect 21269 28203 21327 28209
rect 21269 28169 21281 28203
rect 21315 28200 21327 28203
rect 22922 28200 22928 28212
rect 21315 28172 22928 28200
rect 21315 28169 21327 28172
rect 21269 28163 21327 28169
rect 22922 28160 22928 28172
rect 22980 28160 22986 28212
rect 23750 28200 23756 28212
rect 23124 28172 23756 28200
rect 15749 28135 15807 28141
rect 15749 28132 15761 28135
rect 14691 28036 15424 28064
rect 15488 28104 15761 28132
rect 14691 28033 14703 28036
rect 14645 28027 14703 28033
rect 15488 27996 15516 28104
rect 15749 28101 15761 28104
rect 15795 28101 15807 28135
rect 16298 28132 16304 28144
rect 16259 28104 16304 28132
rect 15749 28095 15807 28101
rect 16298 28092 16304 28104
rect 16356 28092 16362 28144
rect 17862 28132 17868 28144
rect 17823 28104 17868 28132
rect 17862 28092 17868 28104
rect 17920 28092 17926 28144
rect 18785 28135 18843 28141
rect 18785 28101 18797 28135
rect 18831 28132 18843 28135
rect 23124 28132 23152 28172
rect 23750 28160 23756 28172
rect 23808 28200 23814 28212
rect 28994 28200 29000 28212
rect 23808 28172 29000 28200
rect 23808 28160 23814 28172
rect 28994 28160 29000 28172
rect 29052 28160 29058 28212
rect 23290 28132 23296 28144
rect 18831 28104 23152 28132
rect 23251 28104 23296 28132
rect 18831 28101 18843 28104
rect 18785 28095 18843 28101
rect 23290 28092 23296 28104
rect 23348 28092 23354 28144
rect 24854 28132 24860 28144
rect 24815 28104 24860 28132
rect 24854 28092 24860 28104
rect 24912 28092 24918 28144
rect 25774 28132 25780 28144
rect 25735 28104 25780 28132
rect 25774 28092 25780 28104
rect 25832 28092 25838 28144
rect 28626 28132 28632 28144
rect 28587 28104 28632 28132
rect 28626 28092 28632 28104
rect 28684 28092 28690 28144
rect 29086 28092 29092 28144
rect 29144 28132 29150 28144
rect 30101 28135 30159 28141
rect 30101 28132 30113 28135
rect 29144 28104 30113 28132
rect 29144 28092 29150 28104
rect 30101 28101 30113 28104
rect 30147 28101 30159 28135
rect 30101 28095 30159 28101
rect 30193 28135 30251 28141
rect 30193 28101 30205 28135
rect 30239 28132 30251 28135
rect 30466 28132 30472 28144
rect 30239 28104 30472 28132
rect 30239 28101 30251 28104
rect 30193 28095 30251 28101
rect 30466 28092 30472 28104
rect 30524 28092 30530 28144
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28064 16911 28067
rect 16942 28064 16948 28076
rect 16899 28036 16948 28064
rect 16899 28033 16911 28036
rect 16853 28027 16911 28033
rect 16942 28024 16948 28036
rect 17000 28024 17006 28076
rect 18966 28024 18972 28076
rect 19024 28064 19030 28076
rect 19245 28067 19303 28073
rect 19245 28064 19257 28067
rect 19024 28036 19257 28064
rect 19024 28024 19030 28036
rect 19245 28033 19257 28036
rect 19291 28033 19303 28067
rect 19245 28027 19303 28033
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 20165 28067 20223 28073
rect 20165 28064 20177 28067
rect 19392 28036 20177 28064
rect 19392 28024 19398 28036
rect 20165 28033 20177 28036
rect 20211 28064 20223 28067
rect 20622 28064 20628 28076
rect 20211 28036 20628 28064
rect 20211 28033 20223 28036
rect 20165 28027 20223 28033
rect 20622 28024 20628 28036
rect 20680 28024 20686 28076
rect 20990 28024 20996 28076
rect 21048 28064 21054 28076
rect 21453 28067 21511 28073
rect 21453 28064 21465 28067
rect 21048 28036 21465 28064
rect 21048 28024 21054 28036
rect 21453 28033 21465 28036
rect 21499 28033 21511 28067
rect 21453 28027 21511 28033
rect 21542 28024 21548 28076
rect 21600 28064 21606 28076
rect 22002 28064 22008 28076
rect 21600 28036 22008 28064
rect 21600 28024 21606 28036
rect 22002 28024 22008 28036
rect 22060 28064 22066 28076
rect 22097 28067 22155 28073
rect 22097 28064 22109 28067
rect 22060 28036 22109 28064
rect 22060 28024 22066 28036
rect 22097 28033 22109 28036
rect 22143 28033 22155 28067
rect 26234 28064 26240 28076
rect 26195 28036 26240 28064
rect 22097 28027 22155 28033
rect 26234 28024 26240 28036
rect 26292 28064 26298 28076
rect 26510 28064 26516 28076
rect 26292 28036 26516 28064
rect 26292 28024 26298 28036
rect 26510 28024 26516 28036
rect 26568 28024 26574 28076
rect 27154 28064 27160 28076
rect 27115 28036 27160 28064
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27706 28024 27712 28076
rect 27764 28064 27770 28076
rect 27801 28067 27859 28073
rect 27801 28064 27813 28067
rect 27764 28036 27813 28064
rect 27764 28024 27770 28036
rect 27801 28033 27813 28036
rect 27847 28033 27859 28067
rect 27801 28027 27859 28033
rect 15654 27996 15660 28008
rect 14568 27968 15516 27996
rect 15615 27968 15660 27996
rect 14461 27959 14519 27965
rect 14476 27928 14504 27959
rect 15654 27956 15660 27968
rect 15712 27956 15718 28008
rect 16132 27968 17724 27996
rect 16132 27928 16160 27968
rect 14476 27900 16160 27928
rect 17696 27928 17724 27968
rect 17770 27956 17776 28008
rect 17828 27996 17834 28008
rect 23201 27999 23259 28005
rect 17828 27968 17873 27996
rect 17828 27956 17834 27968
rect 23201 27965 23213 27999
rect 23247 27996 23259 27999
rect 23382 27996 23388 28008
rect 23247 27968 23388 27996
rect 23247 27965 23259 27968
rect 23201 27959 23259 27965
rect 23382 27956 23388 27968
rect 23440 27956 23446 28008
rect 23750 27996 23756 28008
rect 23711 27968 23756 27996
rect 23750 27956 23756 27968
rect 23808 27956 23814 28008
rect 24578 27956 24584 28008
rect 24636 27996 24642 28008
rect 24765 27999 24823 28005
rect 24765 27996 24777 27999
rect 24636 27968 24777 27996
rect 24636 27956 24642 27968
rect 24765 27965 24777 27968
rect 24811 27996 24823 27999
rect 26329 27999 26387 28005
rect 26329 27996 26341 27999
rect 24811 27968 26341 27996
rect 24811 27965 24823 27968
rect 24765 27959 24823 27965
rect 26329 27965 26341 27968
rect 26375 27965 26387 27999
rect 26329 27959 26387 27965
rect 28074 27956 28080 28008
rect 28132 27996 28138 28008
rect 28537 27999 28595 28005
rect 28537 27996 28549 27999
rect 28132 27968 28549 27996
rect 28132 27956 28138 27968
rect 28537 27965 28549 27968
rect 28583 27965 28595 27999
rect 28994 27996 29000 28008
rect 28955 27968 29000 27996
rect 28537 27959 28595 27965
rect 28994 27956 29000 27968
rect 29052 27996 29058 28008
rect 29546 27996 29552 28008
rect 29052 27968 29552 27996
rect 29052 27956 29058 27968
rect 29546 27956 29552 27968
rect 29604 27956 29610 28008
rect 30745 27999 30803 28005
rect 30745 27965 30757 27999
rect 30791 27996 30803 27999
rect 33962 27996 33968 28008
rect 30791 27968 33968 27996
rect 30791 27965 30803 27968
rect 30745 27959 30803 27965
rect 33962 27956 33968 27968
rect 34020 27956 34026 28008
rect 25498 27928 25504 27940
rect 17696 27900 25504 27928
rect 25498 27888 25504 27900
rect 25556 27888 25562 27940
rect 11149 27863 11207 27869
rect 11149 27829 11161 27863
rect 11195 27860 11207 27863
rect 11974 27860 11980 27872
rect 11195 27832 11980 27860
rect 11195 27829 11207 27832
rect 11149 27823 11207 27829
rect 11974 27820 11980 27832
rect 12032 27820 12038 27872
rect 12158 27860 12164 27872
rect 12119 27832 12164 27860
rect 12158 27820 12164 27832
rect 12216 27820 12222 27872
rect 14001 27863 14059 27869
rect 14001 27829 14013 27863
rect 14047 27860 14059 27863
rect 14829 27863 14887 27869
rect 14829 27860 14841 27863
rect 14047 27832 14841 27860
rect 14047 27829 14059 27832
rect 14001 27823 14059 27829
rect 14829 27829 14841 27832
rect 14875 27860 14887 27863
rect 15654 27860 15660 27872
rect 14875 27832 15660 27860
rect 14875 27829 14887 27832
rect 14829 27823 14887 27829
rect 15654 27820 15660 27832
rect 15712 27820 15718 27872
rect 16942 27860 16948 27872
rect 16903 27832 16948 27860
rect 16942 27820 16948 27832
rect 17000 27820 17006 27872
rect 19334 27860 19340 27872
rect 19295 27832 19340 27860
rect 19334 27820 19340 27832
rect 19392 27820 19398 27872
rect 20257 27863 20315 27869
rect 20257 27829 20269 27863
rect 20303 27860 20315 27863
rect 20438 27860 20444 27872
rect 20303 27832 20444 27860
rect 20303 27829 20315 27832
rect 20257 27823 20315 27829
rect 20438 27820 20444 27832
rect 20496 27820 20502 27872
rect 22186 27820 22192 27872
rect 22244 27860 22250 27872
rect 22244 27832 22289 27860
rect 22244 27820 22250 27832
rect 26418 27820 26424 27872
rect 26476 27860 26482 27872
rect 27249 27863 27307 27869
rect 27249 27860 27261 27863
rect 26476 27832 27261 27860
rect 26476 27820 26482 27832
rect 27249 27829 27261 27832
rect 27295 27829 27307 27863
rect 27890 27860 27896 27872
rect 27851 27832 27896 27860
rect 27249 27823 27307 27829
rect 27890 27820 27896 27832
rect 27948 27820 27954 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 9766 27616 9772 27668
rect 9824 27656 9830 27668
rect 9953 27659 10011 27665
rect 9953 27656 9965 27659
rect 9824 27628 9965 27656
rect 9824 27616 9830 27628
rect 9953 27625 9965 27628
rect 9999 27625 10011 27659
rect 9953 27619 10011 27625
rect 12268 27628 13676 27656
rect 7466 27520 7472 27532
rect 7427 27492 7472 27520
rect 7466 27480 7472 27492
rect 7524 27480 7530 27532
rect 9968 27520 9996 27619
rect 10781 27523 10839 27529
rect 10781 27520 10793 27523
rect 9968 27492 10793 27520
rect 10781 27489 10793 27492
rect 10827 27489 10839 27523
rect 10781 27483 10839 27489
rect 10962 27480 10968 27532
rect 11020 27520 11026 27532
rect 11057 27523 11115 27529
rect 11057 27520 11069 27523
rect 11020 27492 11069 27520
rect 11020 27480 11026 27492
rect 11057 27489 11069 27492
rect 11103 27520 11115 27523
rect 11103 27492 11560 27520
rect 11103 27489 11115 27492
rect 11057 27483 11115 27489
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27452 1639 27455
rect 4062 27452 4068 27464
rect 1627 27424 4068 27452
rect 1627 27421 1639 27424
rect 1581 27415 1639 27421
rect 4062 27412 4068 27424
rect 4120 27412 4126 27464
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27421 9643 27455
rect 9766 27452 9772 27464
rect 9727 27424 9772 27452
rect 9585 27415 9643 27421
rect 7558 27384 7564 27396
rect 7519 27356 7564 27384
rect 7558 27344 7564 27356
rect 7616 27344 7622 27396
rect 8478 27384 8484 27396
rect 8439 27356 8484 27384
rect 8478 27344 8484 27356
rect 8536 27344 8542 27396
rect 9600 27384 9628 27415
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 10778 27384 10784 27396
rect 9600 27356 10784 27384
rect 10778 27344 10784 27356
rect 10836 27344 10842 27396
rect 10873 27387 10931 27393
rect 10873 27353 10885 27387
rect 10919 27353 10931 27387
rect 11532 27384 11560 27492
rect 12268 27464 12296 27628
rect 12345 27591 12403 27597
rect 12345 27557 12357 27591
rect 12391 27588 12403 27591
rect 13538 27588 13544 27600
rect 12391 27560 13544 27588
rect 12391 27557 12403 27560
rect 12345 27551 12403 27557
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 13648 27588 13676 27628
rect 13814 27616 13820 27668
rect 13872 27656 13878 27668
rect 16850 27656 16856 27668
rect 13872 27628 16856 27656
rect 13872 27616 13878 27628
rect 16850 27616 16856 27628
rect 16908 27616 16914 27668
rect 17589 27659 17647 27665
rect 17589 27625 17601 27659
rect 17635 27656 17647 27659
rect 17862 27656 17868 27668
rect 17635 27628 17868 27656
rect 17635 27625 17647 27628
rect 17589 27619 17647 27625
rect 17862 27616 17868 27628
rect 17920 27616 17926 27668
rect 20714 27616 20720 27668
rect 20772 27656 20778 27668
rect 23658 27656 23664 27668
rect 20772 27628 23664 27656
rect 20772 27616 20778 27628
rect 23658 27616 23664 27628
rect 23716 27656 23722 27668
rect 23716 27628 24440 27656
rect 23716 27616 23722 27628
rect 14550 27588 14556 27600
rect 13648 27560 14556 27588
rect 14550 27548 14556 27560
rect 14608 27548 14614 27600
rect 15010 27548 15016 27600
rect 15068 27588 15074 27600
rect 21542 27588 21548 27600
rect 15068 27560 19380 27588
rect 15068 27548 15074 27560
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 12820 27492 13277 27520
rect 12250 27452 12256 27464
rect 12211 27424 12256 27452
rect 12250 27412 12256 27424
rect 12308 27412 12314 27464
rect 12526 27384 12532 27396
rect 11532 27356 12532 27384
rect 10873 27347 10931 27353
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 10888 27316 10916 27347
rect 12526 27344 12532 27356
rect 12584 27384 12590 27396
rect 12820 27384 12848 27492
rect 13265 27489 13277 27492
rect 13311 27489 13323 27523
rect 13265 27483 13323 27489
rect 13630 27480 13636 27532
rect 13688 27520 13694 27532
rect 14369 27523 14427 27529
rect 14369 27520 14381 27523
rect 13688 27492 14381 27520
rect 13688 27480 13694 27492
rect 14369 27489 14381 27492
rect 14415 27489 14427 27523
rect 16298 27520 16304 27532
rect 16259 27492 16304 27520
rect 14369 27483 14427 27489
rect 16298 27480 16304 27492
rect 16356 27480 16362 27532
rect 15746 27452 15752 27464
rect 15212 27424 15752 27452
rect 12584 27356 12848 27384
rect 12989 27387 13047 27393
rect 12584 27344 12590 27356
rect 12989 27353 13001 27387
rect 13035 27353 13047 27387
rect 12989 27347 13047 27353
rect 13081 27387 13139 27393
rect 13081 27353 13093 27387
rect 13127 27384 13139 27387
rect 14090 27384 14096 27396
rect 13127 27356 14096 27384
rect 13127 27353 13139 27356
rect 13081 27347 13139 27353
rect 11514 27316 11520 27328
rect 10888 27288 11520 27316
rect 11514 27276 11520 27288
rect 11572 27276 11578 27328
rect 13004 27316 13032 27347
rect 14090 27344 14096 27356
rect 14148 27344 14154 27396
rect 14458 27344 14464 27396
rect 14516 27384 14522 27396
rect 14516 27356 14561 27384
rect 14516 27344 14522 27356
rect 15212 27316 15240 27424
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16758 27412 16764 27464
rect 16816 27452 16822 27464
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 16816 27424 17509 27452
rect 16816 27412 16822 27424
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 15381 27387 15439 27393
rect 15381 27353 15393 27387
rect 15427 27384 15439 27387
rect 15654 27384 15660 27396
rect 15427 27356 15660 27384
rect 15427 27353 15439 27356
rect 15381 27347 15439 27353
rect 15654 27344 15660 27356
rect 15712 27344 15718 27396
rect 15930 27384 15936 27396
rect 15891 27356 15936 27384
rect 15930 27344 15936 27356
rect 15988 27344 15994 27396
rect 16025 27387 16083 27393
rect 16025 27353 16037 27387
rect 16071 27353 16083 27387
rect 16025 27347 16083 27353
rect 13004 27288 15240 27316
rect 15470 27276 15476 27328
rect 15528 27316 15534 27328
rect 16040 27316 16068 27347
rect 16942 27344 16948 27396
rect 17000 27384 17006 27396
rect 18233 27387 18291 27393
rect 18233 27384 18245 27387
rect 17000 27356 18245 27384
rect 17000 27344 17006 27356
rect 18233 27353 18245 27356
rect 18279 27353 18291 27387
rect 18233 27347 18291 27353
rect 18325 27387 18383 27393
rect 18325 27353 18337 27387
rect 18371 27353 18383 27387
rect 18325 27347 18383 27353
rect 18877 27387 18935 27393
rect 18877 27353 18889 27387
rect 18923 27384 18935 27387
rect 19242 27384 19248 27396
rect 18923 27356 19248 27384
rect 18923 27353 18935 27356
rect 18877 27347 18935 27353
rect 15528 27288 16068 27316
rect 18340 27316 18368 27347
rect 19242 27344 19248 27356
rect 19300 27344 19306 27396
rect 19352 27384 19380 27560
rect 19444 27560 21548 27588
rect 19444 27461 19472 27560
rect 21542 27548 21548 27560
rect 21600 27548 21606 27600
rect 21818 27548 21824 27600
rect 21876 27588 21882 27600
rect 24412 27588 24440 27628
rect 26234 27616 26240 27668
rect 26292 27656 26298 27668
rect 26292 27628 31754 27656
rect 26292 27616 26298 27628
rect 30466 27588 30472 27600
rect 21876 27560 23612 27588
rect 24412 27560 25912 27588
rect 30427 27560 30472 27588
rect 21876 27548 21882 27560
rect 19521 27523 19579 27529
rect 19521 27489 19533 27523
rect 19567 27520 19579 27523
rect 20346 27520 20352 27532
rect 19567 27492 20352 27520
rect 19567 27489 19579 27492
rect 19521 27483 19579 27489
rect 20346 27480 20352 27492
rect 20404 27480 20410 27532
rect 23017 27523 23075 27529
rect 23017 27520 23029 27523
rect 21192 27492 23029 27520
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 20165 27387 20223 27393
rect 20165 27384 20177 27387
rect 19352 27356 20177 27384
rect 20165 27353 20177 27356
rect 20211 27353 20223 27387
rect 20165 27347 20223 27353
rect 20257 27387 20315 27393
rect 20257 27353 20269 27387
rect 20303 27353 20315 27387
rect 20806 27384 20812 27396
rect 20767 27356 20812 27384
rect 20257 27347 20315 27353
rect 19334 27316 19340 27328
rect 18340 27288 19340 27316
rect 15528 27276 15534 27288
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 20272 27316 20300 27347
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 21192 27316 21220 27492
rect 23017 27489 23029 27492
rect 23063 27489 23075 27523
rect 23584 27520 23612 27560
rect 24673 27523 24731 27529
rect 23584 27492 24072 27520
rect 23017 27483 23075 27489
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23474 27452 23480 27464
rect 22971 27424 23480 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 23569 27455 23627 27461
rect 23569 27421 23581 27455
rect 23615 27452 23627 27455
rect 23934 27452 23940 27464
rect 23615 27424 23940 27452
rect 23615 27421 23627 27424
rect 23569 27415 23627 27421
rect 23934 27412 23940 27424
rect 23992 27412 23998 27464
rect 21818 27384 21824 27396
rect 21779 27356 21824 27384
rect 21818 27344 21824 27356
rect 21876 27344 21882 27396
rect 21913 27387 21971 27393
rect 21913 27353 21925 27387
rect 21959 27353 21971 27387
rect 21913 27347 21971 27353
rect 20272 27288 21220 27316
rect 21928 27316 21956 27347
rect 22002 27344 22008 27396
rect 22060 27384 22066 27396
rect 22465 27387 22523 27393
rect 22465 27384 22477 27387
rect 22060 27356 22477 27384
rect 22060 27344 22066 27356
rect 22465 27353 22477 27356
rect 22511 27353 22523 27387
rect 23661 27387 23719 27393
rect 23661 27384 23673 27387
rect 22465 27347 22523 27353
rect 22848 27356 23673 27384
rect 22848 27316 22876 27356
rect 23661 27353 23673 27356
rect 23707 27353 23719 27387
rect 24044 27384 24072 27492
rect 24673 27489 24685 27523
rect 24719 27520 24731 27523
rect 25774 27520 25780 27532
rect 24719 27492 25780 27520
rect 24719 27489 24731 27492
rect 24673 27483 24731 27489
rect 25774 27480 25780 27492
rect 25832 27480 25838 27532
rect 25884 27520 25912 27560
rect 30466 27548 30472 27560
rect 30524 27548 30530 27600
rect 31726 27588 31754 27628
rect 33870 27588 33876 27600
rect 31726 27560 33876 27588
rect 33870 27548 33876 27560
rect 33928 27548 33934 27600
rect 26237 27523 26295 27529
rect 26237 27520 26249 27523
rect 25884 27492 26249 27520
rect 26237 27489 26249 27492
rect 26283 27489 26295 27523
rect 26694 27520 26700 27532
rect 26655 27492 26700 27520
rect 26237 27483 26295 27489
rect 26694 27480 26700 27492
rect 26752 27520 26758 27532
rect 26752 27492 27200 27520
rect 26752 27480 26758 27492
rect 27172 27452 27200 27492
rect 27246 27480 27252 27532
rect 27304 27520 27310 27532
rect 27801 27523 27859 27529
rect 27801 27520 27813 27523
rect 27304 27492 27813 27520
rect 27304 27480 27310 27492
rect 27801 27489 27813 27492
rect 27847 27489 27859 27523
rect 28166 27520 28172 27532
rect 28127 27492 28172 27520
rect 27801 27483 27859 27489
rect 28166 27480 28172 27492
rect 28224 27520 28230 27532
rect 31754 27520 31760 27532
rect 28224 27492 29592 27520
rect 28224 27480 28230 27492
rect 27338 27452 27344 27464
rect 27172 27424 27344 27452
rect 27338 27412 27344 27424
rect 27396 27412 27402 27464
rect 24670 27384 24676 27396
rect 24044 27356 24676 27384
rect 23661 27347 23719 27353
rect 24670 27344 24676 27356
rect 24728 27344 24734 27396
rect 24762 27344 24768 27396
rect 24820 27384 24826 27396
rect 24820 27356 24865 27384
rect 24820 27344 24826 27356
rect 25314 27344 25320 27396
rect 25372 27384 25378 27396
rect 25685 27387 25743 27393
rect 25685 27384 25697 27387
rect 25372 27356 25697 27384
rect 25372 27344 25378 27356
rect 25685 27353 25697 27356
rect 25731 27353 25743 27387
rect 25685 27347 25743 27353
rect 26329 27387 26387 27393
rect 26329 27353 26341 27387
rect 26375 27384 26387 27387
rect 26418 27384 26424 27396
rect 26375 27356 26424 27384
rect 26375 27353 26387 27356
rect 26329 27347 26387 27353
rect 26418 27344 26424 27356
rect 26476 27344 26482 27396
rect 27890 27344 27896 27396
rect 27948 27384 27954 27396
rect 29564 27384 29592 27492
rect 29748 27492 31760 27520
rect 29748 27464 29776 27492
rect 31754 27480 31760 27492
rect 31812 27480 31818 27532
rect 29730 27452 29736 27464
rect 29691 27424 29736 27452
rect 29730 27412 29736 27424
rect 29788 27412 29794 27464
rect 30374 27452 30380 27464
rect 30335 27424 30380 27452
rect 30374 27412 30380 27424
rect 30432 27412 30438 27464
rect 38286 27452 38292 27464
rect 38247 27424 38292 27452
rect 38286 27412 38292 27424
rect 38344 27412 38350 27464
rect 30466 27384 30472 27396
rect 27948 27356 27993 27384
rect 29564 27356 30472 27384
rect 27948 27344 27954 27356
rect 30466 27344 30472 27356
rect 30524 27344 30530 27396
rect 21928 27288 22876 27316
rect 24394 27276 24400 27328
rect 24452 27316 24458 27328
rect 27706 27316 27712 27328
rect 24452 27288 27712 27316
rect 24452 27276 24458 27288
rect 27706 27276 27712 27288
rect 27764 27276 27770 27328
rect 28074 27276 28080 27328
rect 28132 27316 28138 27328
rect 29825 27319 29883 27325
rect 29825 27316 29837 27319
rect 28132 27288 29837 27316
rect 28132 27276 28138 27288
rect 29825 27285 29837 27288
rect 29871 27285 29883 27319
rect 29825 27279 29883 27285
rect 34514 27276 34520 27328
rect 34572 27316 34578 27328
rect 38105 27319 38163 27325
rect 38105 27316 38117 27319
rect 34572 27288 38117 27316
rect 34572 27276 34578 27288
rect 38105 27285 38117 27288
rect 38151 27285 38163 27319
rect 38105 27279 38163 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1581 27115 1639 27121
rect 1581 27081 1593 27115
rect 1627 27112 1639 27115
rect 8294 27112 8300 27124
rect 1627 27084 8300 27112
rect 1627 27081 1639 27084
rect 1581 27075 1639 27081
rect 8294 27072 8300 27084
rect 8352 27072 8358 27124
rect 9766 27112 9772 27124
rect 9727 27084 9772 27112
rect 9766 27072 9772 27084
rect 9824 27072 9830 27124
rect 10413 27115 10471 27121
rect 10413 27081 10425 27115
rect 10459 27112 10471 27115
rect 10686 27112 10692 27124
rect 10459 27084 10692 27112
rect 10459 27081 10471 27084
rect 10413 27075 10471 27081
rect 10686 27072 10692 27084
rect 10744 27072 10750 27124
rect 11054 27112 11060 27124
rect 11015 27084 11060 27112
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 13924 27084 15056 27112
rect 12250 27044 12256 27056
rect 10336 27016 12256 27044
rect 1762 26976 1768 26988
rect 1723 26948 1768 26976
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 9674 26976 9680 26988
rect 9635 26948 9680 26976
rect 9674 26936 9680 26948
rect 9732 26936 9738 26988
rect 10336 26985 10364 27016
rect 12250 27004 12256 27016
rect 12308 27004 12314 27056
rect 12342 27004 12348 27056
rect 12400 27044 12406 27056
rect 13924 27053 13952 27084
rect 12989 27047 13047 27053
rect 12989 27044 13001 27047
rect 12400 27016 13001 27044
rect 12400 27004 12406 27016
rect 12989 27013 13001 27016
rect 13035 27013 13047 27047
rect 12989 27007 13047 27013
rect 13909 27047 13967 27053
rect 13909 27013 13921 27047
rect 13955 27013 13967 27047
rect 14550 27044 14556 27056
rect 14511 27016 14556 27044
rect 13909 27007 13967 27013
rect 14550 27004 14556 27016
rect 14608 27004 14614 27056
rect 15028 27044 15056 27084
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 20346 27112 20352 27124
rect 15160 27084 20352 27112
rect 15160 27072 15166 27084
rect 20346 27072 20352 27084
rect 20404 27072 20410 27124
rect 26602 27112 26608 27124
rect 22572 27084 26608 27112
rect 15028 27016 16896 27044
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 10686 26936 10692 26988
rect 10744 26976 10750 26988
rect 10870 26976 10876 26988
rect 10744 26948 10876 26976
rect 10744 26936 10750 26948
rect 10870 26936 10876 26948
rect 10928 26976 10934 26988
rect 10965 26979 11023 26985
rect 10965 26976 10977 26979
rect 10928 26948 10977 26976
rect 10928 26936 10934 26948
rect 10965 26945 10977 26948
rect 11011 26945 11023 26979
rect 11885 26979 11943 26985
rect 10965 26939 11023 26945
rect 11256 26948 11836 26976
rect 7374 26868 7380 26920
rect 7432 26908 7438 26920
rect 11256 26908 11284 26948
rect 7432 26880 11284 26908
rect 11701 26911 11759 26917
rect 7432 26868 7438 26880
rect 11701 26877 11713 26911
rect 11747 26877 11759 26911
rect 11808 26908 11836 26948
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12158 26976 12164 26988
rect 11931 26948 12164 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12158 26936 12164 26948
rect 12216 26936 12222 26988
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 14274 26976 14280 26988
rect 14148 26948 14280 26976
rect 14148 26936 14154 26948
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15896 26948 15945 26976
rect 15896 26936 15902 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 11808 26880 12909 26908
rect 11701 26871 11759 26877
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 12897 26871 12955 26877
rect 10778 26732 10784 26784
rect 10836 26772 10842 26784
rect 11716 26772 11744 26871
rect 13998 26868 14004 26920
rect 14056 26908 14062 26920
rect 14461 26911 14519 26917
rect 14461 26908 14473 26911
rect 14056 26880 14473 26908
rect 14056 26868 14062 26880
rect 14461 26877 14473 26880
rect 14507 26908 14519 26911
rect 15010 26908 15016 26920
rect 14507 26880 15016 26908
rect 14507 26877 14519 26880
rect 14461 26871 14519 26877
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 15378 26868 15384 26920
rect 15436 26908 15442 26920
rect 15473 26911 15531 26917
rect 15473 26908 15485 26911
rect 15436 26880 15485 26908
rect 15436 26868 15442 26880
rect 15473 26877 15485 26880
rect 15519 26908 15531 26911
rect 16868 26908 16896 27016
rect 16942 27004 16948 27056
rect 17000 27044 17006 27056
rect 17129 27047 17187 27053
rect 17129 27044 17141 27047
rect 17000 27016 17141 27044
rect 17000 27004 17006 27016
rect 17129 27013 17141 27016
rect 17175 27013 17187 27047
rect 17129 27007 17187 27013
rect 17221 27047 17279 27053
rect 17221 27013 17233 27047
rect 17267 27044 17279 27047
rect 17586 27044 17592 27056
rect 17267 27016 17592 27044
rect 17267 27013 17279 27016
rect 17221 27007 17279 27013
rect 17586 27004 17592 27016
rect 17644 27004 17650 27056
rect 18782 27044 18788 27056
rect 18743 27016 18788 27044
rect 18782 27004 18788 27016
rect 18840 27004 18846 27056
rect 20438 27004 20444 27056
rect 20496 27044 20502 27056
rect 20533 27047 20591 27053
rect 20533 27044 20545 27047
rect 20496 27016 20545 27044
rect 20496 27004 20502 27016
rect 20533 27013 20545 27016
rect 20579 27013 20591 27047
rect 20533 27007 20591 27013
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26976 22063 26979
rect 22370 26976 22376 26988
rect 22051 26948 22376 26976
rect 22051 26945 22063 26948
rect 22005 26939 22063 26945
rect 22370 26936 22376 26948
rect 22428 26936 22434 26988
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 15519 26880 16712 26908
rect 16868 26880 17417 26908
rect 15519 26877 15531 26880
rect 15473 26871 15531 26877
rect 11974 26800 11980 26852
rect 12032 26840 12038 26852
rect 12069 26843 12127 26849
rect 12069 26840 12081 26843
rect 12032 26812 12081 26840
rect 12032 26800 12038 26812
rect 12069 26809 12081 26812
rect 12115 26840 12127 26843
rect 15930 26840 15936 26852
rect 12115 26812 15936 26840
rect 12115 26809 12127 26812
rect 12069 26803 12127 26809
rect 15930 26800 15936 26812
rect 15988 26800 15994 26852
rect 16684 26840 16712 26880
rect 17405 26877 17417 26880
rect 17451 26908 17463 26911
rect 18230 26908 18236 26920
rect 17451 26880 18236 26908
rect 17451 26877 17463 26880
rect 17405 26871 17463 26877
rect 18230 26868 18236 26880
rect 18288 26868 18294 26920
rect 18690 26908 18696 26920
rect 18651 26880 18696 26908
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 20441 26911 20499 26917
rect 20441 26877 20453 26911
rect 20487 26908 20499 26911
rect 20714 26908 20720 26920
rect 20487 26880 20720 26908
rect 20487 26877 20499 26880
rect 20441 26871 20499 26877
rect 20714 26868 20720 26880
rect 20772 26868 20778 26920
rect 20898 26908 20904 26920
rect 20859 26880 20904 26908
rect 20898 26868 20904 26880
rect 20956 26868 20962 26920
rect 22572 26908 22600 27084
rect 26602 27072 26608 27084
rect 26660 27072 26666 27124
rect 29730 27112 29736 27124
rect 27264 27084 29736 27112
rect 22830 27044 22836 27056
rect 22791 27016 22836 27044
rect 22830 27004 22836 27016
rect 22888 27004 22894 27056
rect 24670 27044 24676 27056
rect 24631 27016 24676 27044
rect 24670 27004 24676 27016
rect 24728 27004 24734 27056
rect 24762 27004 24768 27056
rect 24820 27044 24826 27056
rect 26878 27044 26884 27056
rect 24820 27016 26884 27044
rect 24820 27004 24826 27016
rect 26878 27004 26884 27016
rect 26936 27004 26942 27056
rect 27264 27053 27292 27084
rect 29730 27072 29736 27084
rect 29788 27072 29794 27124
rect 33318 27112 33324 27124
rect 33279 27084 33324 27112
rect 33318 27072 33324 27084
rect 33376 27072 33382 27124
rect 27249 27047 27307 27053
rect 27249 27013 27261 27047
rect 27295 27013 27307 27047
rect 27249 27007 27307 27013
rect 27338 27004 27344 27056
rect 27396 27044 27402 27056
rect 28169 27047 28227 27053
rect 27396 27016 27844 27044
rect 27396 27004 27402 27016
rect 26053 26979 26111 26985
rect 26053 26945 26065 26979
rect 26099 26976 26111 26979
rect 26418 26976 26424 26988
rect 26099 26948 26424 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 26418 26936 26424 26948
rect 26476 26976 26482 26988
rect 27430 26976 27436 26988
rect 26476 26948 27436 26976
rect 26476 26936 26482 26948
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 22741 26911 22799 26917
rect 22741 26908 22753 26911
rect 22572 26880 22753 26908
rect 22741 26877 22753 26880
rect 22787 26877 22799 26911
rect 22741 26871 22799 26877
rect 23017 26911 23075 26917
rect 23017 26877 23029 26911
rect 23063 26877 23075 26911
rect 24578 26908 24584 26920
rect 24539 26880 24584 26908
rect 23017 26871 23075 26877
rect 19058 26840 19064 26852
rect 16684 26812 19064 26840
rect 19058 26800 19064 26812
rect 19116 26800 19122 26852
rect 19242 26840 19248 26852
rect 19203 26812 19248 26840
rect 19242 26800 19248 26812
rect 19300 26800 19306 26852
rect 19518 26800 19524 26852
rect 19576 26840 19582 26852
rect 23032 26840 23060 26871
rect 24578 26868 24584 26880
rect 24636 26868 24642 26920
rect 24854 26908 24860 26920
rect 24815 26880 24860 26908
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 27338 26908 27344 26920
rect 24964 26880 27344 26908
rect 19576 26812 23060 26840
rect 19576 26800 19582 26812
rect 24486 26800 24492 26852
rect 24544 26840 24550 26852
rect 24964 26840 24992 26880
rect 27338 26868 27344 26880
rect 27396 26868 27402 26920
rect 24544 26812 24992 26840
rect 24544 26800 24550 26812
rect 27154 26800 27160 26852
rect 27212 26840 27218 26852
rect 27816 26840 27844 27016
rect 28169 27013 28181 27047
rect 28215 27044 28227 27047
rect 29641 27047 29699 27053
rect 29641 27044 29653 27047
rect 28215 27016 29653 27044
rect 28215 27013 28227 27016
rect 28169 27007 28227 27013
rect 29641 27013 29653 27016
rect 29687 27013 29699 27047
rect 29641 27007 29699 27013
rect 29454 26936 29460 26988
rect 29512 26976 29518 26988
rect 29549 26979 29607 26985
rect 29549 26976 29561 26979
rect 29512 26948 29561 26976
rect 29512 26936 29518 26948
rect 29549 26945 29561 26948
rect 29595 26976 29607 26979
rect 30374 26976 30380 26988
rect 29595 26948 30380 26976
rect 29595 26945 29607 26948
rect 29549 26939 29607 26945
rect 30374 26936 30380 26948
rect 30432 26936 30438 26988
rect 32677 26979 32735 26985
rect 32677 26945 32689 26979
rect 32723 26945 32735 26979
rect 32677 26939 32735 26945
rect 33229 26979 33287 26985
rect 33229 26945 33241 26979
rect 33275 26976 33287 26979
rect 33594 26976 33600 26988
rect 33275 26948 33600 26976
rect 33275 26945 33287 26948
rect 33229 26939 33287 26945
rect 28074 26908 28080 26920
rect 28035 26880 28080 26908
rect 28074 26868 28080 26880
rect 28132 26868 28138 26920
rect 28353 26911 28411 26917
rect 28353 26877 28365 26911
rect 28399 26877 28411 26911
rect 28353 26871 28411 26877
rect 28368 26840 28396 26871
rect 31938 26868 31944 26920
rect 31996 26908 32002 26920
rect 32692 26908 32720 26939
rect 33594 26936 33600 26948
rect 33652 26936 33658 26988
rect 38286 26976 38292 26988
rect 38247 26948 38292 26976
rect 38286 26936 38292 26948
rect 38344 26936 38350 26988
rect 34698 26908 34704 26920
rect 31996 26880 34704 26908
rect 31996 26868 32002 26880
rect 34698 26868 34704 26880
rect 34756 26868 34762 26920
rect 27212 26812 27752 26840
rect 27816 26812 28396 26840
rect 32493 26843 32551 26849
rect 27212 26800 27218 26812
rect 14826 26772 14832 26784
rect 10836 26744 14832 26772
rect 10836 26732 10842 26744
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 15838 26732 15844 26784
rect 15896 26772 15902 26784
rect 16025 26775 16083 26781
rect 16025 26772 16037 26775
rect 15896 26744 16037 26772
rect 15896 26732 15902 26744
rect 16025 26741 16037 26744
rect 16071 26741 16083 26775
rect 16025 26735 16083 26741
rect 18046 26732 18052 26784
rect 18104 26772 18110 26784
rect 21174 26772 21180 26784
rect 18104 26744 21180 26772
rect 18104 26732 18110 26744
rect 21174 26732 21180 26744
rect 21232 26732 21238 26784
rect 21358 26732 21364 26784
rect 21416 26772 21422 26784
rect 22097 26775 22155 26781
rect 22097 26772 22109 26775
rect 21416 26744 22109 26772
rect 21416 26732 21422 26744
rect 22097 26741 22109 26744
rect 22143 26741 22155 26775
rect 22097 26735 22155 26741
rect 24762 26732 24768 26784
rect 24820 26772 24826 26784
rect 26145 26775 26203 26781
rect 26145 26772 26157 26775
rect 24820 26744 26157 26772
rect 24820 26732 24826 26744
rect 26145 26741 26157 26744
rect 26191 26741 26203 26775
rect 26145 26735 26203 26741
rect 26786 26732 26792 26784
rect 26844 26772 26850 26784
rect 27341 26775 27399 26781
rect 27341 26772 27353 26775
rect 26844 26744 27353 26772
rect 26844 26732 26850 26744
rect 27341 26741 27353 26744
rect 27387 26741 27399 26775
rect 27724 26772 27752 26812
rect 32493 26809 32505 26843
rect 32539 26840 32551 26843
rect 35342 26840 35348 26852
rect 32539 26812 35348 26840
rect 32539 26809 32551 26812
rect 32493 26803 32551 26809
rect 35342 26800 35348 26812
rect 35400 26800 35406 26852
rect 29362 26772 29368 26784
rect 27724 26744 29368 26772
rect 27341 26735 27399 26741
rect 29362 26732 29368 26744
rect 29420 26772 29426 26784
rect 31294 26772 31300 26784
rect 29420 26744 31300 26772
rect 29420 26732 29426 26744
rect 31294 26732 31300 26744
rect 31352 26732 31358 26784
rect 37274 26732 37280 26784
rect 37332 26772 37338 26784
rect 38105 26775 38163 26781
rect 38105 26772 38117 26775
rect 37332 26744 38117 26772
rect 37332 26732 37338 26744
rect 38105 26741 38117 26744
rect 38151 26741 38163 26775
rect 38105 26735 38163 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 7558 26528 7564 26580
rect 7616 26568 7622 26580
rect 10137 26571 10195 26577
rect 10137 26568 10149 26571
rect 7616 26540 10149 26568
rect 7616 26528 7622 26540
rect 10137 26537 10149 26540
rect 10183 26537 10195 26571
rect 10778 26568 10784 26580
rect 10739 26540 10784 26568
rect 10137 26531 10195 26537
rect 10778 26528 10784 26540
rect 10836 26528 10842 26580
rect 12069 26571 12127 26577
rect 12069 26537 12081 26571
rect 12115 26568 12127 26571
rect 14550 26568 14556 26580
rect 12115 26540 14556 26568
rect 12115 26537 12127 26540
rect 12069 26531 12127 26537
rect 14550 26528 14556 26540
rect 14608 26528 14614 26580
rect 14918 26568 14924 26580
rect 14879 26540 14924 26568
rect 14918 26528 14924 26540
rect 14976 26528 14982 26580
rect 18782 26568 18788 26580
rect 18743 26540 18788 26568
rect 18782 26528 18788 26540
rect 18840 26528 18846 26580
rect 18892 26540 20392 26568
rect 9674 26460 9680 26512
rect 9732 26500 9738 26512
rect 10594 26500 10600 26512
rect 9732 26472 10600 26500
rect 9732 26460 9738 26472
rect 10594 26460 10600 26472
rect 10652 26460 10658 26512
rect 11425 26503 11483 26509
rect 11425 26469 11437 26503
rect 11471 26500 11483 26503
rect 12342 26500 12348 26512
rect 11471 26472 12348 26500
rect 11471 26469 11483 26472
rect 11425 26463 11483 26469
rect 12342 26460 12348 26472
rect 12400 26460 12406 26512
rect 13078 26500 13084 26512
rect 12452 26472 13084 26500
rect 12452 26432 12480 26472
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 15378 26500 15384 26512
rect 13648 26472 15384 26500
rect 12710 26432 12716 26444
rect 10060 26404 12480 26432
rect 12671 26404 12716 26432
rect 10060 26373 10088 26404
rect 12710 26392 12716 26404
rect 12768 26392 12774 26444
rect 12894 26392 12900 26444
rect 12952 26432 12958 26444
rect 12989 26435 13047 26441
rect 12989 26432 13001 26435
rect 12952 26404 13001 26432
rect 12952 26392 12958 26404
rect 12989 26401 13001 26404
rect 13035 26401 13047 26435
rect 13648 26432 13676 26472
rect 15378 26460 15384 26472
rect 15436 26460 15442 26512
rect 15746 26460 15752 26512
rect 15804 26500 15810 26512
rect 16485 26503 16543 26509
rect 16485 26500 16497 26503
rect 15804 26472 16497 26500
rect 15804 26460 15810 26472
rect 16485 26469 16497 26472
rect 16531 26469 16543 26503
rect 16485 26463 16543 26469
rect 17402 26460 17408 26512
rect 17460 26500 17466 26512
rect 18892 26500 18920 26540
rect 17460 26472 18920 26500
rect 17460 26460 17466 26472
rect 19242 26460 19248 26512
rect 19300 26500 19306 26512
rect 20162 26500 20168 26512
rect 19300 26472 20168 26500
rect 19300 26460 19306 26472
rect 20162 26460 20168 26472
rect 20220 26460 20226 26512
rect 12989 26395 13047 26401
rect 13556 26404 13676 26432
rect 10045 26367 10103 26373
rect 10045 26333 10057 26367
rect 10091 26333 10103 26367
rect 10045 26327 10103 26333
rect 10502 26324 10508 26376
rect 10560 26364 10566 26376
rect 10689 26367 10747 26373
rect 10689 26364 10701 26367
rect 10560 26336 10701 26364
rect 10560 26324 10566 26336
rect 10689 26333 10701 26336
rect 10735 26364 10747 26367
rect 10778 26364 10784 26376
rect 10735 26336 10784 26364
rect 10735 26333 10747 26336
rect 10689 26327 10747 26333
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 11330 26364 11336 26376
rect 11291 26336 11336 26364
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 11790 26324 11796 26376
rect 11848 26364 11854 26376
rect 11977 26367 12035 26373
rect 11977 26364 11989 26367
rect 11848 26336 11989 26364
rect 11848 26324 11854 26336
rect 11977 26333 11989 26336
rect 12023 26333 12035 26367
rect 11977 26327 12035 26333
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 12802 26296 12808 26308
rect 8536 26268 12664 26296
rect 12763 26268 12808 26296
rect 8536 26256 8542 26268
rect 12636 26228 12664 26268
rect 12802 26256 12808 26268
rect 12860 26256 12866 26308
rect 13556 26296 13584 26404
rect 14366 26392 14372 26444
rect 14424 26432 14430 26444
rect 14461 26435 14519 26441
rect 14461 26432 14473 26435
rect 14424 26404 14473 26432
rect 14424 26392 14430 26404
rect 14461 26401 14473 26404
rect 14507 26401 14519 26435
rect 14461 26395 14519 26401
rect 15933 26435 15991 26441
rect 15933 26401 15945 26435
rect 15979 26432 15991 26435
rect 15979 26404 16896 26432
rect 15979 26401 15991 26404
rect 15933 26395 15991 26401
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26364 14335 26367
rect 14550 26364 14556 26376
rect 14323 26336 14556 26364
rect 14323 26333 14335 26336
rect 14277 26327 14335 26333
rect 14550 26324 14556 26336
rect 14608 26364 14614 26376
rect 15102 26364 15108 26376
rect 14608 26336 15108 26364
rect 14608 26324 14614 26336
rect 15102 26324 15108 26336
rect 15160 26324 15166 26376
rect 16022 26305 16028 26308
rect 12912 26268 13584 26296
rect 12912 26228 12940 26268
rect 16018 26259 16028 26305
rect 16080 26296 16086 26308
rect 16868 26296 16896 26404
rect 16942 26392 16948 26444
rect 17000 26432 17006 26444
rect 17221 26435 17279 26441
rect 17221 26432 17233 26435
rect 17000 26404 17233 26432
rect 17000 26392 17006 26404
rect 17221 26401 17233 26404
rect 17267 26401 17279 26435
rect 17221 26395 17279 26401
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19797 26435 19855 26441
rect 19797 26432 19809 26435
rect 19392 26404 19809 26432
rect 19392 26392 19398 26404
rect 19797 26401 19809 26404
rect 19843 26432 19855 26435
rect 20070 26432 20076 26444
rect 19843 26404 20076 26432
rect 19843 26401 19855 26404
rect 19797 26395 19855 26401
rect 20070 26392 20076 26404
rect 20128 26392 20134 26444
rect 20364 26432 20392 26540
rect 24670 26528 24676 26580
rect 24728 26568 24734 26580
rect 27801 26571 27859 26577
rect 27801 26568 27813 26571
rect 24728 26540 27813 26568
rect 24728 26528 24734 26540
rect 27801 26537 27813 26540
rect 27847 26537 27859 26571
rect 27801 26531 27859 26537
rect 30466 26528 30472 26580
rect 30524 26568 30530 26580
rect 31386 26568 31392 26580
rect 30524 26540 31392 26568
rect 30524 26528 30530 26540
rect 31386 26528 31392 26540
rect 31444 26528 31450 26580
rect 32677 26571 32735 26577
rect 32677 26537 32689 26571
rect 32723 26568 32735 26571
rect 34606 26568 34612 26580
rect 32723 26540 34612 26568
rect 32723 26537 32735 26540
rect 32677 26531 32735 26537
rect 34606 26528 34612 26540
rect 34664 26528 34670 26580
rect 24946 26460 24952 26512
rect 25004 26500 25010 26512
rect 25225 26503 25283 26509
rect 25225 26500 25237 26503
rect 25004 26472 25237 26500
rect 25004 26460 25010 26472
rect 25225 26469 25237 26472
rect 25271 26469 25283 26503
rect 25225 26463 25283 26469
rect 25314 26460 25320 26512
rect 25372 26500 25378 26512
rect 26142 26500 26148 26512
rect 25372 26472 26148 26500
rect 25372 26460 25378 26472
rect 26142 26460 26148 26472
rect 26200 26460 26206 26512
rect 27246 26500 27252 26512
rect 26252 26472 27252 26500
rect 21269 26435 21327 26441
rect 21269 26432 21281 26435
rect 20364 26404 21281 26432
rect 21269 26401 21281 26404
rect 21315 26401 21327 26435
rect 21269 26395 21327 26401
rect 22833 26435 22891 26441
rect 22833 26401 22845 26435
rect 22879 26432 22891 26435
rect 25774 26432 25780 26444
rect 22879 26404 25780 26432
rect 22879 26401 22891 26404
rect 22833 26395 22891 26401
rect 25774 26392 25780 26404
rect 25832 26392 25838 26444
rect 26252 26441 26280 26472
rect 27246 26460 27252 26472
rect 27304 26460 27310 26512
rect 27338 26460 27344 26512
rect 27396 26500 27402 26512
rect 32033 26503 32091 26509
rect 32033 26500 32045 26503
rect 27396 26472 32045 26500
rect 27396 26460 27402 26472
rect 32033 26469 32045 26472
rect 32079 26469 32091 26503
rect 32033 26463 32091 26469
rect 26237 26435 26295 26441
rect 26237 26401 26249 26435
rect 26283 26401 26295 26435
rect 26237 26395 26295 26401
rect 26326 26392 26332 26444
rect 26384 26432 26390 26444
rect 26513 26435 26571 26441
rect 26513 26432 26525 26435
rect 26384 26404 26525 26432
rect 26384 26392 26390 26404
rect 26513 26401 26525 26404
rect 26559 26401 26571 26435
rect 26513 26395 26571 26401
rect 26694 26392 26700 26444
rect 26752 26432 26758 26444
rect 27062 26432 27068 26444
rect 26752 26404 27068 26432
rect 26752 26392 26758 26404
rect 27062 26392 27068 26404
rect 27120 26392 27126 26444
rect 28445 26435 28503 26441
rect 28445 26432 28457 26435
rect 27172 26404 28457 26432
rect 18598 26324 18604 26376
rect 18656 26364 18662 26376
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18656 26336 18705 26364
rect 18656 26324 18662 26336
rect 18693 26333 18705 26336
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 17218 26296 17224 26308
rect 16080 26268 16118 26296
rect 16868 26268 17224 26296
rect 16022 26256 16028 26259
rect 16080 26256 16086 26268
rect 17218 26256 17224 26268
rect 17276 26256 17282 26308
rect 17310 26256 17316 26308
rect 17368 26296 17374 26308
rect 17368 26268 17413 26296
rect 17368 26256 17374 26268
rect 18046 26256 18052 26308
rect 18104 26296 18110 26308
rect 18233 26299 18291 26305
rect 18233 26296 18245 26299
rect 18104 26268 18245 26296
rect 18104 26256 18110 26268
rect 18233 26265 18245 26268
rect 18279 26265 18291 26299
rect 18233 26259 18291 26265
rect 12636 26200 12940 26228
rect 18708 26228 18736 26327
rect 18782 26256 18788 26308
rect 18840 26296 18846 26308
rect 19518 26296 19524 26308
rect 18840 26268 19524 26296
rect 18840 26256 18846 26268
rect 19518 26256 19524 26268
rect 19576 26256 19582 26308
rect 19613 26299 19671 26305
rect 19613 26265 19625 26299
rect 19659 26296 19671 26299
rect 20162 26296 20168 26308
rect 19659 26268 20168 26296
rect 19659 26265 19671 26268
rect 19613 26259 19671 26265
rect 20162 26256 20168 26268
rect 20220 26256 20226 26308
rect 21358 26256 21364 26308
rect 21416 26296 21422 26308
rect 22281 26299 22339 26305
rect 21416 26268 21461 26296
rect 21416 26256 21422 26268
rect 22281 26265 22293 26299
rect 22327 26296 22339 26299
rect 22830 26296 22836 26308
rect 22327 26268 22836 26296
rect 22327 26265 22339 26268
rect 22281 26259 22339 26265
rect 22830 26256 22836 26268
rect 22888 26256 22894 26308
rect 22922 26256 22928 26308
rect 22980 26296 22986 26308
rect 23845 26299 23903 26305
rect 22980 26268 23025 26296
rect 22980 26256 22986 26268
rect 23845 26265 23857 26299
rect 23891 26296 23903 26299
rect 24118 26296 24124 26308
rect 23891 26268 24124 26296
rect 23891 26265 23903 26268
rect 23845 26259 23903 26265
rect 24118 26256 24124 26268
rect 24176 26256 24182 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 24673 26299 24731 26305
rect 24673 26296 24685 26299
rect 24544 26268 24685 26296
rect 24544 26256 24550 26268
rect 24673 26265 24685 26268
rect 24719 26265 24731 26299
rect 24673 26259 24731 26265
rect 24762 26256 24768 26308
rect 24820 26296 24826 26308
rect 26329 26299 26387 26305
rect 24820 26268 24865 26296
rect 24820 26256 24826 26268
rect 26329 26265 26341 26299
rect 26375 26296 26387 26299
rect 27172 26296 27200 26404
rect 28445 26401 28457 26404
rect 28491 26401 28503 26435
rect 30466 26432 30472 26444
rect 30427 26404 30472 26432
rect 28445 26395 28503 26401
rect 30466 26392 30472 26404
rect 30524 26392 30530 26444
rect 31018 26392 31024 26444
rect 31076 26432 31082 26444
rect 31076 26404 32628 26432
rect 31076 26392 31082 26404
rect 27706 26364 27712 26376
rect 27667 26336 27712 26364
rect 27706 26324 27712 26336
rect 27764 26324 27770 26376
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26333 28411 26367
rect 28353 26327 28411 26333
rect 26375 26268 27200 26296
rect 26375 26265 26387 26268
rect 26329 26259 26387 26265
rect 27430 26256 27436 26308
rect 27488 26296 27494 26308
rect 28368 26296 28396 26327
rect 28534 26324 28540 26376
rect 28592 26364 28598 26376
rect 28997 26367 29055 26373
rect 28997 26364 29009 26367
rect 28592 26336 29009 26364
rect 28592 26324 28598 26336
rect 28997 26333 29009 26336
rect 29043 26333 29055 26367
rect 31294 26364 31300 26376
rect 31255 26336 31300 26364
rect 28997 26327 29055 26333
rect 31294 26324 31300 26336
rect 31352 26324 31358 26376
rect 31938 26364 31944 26376
rect 31899 26336 31944 26364
rect 31938 26324 31944 26336
rect 31996 26324 32002 26376
rect 32600 26373 32628 26404
rect 32585 26367 32643 26373
rect 32585 26333 32597 26367
rect 32631 26333 32643 26367
rect 32585 26327 32643 26333
rect 27488 26268 28396 26296
rect 29089 26299 29147 26305
rect 27488 26256 27494 26268
rect 29089 26265 29101 26299
rect 29135 26296 29147 26299
rect 29822 26296 29828 26308
rect 29135 26268 29684 26296
rect 29783 26268 29828 26296
rect 29135 26265 29147 26268
rect 29089 26259 29147 26265
rect 27154 26228 27160 26240
rect 18708 26200 27160 26228
rect 27154 26188 27160 26200
rect 27212 26188 27218 26240
rect 29656 26228 29684 26268
rect 29822 26256 29828 26268
rect 29880 26256 29886 26308
rect 29917 26299 29975 26305
rect 29917 26265 29929 26299
rect 29963 26265 29975 26299
rect 29917 26259 29975 26265
rect 29932 26228 29960 26259
rect 29656 26200 29960 26228
rect 31389 26231 31447 26237
rect 31389 26197 31401 26231
rect 31435 26228 31447 26231
rect 31570 26228 31576 26240
rect 31435 26200 31576 26228
rect 31435 26197 31447 26200
rect 31389 26191 31447 26197
rect 31570 26188 31576 26200
rect 31628 26188 31634 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 12618 26024 12624 26036
rect 12406 25996 12624 26024
rect 11977 25959 12035 25965
rect 11977 25925 11989 25959
rect 12023 25956 12035 25959
rect 12406 25956 12434 25996
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 12986 25984 12992 26036
rect 13044 26024 13050 26036
rect 16945 26027 17003 26033
rect 13044 25996 15240 26024
rect 13044 25984 13050 25996
rect 12526 25956 12532 25968
rect 12023 25928 12434 25956
rect 12487 25928 12532 25956
rect 12023 25925 12035 25928
rect 11977 25919 12035 25925
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 15102 25956 15108 25968
rect 15063 25928 15108 25956
rect 15102 25916 15108 25928
rect 15160 25916 15166 25968
rect 15212 25956 15240 25996
rect 16945 25993 16957 26027
rect 16991 26024 17003 26027
rect 17310 26024 17316 26036
rect 16991 25996 17316 26024
rect 16991 25993 17003 25996
rect 16945 25987 17003 25993
rect 17310 25984 17316 25996
rect 17368 25984 17374 26036
rect 17586 26024 17592 26036
rect 17547 25996 17592 26024
rect 17586 25984 17592 25996
rect 17644 25984 17650 26036
rect 17678 25984 17684 26036
rect 17736 26024 17742 26036
rect 17736 25996 20208 26024
rect 17736 25984 17742 25996
rect 18877 25959 18935 25965
rect 15212 25928 17540 25956
rect 9861 25891 9919 25897
rect 9861 25857 9873 25891
rect 9907 25857 9919 25891
rect 9861 25851 9919 25857
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25888 10011 25891
rect 10689 25891 10747 25897
rect 10689 25888 10701 25891
rect 9999 25860 10701 25888
rect 9999 25857 10011 25860
rect 9953 25851 10011 25857
rect 10689 25857 10701 25860
rect 10735 25857 10747 25891
rect 13078 25888 13084 25900
rect 13039 25860 13084 25888
rect 10689 25851 10747 25857
rect 9876 25684 9904 25851
rect 13078 25848 13084 25860
rect 13136 25848 13142 25900
rect 13909 25891 13967 25897
rect 13909 25888 13921 25891
rect 13188 25860 13921 25888
rect 10505 25823 10563 25829
rect 10505 25789 10517 25823
rect 10551 25820 10563 25823
rect 10962 25820 10968 25832
rect 10551 25792 10968 25820
rect 10551 25789 10563 25792
rect 10505 25783 10563 25789
rect 10962 25780 10968 25792
rect 11020 25780 11026 25832
rect 11149 25823 11207 25829
rect 11149 25789 11161 25823
rect 11195 25820 11207 25823
rect 11882 25820 11888 25832
rect 11195 25792 11888 25820
rect 11195 25789 11207 25792
rect 11149 25783 11207 25789
rect 11882 25780 11888 25792
rect 11940 25780 11946 25832
rect 13188 25820 13216 25860
rect 13909 25857 13921 25860
rect 13955 25857 13967 25891
rect 13909 25851 13967 25857
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25888 16911 25891
rect 17402 25888 17408 25900
rect 16899 25860 17408 25888
rect 16899 25857 16911 25860
rect 16853 25851 16911 25857
rect 17402 25848 17408 25860
rect 17460 25848 17466 25900
rect 17512 25897 17540 25928
rect 18877 25925 18889 25959
rect 18923 25956 18935 25959
rect 20070 25956 20076 25968
rect 18923 25928 20076 25956
rect 18923 25925 18935 25928
rect 18877 25919 18935 25925
rect 20070 25916 20076 25928
rect 20128 25916 20134 25968
rect 17497 25891 17555 25897
rect 17497 25857 17509 25891
rect 17543 25857 17555 25891
rect 17497 25851 17555 25857
rect 12406 25792 13216 25820
rect 13725 25823 13783 25829
rect 10870 25712 10876 25764
rect 10928 25752 10934 25764
rect 12406 25752 12434 25792
rect 13725 25789 13737 25823
rect 13771 25820 13783 25823
rect 14550 25820 14556 25832
rect 13771 25792 14556 25820
rect 13771 25789 13783 25792
rect 13725 25783 13783 25789
rect 14550 25780 14556 25792
rect 14608 25780 14614 25832
rect 15010 25820 15016 25832
rect 14923 25792 15016 25820
rect 15010 25780 15016 25792
rect 15068 25780 15074 25832
rect 15654 25820 15660 25832
rect 15615 25792 15660 25820
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 10928 25724 12434 25752
rect 13173 25755 13231 25761
rect 10928 25712 10934 25724
rect 13173 25721 13185 25755
rect 13219 25752 13231 25755
rect 14458 25752 14464 25764
rect 13219 25724 14464 25752
rect 13219 25721 13231 25724
rect 13173 25715 13231 25721
rect 14458 25712 14464 25724
rect 14516 25712 14522 25764
rect 15028 25752 15056 25780
rect 17126 25752 17132 25764
rect 15028 25724 17132 25752
rect 17126 25712 17132 25724
rect 17184 25712 17190 25764
rect 17512 25752 17540 25851
rect 18785 25823 18843 25829
rect 18785 25789 18797 25823
rect 18831 25820 18843 25823
rect 19242 25820 19248 25832
rect 18831 25792 19248 25820
rect 18831 25789 18843 25792
rect 18785 25783 18843 25789
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 19797 25823 19855 25829
rect 19797 25789 19809 25823
rect 19843 25820 19855 25823
rect 20180 25820 20208 25996
rect 20806 25984 20812 26036
rect 20864 26024 20870 26036
rect 22002 26024 22008 26036
rect 20864 25996 22008 26024
rect 20864 25984 20870 25996
rect 22002 25984 22008 25996
rect 22060 25984 22066 26036
rect 22112 25996 27476 26024
rect 21269 25891 21327 25897
rect 21269 25857 21281 25891
rect 21315 25888 21327 25891
rect 21818 25888 21824 25900
rect 21315 25860 21824 25888
rect 21315 25857 21327 25860
rect 21269 25851 21327 25857
rect 20806 25820 20812 25832
rect 19843 25792 20812 25820
rect 19843 25789 19855 25792
rect 19797 25783 19855 25789
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 21284 25752 21312 25851
rect 21818 25848 21824 25860
rect 21876 25848 21882 25900
rect 22112 25897 22140 25996
rect 23106 25956 23112 25968
rect 23067 25928 23112 25956
rect 23106 25916 23112 25928
rect 23164 25916 23170 25968
rect 24578 25956 24584 25968
rect 24539 25928 24584 25956
rect 24578 25916 24584 25928
rect 24636 25916 24642 25968
rect 24673 25959 24731 25965
rect 24673 25925 24685 25959
rect 24719 25956 24731 25959
rect 26142 25956 26148 25968
rect 24719 25928 26148 25956
rect 24719 25925 24731 25928
rect 24673 25919 24731 25925
rect 26142 25916 26148 25928
rect 26200 25916 26206 25968
rect 26421 25959 26479 25965
rect 26421 25956 26433 25959
rect 26252 25928 26433 25956
rect 22097 25891 22155 25897
rect 22097 25857 22109 25891
rect 22143 25857 22155 25891
rect 25682 25888 25688 25900
rect 25643 25860 25688 25888
rect 22097 25851 22155 25857
rect 25682 25848 25688 25860
rect 25740 25848 25746 25900
rect 26252 25888 26280 25928
rect 26421 25925 26433 25928
rect 26467 25925 26479 25959
rect 27448 25956 27476 25996
rect 27522 25984 27528 26036
rect 27580 26024 27586 26036
rect 27801 26027 27859 26033
rect 27801 26024 27813 26027
rect 27580 25996 27813 26024
rect 27580 25984 27586 25996
rect 27801 25993 27813 25996
rect 27847 25993 27859 26027
rect 30745 26027 30803 26033
rect 30745 26024 30757 26027
rect 27801 25987 27859 25993
rect 29288 25996 30757 26024
rect 28902 25956 28908 25968
rect 27448 25928 28908 25956
rect 26421 25919 26479 25925
rect 28902 25916 28908 25928
rect 28960 25916 28966 25968
rect 29288 25965 29316 25996
rect 30745 25993 30757 25996
rect 30791 25993 30803 26027
rect 30745 25987 30803 25993
rect 31389 26027 31447 26033
rect 31389 25993 31401 26027
rect 31435 26024 31447 26027
rect 38010 26024 38016 26036
rect 31435 25996 38016 26024
rect 31435 25993 31447 25996
rect 31389 25987 31447 25993
rect 38010 25984 38016 25996
rect 38068 25984 38074 26036
rect 29273 25959 29331 25965
rect 29273 25925 29285 25959
rect 29319 25925 29331 25959
rect 29273 25919 29331 25925
rect 29365 25959 29423 25965
rect 29365 25925 29377 25959
rect 29411 25956 29423 25959
rect 29730 25956 29736 25968
rect 29411 25928 29736 25956
rect 29411 25925 29423 25928
rect 29365 25919 29423 25925
rect 29730 25916 29736 25928
rect 29788 25916 29794 25968
rect 30098 25916 30104 25968
rect 30156 25956 30162 25968
rect 38194 25956 38200 25968
rect 30156 25928 38200 25956
rect 30156 25916 30162 25928
rect 38194 25916 38200 25928
rect 38252 25916 38258 25968
rect 25792 25860 26280 25888
rect 26329 25891 26387 25897
rect 23017 25823 23075 25829
rect 23017 25789 23029 25823
rect 23063 25820 23075 25823
rect 23382 25820 23388 25832
rect 23063 25792 23388 25820
rect 23063 25789 23075 25792
rect 23017 25783 23075 25789
rect 23382 25780 23388 25792
rect 23440 25780 23446 25832
rect 24026 25820 24032 25832
rect 23987 25792 24032 25820
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 24946 25820 24952 25832
rect 24907 25792 24952 25820
rect 24946 25780 24952 25792
rect 25004 25780 25010 25832
rect 25498 25820 25504 25832
rect 25056 25792 25504 25820
rect 17512 25724 21312 25752
rect 21361 25755 21419 25761
rect 21361 25721 21373 25755
rect 21407 25752 21419 25755
rect 22922 25752 22928 25764
rect 21407 25724 22928 25752
rect 21407 25721 21419 25724
rect 21361 25715 21419 25721
rect 22922 25712 22928 25724
rect 22980 25712 22986 25764
rect 23106 25712 23112 25764
rect 23164 25752 23170 25764
rect 25056 25752 25084 25792
rect 25498 25780 25504 25792
rect 25556 25820 25562 25832
rect 25792 25820 25820 25860
rect 26329 25857 26341 25891
rect 26375 25857 26387 25891
rect 27154 25888 27160 25900
rect 27115 25860 27160 25888
rect 26329 25851 26387 25857
rect 25556 25792 25820 25820
rect 26344 25820 26372 25851
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 27985 25891 28043 25897
rect 27985 25857 27997 25891
rect 28031 25857 28043 25891
rect 28534 25888 28540 25900
rect 28495 25860 28540 25888
rect 27985 25851 28043 25857
rect 28000 25820 28028 25851
rect 28534 25848 28540 25860
rect 28592 25848 28598 25900
rect 30190 25848 30196 25900
rect 30248 25888 30254 25900
rect 31573 25891 31631 25897
rect 31573 25888 31585 25891
rect 30248 25860 31585 25888
rect 30248 25848 30254 25860
rect 31573 25857 31585 25860
rect 31619 25857 31631 25891
rect 31573 25851 31631 25857
rect 34149 25891 34207 25897
rect 34149 25857 34161 25891
rect 34195 25888 34207 25891
rect 34514 25888 34520 25900
rect 34195 25860 34520 25888
rect 34195 25857 34207 25860
rect 34149 25851 34207 25857
rect 34514 25848 34520 25860
rect 34572 25848 34578 25900
rect 30282 25820 30288 25832
rect 26344 25792 30052 25820
rect 30243 25792 30288 25820
rect 25556 25780 25562 25792
rect 27249 25755 27307 25761
rect 23164 25724 25084 25752
rect 25332 25724 27200 25752
rect 23164 25712 23170 25724
rect 25332 25696 25360 25724
rect 11146 25684 11152 25696
rect 9876 25656 11152 25684
rect 11146 25644 11152 25656
rect 11204 25684 11210 25696
rect 12342 25684 12348 25696
rect 11204 25656 12348 25684
rect 11204 25644 11210 25656
rect 12342 25644 12348 25656
rect 12400 25644 12406 25696
rect 13722 25644 13728 25696
rect 13780 25684 13786 25696
rect 14093 25687 14151 25693
rect 14093 25684 14105 25687
rect 13780 25656 14105 25684
rect 13780 25644 13786 25656
rect 14093 25653 14105 25656
rect 14139 25653 14151 25687
rect 14093 25647 14151 25653
rect 16114 25644 16120 25696
rect 16172 25684 16178 25696
rect 21082 25684 21088 25696
rect 16172 25656 21088 25684
rect 16172 25644 16178 25656
rect 21082 25644 21088 25656
rect 21140 25644 21146 25696
rect 21450 25644 21456 25696
rect 21508 25684 21514 25696
rect 22189 25687 22247 25693
rect 22189 25684 22201 25687
rect 21508 25656 22201 25684
rect 21508 25644 21514 25656
rect 22189 25653 22201 25656
rect 22235 25653 22247 25687
rect 22189 25647 22247 25653
rect 24946 25644 24952 25696
rect 25004 25684 25010 25696
rect 25314 25684 25320 25696
rect 25004 25656 25320 25684
rect 25004 25644 25010 25656
rect 25314 25644 25320 25656
rect 25372 25644 25378 25696
rect 25774 25684 25780 25696
rect 25735 25656 25780 25684
rect 25774 25644 25780 25656
rect 25832 25644 25838 25696
rect 27172 25684 27200 25724
rect 27249 25721 27261 25755
rect 27295 25752 27307 25755
rect 29914 25752 29920 25764
rect 27295 25724 29920 25752
rect 27295 25721 27307 25724
rect 27249 25715 27307 25721
rect 29914 25712 29920 25724
rect 29972 25712 29978 25764
rect 30024 25752 30052 25792
rect 30282 25780 30288 25792
rect 30340 25780 30346 25832
rect 34422 25752 34428 25764
rect 30024 25724 34428 25752
rect 34422 25712 34428 25724
rect 34480 25712 34486 25764
rect 28442 25684 28448 25696
rect 27172 25656 28448 25684
rect 28442 25644 28448 25656
rect 28500 25644 28506 25696
rect 28629 25687 28687 25693
rect 28629 25653 28641 25687
rect 28675 25684 28687 25687
rect 28810 25684 28816 25696
rect 28675 25656 28816 25684
rect 28675 25653 28687 25656
rect 28629 25647 28687 25653
rect 28810 25644 28816 25656
rect 28868 25644 28874 25696
rect 28902 25644 28908 25696
rect 28960 25684 28966 25696
rect 31846 25684 31852 25696
rect 28960 25656 31852 25684
rect 28960 25644 28966 25656
rect 31846 25644 31852 25656
rect 31904 25644 31910 25696
rect 33686 25644 33692 25696
rect 33744 25684 33750 25696
rect 34241 25687 34299 25693
rect 34241 25684 34253 25687
rect 33744 25656 34253 25684
rect 33744 25644 33750 25656
rect 34241 25653 34253 25656
rect 34287 25653 34299 25687
rect 34241 25647 34299 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 10870 25480 10876 25492
rect 10831 25452 10876 25480
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 11882 25440 11888 25492
rect 11940 25480 11946 25492
rect 13722 25480 13728 25492
rect 11940 25452 13728 25480
rect 11940 25440 11946 25452
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 14090 25440 14096 25492
rect 14148 25480 14154 25492
rect 30190 25480 30196 25492
rect 14148 25452 30196 25480
rect 14148 25440 14154 25452
rect 30190 25440 30196 25452
rect 30248 25440 30254 25492
rect 2746 25384 12434 25412
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25276 1639 25279
rect 2746 25276 2774 25384
rect 9585 25347 9643 25353
rect 9585 25313 9597 25347
rect 9631 25344 9643 25347
rect 11609 25347 11667 25353
rect 11609 25344 11621 25347
rect 9631 25316 11621 25344
rect 9631 25313 9643 25316
rect 9585 25307 9643 25313
rect 11609 25313 11621 25316
rect 11655 25313 11667 25347
rect 11609 25307 11667 25313
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 12069 25347 12127 25353
rect 12069 25344 12081 25347
rect 12032 25316 12081 25344
rect 12032 25304 12038 25316
rect 12069 25313 12081 25316
rect 12115 25313 12127 25347
rect 12406 25344 12434 25384
rect 14182 25372 14188 25424
rect 14240 25412 14246 25424
rect 16850 25412 16856 25424
rect 14240 25384 16856 25412
rect 14240 25372 14246 25384
rect 16850 25372 16856 25384
rect 16908 25372 16914 25424
rect 25682 25412 25688 25424
rect 18432 25384 25688 25412
rect 12406 25316 18000 25344
rect 12069 25307 12127 25313
rect 9490 25276 9496 25288
rect 1627 25248 2774 25276
rect 9451 25248 9496 25276
rect 1627 25245 1639 25248
rect 1581 25239 1639 25245
rect 9490 25236 9496 25248
rect 9548 25236 9554 25288
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 10152 25208 10180 25239
rect 10686 25236 10692 25288
rect 10744 25276 10750 25288
rect 10781 25279 10839 25285
rect 10781 25276 10793 25279
rect 10744 25248 10793 25276
rect 10744 25236 10750 25248
rect 10781 25245 10793 25248
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 10962 25236 10968 25288
rect 11020 25276 11026 25288
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 11020 25248 11437 25276
rect 11020 25236 11026 25248
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25245 13139 25279
rect 13262 25276 13268 25288
rect 13223 25248 13268 25276
rect 13081 25239 13139 25245
rect 10152 25180 12204 25208
rect 1762 25140 1768 25152
rect 1723 25112 1768 25140
rect 1762 25100 1768 25112
rect 1820 25100 1826 25152
rect 5994 25100 6000 25152
rect 6052 25140 6058 25152
rect 9858 25140 9864 25152
rect 6052 25112 9864 25140
rect 6052 25100 6058 25112
rect 9858 25100 9864 25112
rect 9916 25100 9922 25152
rect 10229 25143 10287 25149
rect 10229 25109 10241 25143
rect 10275 25140 10287 25143
rect 11974 25140 11980 25152
rect 10275 25112 11980 25140
rect 10275 25109 10287 25112
rect 10229 25103 10287 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12176 25140 12204 25180
rect 12986 25140 12992 25152
rect 12176 25112 12992 25140
rect 12986 25100 12992 25112
rect 13044 25100 13050 25152
rect 13096 25140 13124 25239
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 16114 25276 16120 25288
rect 16075 25248 16120 25276
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 14182 25168 14188 25220
rect 14240 25208 14246 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 14240 25180 14381 25208
rect 14240 25168 14246 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 14458 25168 14464 25220
rect 14516 25208 14522 25220
rect 15381 25211 15439 25217
rect 14516 25180 14561 25208
rect 14516 25168 14522 25180
rect 15381 25177 15393 25211
rect 15427 25208 15439 25211
rect 16574 25208 16580 25220
rect 15427 25180 16580 25208
rect 15427 25177 15439 25180
rect 15381 25171 15439 25177
rect 16574 25168 16580 25180
rect 16632 25168 16638 25220
rect 16850 25208 16856 25220
rect 16811 25180 16856 25208
rect 16850 25168 16856 25180
rect 16908 25168 16914 25220
rect 16945 25211 17003 25217
rect 16945 25177 16957 25211
rect 16991 25177 17003 25211
rect 16945 25171 17003 25177
rect 15746 25140 15752 25152
rect 13096 25112 15752 25140
rect 15746 25100 15752 25112
rect 15804 25100 15810 25152
rect 16022 25100 16028 25152
rect 16080 25140 16086 25152
rect 16209 25143 16267 25149
rect 16209 25140 16221 25143
rect 16080 25112 16221 25140
rect 16080 25100 16086 25112
rect 16209 25109 16221 25112
rect 16255 25109 16267 25143
rect 16960 25140 16988 25171
rect 17034 25168 17040 25220
rect 17092 25208 17098 25220
rect 17865 25211 17923 25217
rect 17865 25208 17877 25211
rect 17092 25180 17877 25208
rect 17092 25168 17098 25180
rect 17865 25177 17877 25180
rect 17911 25177 17923 25211
rect 17972 25208 18000 25316
rect 18432 25285 18460 25384
rect 25682 25372 25688 25384
rect 25740 25412 25746 25424
rect 37642 25412 37648 25424
rect 25740 25384 37648 25412
rect 25740 25372 25746 25384
rect 37642 25372 37648 25384
rect 37700 25372 37706 25424
rect 24857 25347 24915 25353
rect 24857 25344 24869 25347
rect 18524 25316 24869 25344
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18524 25208 18552 25316
rect 24857 25313 24869 25316
rect 24903 25313 24915 25347
rect 24857 25307 24915 25313
rect 25409 25347 25467 25353
rect 25409 25313 25421 25347
rect 25455 25344 25467 25347
rect 26973 25347 27031 25353
rect 25455 25316 26832 25344
rect 25455 25313 25467 25316
rect 25409 25307 25467 25313
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25276 20039 25279
rect 20254 25276 20260 25288
rect 20027 25248 20260 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20254 25236 20260 25248
rect 20312 25236 20318 25288
rect 20622 25276 20628 25288
rect 20583 25248 20628 25276
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 24210 25236 24216 25288
rect 24268 25276 24274 25288
rect 24762 25276 24768 25288
rect 24268 25248 24768 25276
rect 24268 25236 24274 25248
rect 24762 25236 24768 25248
rect 24820 25236 24826 25288
rect 17972 25180 18552 25208
rect 20073 25211 20131 25217
rect 17865 25171 17923 25177
rect 20073 25177 20085 25211
rect 20119 25208 20131 25211
rect 20530 25208 20536 25220
rect 20119 25180 20536 25208
rect 20119 25177 20131 25180
rect 20073 25171 20131 25177
rect 20530 25168 20536 25180
rect 20588 25208 20594 25220
rect 21361 25211 21419 25217
rect 21361 25208 21373 25211
rect 20588 25180 21373 25208
rect 20588 25168 20594 25180
rect 21361 25177 21373 25180
rect 21407 25177 21419 25211
rect 21361 25171 21419 25177
rect 21450 25168 21456 25220
rect 21508 25208 21514 25220
rect 22002 25208 22008 25220
rect 21508 25180 21553 25208
rect 21963 25180 22008 25208
rect 21508 25168 21514 25180
rect 22002 25168 22008 25180
rect 22060 25208 22066 25220
rect 22741 25211 22799 25217
rect 22741 25208 22753 25211
rect 22060 25180 22753 25208
rect 22060 25168 22066 25180
rect 22741 25177 22753 25180
rect 22787 25177 22799 25211
rect 22741 25171 22799 25177
rect 22833 25211 22891 25217
rect 22833 25177 22845 25211
rect 22879 25208 22891 25211
rect 23566 25208 23572 25220
rect 22879 25180 23572 25208
rect 22879 25177 22891 25180
rect 22833 25171 22891 25177
rect 23566 25168 23572 25180
rect 23624 25168 23630 25220
rect 23753 25211 23811 25217
rect 23753 25177 23765 25211
rect 23799 25208 23811 25211
rect 24578 25208 24584 25220
rect 23799 25180 24584 25208
rect 23799 25177 23811 25180
rect 23753 25171 23811 25177
rect 24578 25168 24584 25180
rect 24636 25168 24642 25220
rect 24673 25211 24731 25217
rect 24673 25177 24685 25211
rect 24719 25177 24731 25211
rect 24673 25171 24731 25177
rect 18322 25140 18328 25152
rect 16960 25112 18328 25140
rect 16209 25103 16267 25109
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 18506 25140 18512 25152
rect 18467 25112 18512 25140
rect 18506 25100 18512 25112
rect 18564 25100 18570 25152
rect 20717 25143 20775 25149
rect 20717 25109 20729 25143
rect 20763 25140 20775 25143
rect 21174 25140 21180 25152
rect 20763 25112 21180 25140
rect 20763 25109 20775 25112
rect 20717 25103 20775 25109
rect 21174 25100 21180 25112
rect 21232 25100 21238 25152
rect 24688 25140 24716 25171
rect 25498 25168 25504 25220
rect 25556 25208 25562 25220
rect 26421 25211 26479 25217
rect 25556 25180 25601 25208
rect 25556 25168 25562 25180
rect 26421 25177 26433 25211
rect 26467 25208 26479 25211
rect 26694 25208 26700 25220
rect 26467 25180 26700 25208
rect 26467 25177 26479 25180
rect 26421 25171 26479 25177
rect 26694 25168 26700 25180
rect 26752 25168 26758 25220
rect 26510 25140 26516 25152
rect 24688 25112 26516 25140
rect 26510 25100 26516 25112
rect 26568 25100 26574 25152
rect 26804 25140 26832 25316
rect 26973 25313 26985 25347
rect 27019 25344 27031 25347
rect 27246 25344 27252 25356
rect 27019 25316 27252 25344
rect 27019 25313 27031 25316
rect 26973 25307 27031 25313
rect 27246 25304 27252 25316
rect 27304 25304 27310 25356
rect 27614 25344 27620 25356
rect 27575 25316 27620 25344
rect 27614 25304 27620 25316
rect 27672 25304 27678 25356
rect 28534 25304 28540 25356
rect 28592 25344 28598 25356
rect 30098 25344 30104 25356
rect 28592 25316 30104 25344
rect 28592 25304 28598 25316
rect 30098 25304 30104 25316
rect 30156 25304 30162 25356
rect 31754 25344 31760 25356
rect 31715 25316 31760 25344
rect 31754 25304 31760 25316
rect 31812 25304 31818 25356
rect 33686 25344 33692 25356
rect 33647 25316 33692 25344
rect 33686 25304 33692 25316
rect 33744 25304 33750 25356
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 27065 25211 27123 25217
rect 27065 25177 27077 25211
rect 27111 25208 27123 25211
rect 27798 25208 27804 25220
rect 27111 25180 27804 25208
rect 27111 25177 27123 25180
rect 27065 25171 27123 25177
rect 27798 25168 27804 25180
rect 27856 25168 27862 25220
rect 28810 25168 28816 25220
rect 28868 25208 28874 25220
rect 29822 25208 29828 25220
rect 28868 25180 29828 25208
rect 28868 25168 28874 25180
rect 29822 25168 29828 25180
rect 29880 25168 29886 25220
rect 29914 25168 29920 25220
rect 29972 25208 29978 25220
rect 30837 25211 30895 25217
rect 29972 25180 30017 25208
rect 29972 25168 29978 25180
rect 30837 25177 30849 25211
rect 30883 25177 30895 25211
rect 31478 25208 31484 25220
rect 31439 25180 31484 25208
rect 30837 25171 30895 25177
rect 28074 25140 28080 25152
rect 26804 25112 28080 25140
rect 28074 25100 28080 25112
rect 28132 25100 28138 25152
rect 28442 25100 28448 25152
rect 28500 25140 28506 25152
rect 30852 25140 30880 25171
rect 31478 25168 31484 25180
rect 31536 25168 31542 25220
rect 31570 25168 31576 25220
rect 31628 25208 31634 25220
rect 33778 25208 33784 25220
rect 31628 25180 31673 25208
rect 33739 25180 33784 25208
rect 31628 25168 31634 25180
rect 33778 25168 33784 25180
rect 33836 25168 33842 25220
rect 34333 25211 34391 25217
rect 34333 25177 34345 25211
rect 34379 25177 34391 25211
rect 34333 25171 34391 25177
rect 30926 25140 30932 25152
rect 28500 25112 30932 25140
rect 28500 25100 28506 25112
rect 30926 25100 30932 25112
rect 30984 25100 30990 25152
rect 33410 25100 33416 25152
rect 33468 25140 33474 25152
rect 33962 25140 33968 25152
rect 33468 25112 33968 25140
rect 33468 25100 33474 25112
rect 33962 25100 33968 25112
rect 34020 25140 34026 25152
rect 34348 25140 34376 25171
rect 34422 25168 34428 25220
rect 34480 25208 34486 25220
rect 38654 25208 38660 25220
rect 34480 25180 38660 25208
rect 34480 25168 34486 25180
rect 38654 25168 38660 25180
rect 38712 25168 38718 25220
rect 38194 25140 38200 25152
rect 34020 25112 34376 25140
rect 38155 25112 38200 25140
rect 34020 25100 34026 25112
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7282 24896 7288 24948
rect 7340 24936 7346 24948
rect 10686 24936 10692 24948
rect 7340 24908 10692 24936
rect 7340 24896 7346 24908
rect 10686 24896 10692 24908
rect 10744 24896 10750 24948
rect 16482 24936 16488 24948
rect 13280 24908 16488 24936
rect 9493 24871 9551 24877
rect 9493 24837 9505 24871
rect 9539 24868 9551 24871
rect 9674 24868 9680 24880
rect 9539 24840 9680 24868
rect 9539 24837 9551 24840
rect 9493 24831 9551 24837
rect 9674 24828 9680 24840
rect 9732 24828 9738 24880
rect 12158 24868 12164 24880
rect 10888 24840 11100 24868
rect 12119 24840 12164 24868
rect 1762 24800 1768 24812
rect 1723 24772 1768 24800
rect 1762 24760 1768 24772
rect 1820 24760 1826 24812
rect 10888 24800 10916 24840
rect 10244 24772 10916 24800
rect 10965 24803 11023 24809
rect 9398 24732 9404 24744
rect 9359 24704 9404 24732
rect 9398 24692 9404 24704
rect 9456 24692 9462 24744
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 9677 24735 9735 24741
rect 9677 24732 9689 24735
rect 9640 24704 9689 24732
rect 9640 24692 9646 24704
rect 9677 24701 9689 24704
rect 9723 24701 9735 24735
rect 9677 24695 9735 24701
rect 8202 24624 8208 24676
rect 8260 24664 8266 24676
rect 10244 24664 10272 24772
rect 10965 24769 10977 24803
rect 11011 24769 11023 24803
rect 11072 24800 11100 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 12544 24840 12848 24868
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11072 24772 12081 24800
rect 10965 24763 11023 24769
rect 12069 24769 12081 24772
rect 12115 24800 12127 24803
rect 12544 24800 12572 24840
rect 12710 24800 12716 24812
rect 12115 24772 12572 24800
rect 12671 24772 12716 24800
rect 12115 24769 12127 24772
rect 12069 24763 12127 24769
rect 10594 24692 10600 24744
rect 10652 24732 10658 24744
rect 10980 24732 11008 24763
rect 12710 24760 12716 24772
rect 12768 24760 12774 24812
rect 12820 24800 12848 24840
rect 13280 24800 13308 24908
rect 16482 24896 16488 24908
rect 16540 24896 16546 24948
rect 26694 24936 26700 24948
rect 16592 24908 17816 24936
rect 15120 24840 15332 24868
rect 12820 24772 13308 24800
rect 13357 24803 13415 24809
rect 13357 24769 13369 24803
rect 13403 24800 13415 24803
rect 13446 24800 13452 24812
rect 13403 24772 13452 24800
rect 13403 24769 13415 24772
rect 13357 24763 13415 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 13998 24760 14004 24812
rect 14056 24800 14062 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 14056 24772 14565 24800
rect 14056 24760 14062 24772
rect 14553 24769 14565 24772
rect 14599 24800 14611 24803
rect 15120 24800 15148 24840
rect 14599 24772 15148 24800
rect 15197 24803 15255 24809
rect 14599 24769 14611 24772
rect 14553 24763 14611 24769
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 10652 24704 11008 24732
rect 11057 24735 11115 24741
rect 10652 24692 10658 24704
rect 11057 24701 11069 24735
rect 11103 24701 11115 24735
rect 13262 24732 13268 24744
rect 11057 24695 11115 24701
rect 12406 24704 13268 24732
rect 8260 24636 10272 24664
rect 11072 24664 11100 24695
rect 12406 24664 12434 24704
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 11072 24636 12434 24664
rect 12805 24667 12863 24673
rect 8260 24624 8266 24636
rect 12805 24633 12817 24667
rect 12851 24664 12863 24667
rect 15102 24664 15108 24676
rect 12851 24636 15108 24664
rect 12851 24633 12863 24636
rect 12805 24627 12863 24633
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 15212 24664 15240 24763
rect 15304 24732 15332 24840
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 16117 24803 16175 24809
rect 16117 24800 16129 24803
rect 15436 24772 16129 24800
rect 15436 24760 15442 24772
rect 16117 24769 16129 24772
rect 16163 24800 16175 24803
rect 16592 24800 16620 24908
rect 17037 24871 17095 24877
rect 17037 24868 17049 24871
rect 16776 24840 17049 24868
rect 16163 24772 16620 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 16776 24800 16804 24840
rect 17037 24837 17049 24840
rect 17083 24837 17095 24871
rect 17037 24831 17095 24837
rect 16724 24772 16804 24800
rect 17788 24800 17816 24908
rect 22066 24908 26700 24936
rect 19981 24871 20039 24877
rect 19981 24868 19993 24871
rect 18248 24840 18552 24868
rect 18248 24800 18276 24840
rect 18414 24800 18420 24812
rect 17788 24772 18276 24800
rect 18375 24772 18420 24800
rect 16724 24760 16730 24772
rect 18414 24760 18420 24772
rect 18472 24760 18478 24812
rect 18524 24800 18552 24840
rect 19720 24840 19993 24868
rect 19150 24800 19156 24812
rect 18524 24772 18644 24800
rect 19111 24772 19156 24800
rect 16758 24732 16764 24744
rect 15304 24704 16764 24732
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 16945 24735 17003 24741
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 17126 24732 17132 24744
rect 16991 24704 17132 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 17310 24732 17316 24744
rect 17271 24704 17316 24732
rect 17310 24692 17316 24704
rect 17368 24732 17374 24744
rect 17586 24732 17592 24744
rect 17368 24704 17592 24732
rect 17368 24692 17374 24704
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 18322 24692 18328 24744
rect 18380 24732 18386 24744
rect 18509 24735 18567 24741
rect 18509 24732 18521 24735
rect 18380 24704 18521 24732
rect 18380 24692 18386 24704
rect 18509 24701 18521 24704
rect 18555 24701 18567 24735
rect 18616 24732 18644 24772
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19720 24800 19748 24840
rect 19981 24837 19993 24840
rect 20027 24837 20039 24871
rect 20898 24868 20904 24880
rect 20859 24840 20904 24868
rect 19981 24831 20039 24837
rect 20898 24828 20904 24840
rect 20956 24868 20962 24880
rect 22066 24868 22094 24908
rect 26694 24896 26700 24908
rect 26752 24936 26758 24948
rect 27890 24936 27896 24948
rect 26752 24908 27896 24936
rect 26752 24896 26758 24908
rect 27890 24896 27896 24908
rect 27948 24896 27954 24948
rect 20956 24840 22094 24868
rect 22649 24871 22707 24877
rect 20956 24828 20962 24840
rect 22649 24837 22661 24871
rect 22695 24868 22707 24871
rect 24210 24868 24216 24880
rect 22695 24840 23428 24868
rect 24171 24840 24216 24868
rect 22695 24837 22707 24840
rect 22649 24831 22707 24837
rect 19291 24772 19748 24800
rect 23400 24800 23428 24840
rect 24210 24828 24216 24840
rect 24268 24828 24274 24880
rect 27341 24871 27399 24877
rect 27341 24868 27353 24871
rect 27172 24840 27353 24868
rect 23934 24800 23940 24812
rect 23400 24772 23940 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 25406 24800 25412 24812
rect 25148 24772 25412 24800
rect 19889 24735 19947 24741
rect 18616 24704 19840 24732
rect 18509 24695 18567 24701
rect 19702 24664 19708 24676
rect 15212 24636 19708 24664
rect 19702 24624 19708 24636
rect 19760 24624 19766 24676
rect 19812 24664 19840 24704
rect 19889 24701 19901 24735
rect 19935 24732 19947 24735
rect 20714 24732 20720 24744
rect 19935 24704 20720 24732
rect 19935 24701 19947 24704
rect 19889 24695 19947 24701
rect 20714 24692 20720 24704
rect 20772 24732 20778 24744
rect 22557 24735 22615 24741
rect 22557 24732 22569 24735
rect 20772 24704 22569 24732
rect 20772 24692 20778 24704
rect 22557 24701 22569 24704
rect 22603 24701 22615 24735
rect 22830 24732 22836 24744
rect 22791 24704 22836 24732
rect 22557 24695 22615 24701
rect 22830 24692 22836 24704
rect 22888 24692 22894 24744
rect 23014 24692 23020 24744
rect 23072 24732 23078 24744
rect 24121 24735 24179 24741
rect 24121 24732 24133 24735
rect 23072 24704 24133 24732
rect 23072 24692 23078 24704
rect 24121 24701 24133 24704
rect 24167 24732 24179 24735
rect 24486 24732 24492 24744
rect 24167 24704 24492 24732
rect 24167 24701 24179 24704
rect 24121 24695 24179 24701
rect 24486 24692 24492 24704
rect 24544 24692 24550 24744
rect 25148 24741 25176 24772
rect 25406 24760 25412 24772
rect 25464 24760 25470 24812
rect 25593 24803 25651 24809
rect 25593 24769 25605 24803
rect 25639 24800 25651 24803
rect 25682 24800 25688 24812
rect 25639 24772 25688 24800
rect 25639 24769 25651 24772
rect 25593 24763 25651 24769
rect 25682 24760 25688 24772
rect 25740 24760 25746 24812
rect 26237 24803 26295 24809
rect 26237 24769 26249 24803
rect 26283 24769 26295 24803
rect 26237 24763 26295 24769
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24701 25191 24735
rect 25424 24732 25452 24760
rect 25958 24732 25964 24744
rect 25424 24704 25964 24732
rect 25133 24695 25191 24701
rect 25958 24692 25964 24704
rect 26016 24692 26022 24744
rect 26252 24720 26280 24763
rect 26326 24760 26332 24812
rect 26384 24800 26390 24812
rect 27172 24800 27200 24840
rect 27341 24837 27353 24840
rect 27387 24837 27399 24871
rect 27341 24831 27399 24837
rect 27430 24828 27436 24880
rect 27488 24868 27494 24880
rect 29914 24868 29920 24880
rect 27488 24840 29920 24868
rect 27488 24828 27494 24840
rect 29914 24828 29920 24840
rect 29972 24828 29978 24880
rect 30282 24868 30288 24880
rect 30243 24840 30288 24868
rect 30282 24828 30288 24840
rect 30340 24828 30346 24880
rect 29822 24800 29828 24812
rect 26384 24772 26429 24800
rect 26804 24772 27200 24800
rect 28552 24772 29828 24800
rect 26384 24760 26390 24772
rect 26694 24732 26700 24744
rect 26344 24720 26700 24732
rect 26252 24704 26700 24720
rect 26252 24692 26372 24704
rect 26694 24692 26700 24704
rect 26752 24692 26758 24744
rect 23842 24664 23848 24676
rect 19812 24636 21956 24664
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 1854 24596 1860 24608
rect 1627 24568 1860 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 1854 24556 1860 24568
rect 1912 24556 1918 24608
rect 9582 24556 9588 24608
rect 9640 24596 9646 24608
rect 13262 24596 13268 24608
rect 9640 24568 13268 24596
rect 9640 24556 9646 24568
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 13449 24599 13507 24605
rect 13449 24596 13461 24599
rect 13412 24568 13461 24596
rect 13412 24556 13418 24568
rect 13449 24565 13461 24568
rect 13495 24565 13507 24599
rect 14642 24596 14648 24608
rect 14603 24568 14648 24596
rect 13449 24559 13507 24565
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 15286 24596 15292 24608
rect 15247 24568 15292 24596
rect 15286 24556 15292 24568
rect 15344 24556 15350 24608
rect 15930 24556 15936 24608
rect 15988 24596 15994 24608
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 15988 24568 16221 24596
rect 15988 24556 15994 24568
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 21928 24596 21956 24636
rect 22066 24636 23848 24664
rect 22066 24596 22094 24636
rect 23842 24624 23848 24636
rect 23900 24624 23906 24676
rect 24302 24624 24308 24676
rect 24360 24664 24366 24676
rect 26804 24664 26832 24772
rect 27157 24735 27215 24741
rect 27157 24701 27169 24735
rect 27203 24732 27215 24735
rect 27203 24720 27292 24732
rect 27203 24716 27384 24720
rect 27203 24704 27476 24716
rect 27203 24701 27215 24704
rect 27157 24695 27215 24701
rect 27264 24692 27476 24704
rect 27982 24692 27988 24744
rect 28040 24732 28046 24744
rect 28552 24732 28580 24772
rect 29822 24760 29828 24772
rect 29880 24760 29886 24812
rect 32858 24760 32864 24812
rect 32916 24800 32922 24812
rect 32953 24803 33011 24809
rect 32953 24800 32965 24803
rect 32916 24772 32965 24800
rect 32916 24760 32922 24772
rect 32953 24769 32965 24772
rect 32999 24769 33011 24803
rect 32953 24763 33011 24769
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24800 33103 24803
rect 33778 24800 33784 24812
rect 33091 24772 33784 24800
rect 33091 24769 33103 24772
rect 33045 24763 33103 24769
rect 33778 24760 33784 24772
rect 33836 24760 33842 24812
rect 35342 24760 35348 24812
rect 35400 24800 35406 24812
rect 38013 24803 38071 24809
rect 38013 24800 38025 24803
rect 35400 24772 38025 24800
rect 35400 24760 35406 24772
rect 38013 24769 38025 24772
rect 38059 24769 38071 24803
rect 38013 24763 38071 24769
rect 28994 24732 29000 24744
rect 28040 24704 28580 24732
rect 28955 24704 29000 24732
rect 28040 24692 28046 24704
rect 28994 24692 29000 24704
rect 29052 24692 29058 24744
rect 29457 24735 29515 24741
rect 29457 24701 29469 24735
rect 29503 24732 29515 24735
rect 30006 24732 30012 24744
rect 29503 24704 30012 24732
rect 29503 24701 29515 24704
rect 29457 24695 29515 24701
rect 30006 24692 30012 24704
rect 30064 24692 30070 24744
rect 30190 24732 30196 24744
rect 30151 24704 30196 24732
rect 30190 24692 30196 24704
rect 30248 24692 30254 24744
rect 30837 24735 30895 24741
rect 30837 24701 30849 24735
rect 30883 24732 30895 24735
rect 32030 24732 32036 24744
rect 30883 24704 32036 24732
rect 30883 24701 30895 24704
rect 30837 24695 30895 24701
rect 32030 24692 32036 24704
rect 32088 24692 32094 24744
rect 27356 24688 27476 24692
rect 24360 24636 26832 24664
rect 27448 24664 27476 24688
rect 29178 24664 29184 24676
rect 27448 24636 29184 24664
rect 24360 24624 24366 24636
rect 29178 24624 29184 24636
rect 29236 24664 29242 24676
rect 30208 24664 30236 24692
rect 29236 24636 30236 24664
rect 29236 24624 29242 24636
rect 21928 24568 22094 24596
rect 16209 24559 16267 24565
rect 23474 24556 23480 24608
rect 23532 24596 23538 24608
rect 25685 24599 25743 24605
rect 25685 24596 25697 24599
rect 23532 24568 25697 24596
rect 23532 24556 23538 24568
rect 25685 24565 25697 24568
rect 25731 24565 25743 24599
rect 25685 24559 25743 24565
rect 26050 24556 26056 24608
rect 26108 24596 26114 24608
rect 27614 24596 27620 24608
rect 26108 24568 27620 24596
rect 26108 24556 26114 24568
rect 27614 24556 27620 24568
rect 27672 24596 27678 24608
rect 29086 24596 29092 24608
rect 27672 24568 29092 24596
rect 27672 24556 27678 24568
rect 29086 24556 29092 24568
rect 29144 24556 29150 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 10594 24392 10600 24404
rect 9916 24364 10600 24392
rect 9916 24352 9922 24364
rect 10594 24352 10600 24364
rect 10652 24352 10658 24404
rect 11422 24352 11428 24404
rect 11480 24392 11486 24404
rect 11974 24392 11980 24404
rect 11480 24364 11980 24392
rect 11480 24352 11486 24364
rect 11974 24352 11980 24364
rect 12032 24352 12038 24404
rect 13262 24352 13268 24404
rect 13320 24392 13326 24404
rect 15010 24392 15016 24404
rect 13320 24364 15016 24392
rect 13320 24352 13326 24364
rect 15010 24352 15016 24364
rect 15068 24352 15074 24404
rect 20254 24392 20260 24404
rect 15120 24364 20260 24392
rect 12158 24324 12164 24336
rect 10152 24296 12164 24324
rect 9398 24256 9404 24268
rect 9359 24228 9404 24256
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 10152 24265 10180 24296
rect 12158 24284 12164 24296
rect 12216 24324 12222 24336
rect 14550 24324 14556 24336
rect 12216 24296 14556 24324
rect 12216 24284 12222 24296
rect 14550 24284 14556 24296
rect 14608 24284 14614 24336
rect 10137 24259 10195 24265
rect 10137 24225 10149 24259
rect 10183 24225 10195 24259
rect 10137 24219 10195 24225
rect 11149 24259 11207 24265
rect 11149 24225 11161 24259
rect 11195 24256 11207 24259
rect 11238 24256 11244 24268
rect 11195 24228 11244 24256
rect 11195 24225 11207 24228
rect 11149 24219 11207 24225
rect 11238 24216 11244 24228
rect 11296 24256 11302 24268
rect 12342 24256 12348 24268
rect 11296 24228 12348 24256
rect 11296 24216 11302 24228
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 12526 24256 12532 24268
rect 12487 24228 12532 24256
rect 12526 24216 12532 24228
rect 12584 24256 12590 24268
rect 13262 24256 13268 24268
rect 12584 24228 13268 24256
rect 12584 24216 12590 24228
rect 13262 24216 13268 24228
rect 13320 24216 13326 24268
rect 15120 24256 15148 24364
rect 20254 24352 20260 24364
rect 20312 24352 20318 24404
rect 24210 24352 24216 24404
rect 24268 24392 24274 24404
rect 24673 24395 24731 24401
rect 24673 24392 24685 24395
rect 24268 24364 24685 24392
rect 24268 24352 24274 24364
rect 24673 24361 24685 24364
rect 24719 24361 24731 24395
rect 24673 24355 24731 24361
rect 24762 24352 24768 24404
rect 24820 24392 24826 24404
rect 24820 24364 25268 24392
rect 24820 24352 24826 24364
rect 19886 24324 19892 24336
rect 14384 24228 15148 24256
rect 15212 24296 19892 24324
rect 14277 24201 14335 24207
rect 1762 24188 1768 24200
rect 1723 24160 1768 24188
rect 1762 24148 1768 24160
rect 1820 24148 1826 24200
rect 1854 24148 1860 24200
rect 1912 24188 1918 24200
rect 8297 24191 8355 24197
rect 8297 24188 8309 24191
rect 1912 24160 8309 24188
rect 1912 24148 1918 24160
rect 8297 24157 8309 24160
rect 8343 24157 8355 24191
rect 8297 24151 8355 24157
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13722 24188 13728 24200
rect 13587 24160 13728 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 14277 24167 14289 24201
rect 14323 24198 14335 24201
rect 14384 24198 14412 24228
rect 15212 24207 15240 24296
rect 19886 24284 19892 24296
rect 19944 24284 19950 24336
rect 24118 24324 24124 24336
rect 20456 24296 24124 24324
rect 15930 24256 15936 24268
rect 15891 24228 15936 24256
rect 15930 24216 15936 24228
rect 15988 24216 15994 24268
rect 16850 24216 16856 24268
rect 16908 24256 16914 24268
rect 17589 24259 17647 24265
rect 17589 24256 17601 24259
rect 16908 24228 17601 24256
rect 16908 24216 16914 24228
rect 17589 24225 17601 24228
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 17770 24216 17776 24268
rect 17828 24256 17834 24268
rect 17957 24259 18015 24265
rect 17957 24256 17969 24259
rect 17828 24228 17969 24256
rect 17828 24216 17834 24228
rect 17957 24225 17969 24228
rect 18003 24225 18015 24259
rect 17957 24219 18015 24225
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 20456 24256 20484 24296
rect 24118 24284 24124 24296
rect 24176 24324 24182 24336
rect 24854 24324 24860 24336
rect 24176 24296 24860 24324
rect 24176 24284 24182 24296
rect 24854 24284 24860 24296
rect 24912 24284 24918 24336
rect 18288 24228 20484 24256
rect 18288 24216 18294 24228
rect 20530 24216 20536 24268
rect 20588 24256 20594 24268
rect 21085 24259 21143 24265
rect 21085 24256 21097 24259
rect 20588 24228 21097 24256
rect 20588 24216 20594 24228
rect 21085 24225 21097 24228
rect 21131 24225 21143 24259
rect 21085 24219 21143 24225
rect 21266 24216 21272 24268
rect 21324 24256 21330 24268
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 21324 24228 21373 24256
rect 21324 24216 21330 24228
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 21361 24219 21419 24225
rect 25240 24256 25268 24364
rect 25498 24352 25504 24404
rect 25556 24392 25562 24404
rect 25961 24395 26019 24401
rect 25961 24392 25973 24395
rect 25556 24364 25973 24392
rect 25556 24352 25562 24364
rect 25961 24361 25973 24364
rect 26007 24361 26019 24395
rect 26510 24392 26516 24404
rect 26423 24364 26516 24392
rect 25961 24355 26019 24361
rect 26510 24352 26516 24364
rect 26568 24392 26574 24404
rect 37458 24392 37464 24404
rect 26568 24364 37464 24392
rect 26568 24352 26574 24364
rect 37458 24352 37464 24364
rect 37516 24352 37522 24404
rect 25682 24284 25688 24336
rect 25740 24324 25746 24336
rect 26418 24324 26424 24336
rect 25740 24296 26424 24324
rect 25740 24284 25746 24296
rect 26418 24284 26424 24296
rect 26476 24284 26482 24336
rect 25498 24256 25504 24268
rect 25240 24228 25504 24256
rect 14323 24170 14412 24198
rect 15197 24201 15255 24207
rect 14323 24167 14335 24170
rect 14277 24161 14335 24167
rect 15197 24167 15209 24201
rect 15243 24167 15255 24201
rect 15197 24161 15255 24167
rect 19702 24148 19708 24200
rect 19760 24188 19766 24200
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 19760 24160 19809 24188
rect 19760 24148 19766 24160
rect 19797 24157 19809 24160
rect 19843 24188 19855 24191
rect 20438 24188 20444 24200
rect 19843 24160 20444 24188
rect 19843 24157 19855 24160
rect 19797 24151 19855 24157
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 25240 24197 25268 24228
rect 25498 24216 25504 24228
rect 25556 24216 25562 24268
rect 24581 24191 24639 24197
rect 24581 24188 24593 24191
rect 23860 24160 24593 24188
rect 23860 24132 23888 24160
rect 24581 24157 24593 24160
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 25225 24191 25283 24197
rect 25225 24157 25237 24191
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 25314 24148 25320 24200
rect 25372 24188 25378 24200
rect 25869 24191 25927 24197
rect 25869 24188 25881 24191
rect 25372 24160 25881 24188
rect 25372 24148 25378 24160
rect 25869 24157 25881 24160
rect 25915 24188 25927 24191
rect 26418 24188 26424 24200
rect 25915 24160 26424 24188
rect 25915 24157 25927 24160
rect 25869 24151 25927 24157
rect 26418 24148 26424 24160
rect 26476 24148 26482 24200
rect 26528 24197 26556 24352
rect 26602 24284 26608 24336
rect 26660 24324 26666 24336
rect 26660 24296 26705 24324
rect 26660 24284 26666 24296
rect 27982 24284 27988 24336
rect 28040 24324 28046 24336
rect 30558 24324 30564 24336
rect 28040 24296 30564 24324
rect 28040 24284 28046 24296
rect 30558 24284 30564 24296
rect 30616 24284 30622 24336
rect 31754 24284 31760 24336
rect 31812 24324 31818 24336
rect 31812 24296 32444 24324
rect 31812 24284 31818 24296
rect 28442 24256 28448 24268
rect 28403 24228 28448 24256
rect 28442 24216 28448 24228
rect 28500 24216 28506 24268
rect 30006 24256 30012 24268
rect 29967 24228 30012 24256
rect 30006 24216 30012 24228
rect 30064 24216 30070 24268
rect 31018 24256 31024 24268
rect 30979 24228 31024 24256
rect 31018 24216 31024 24228
rect 31076 24256 31082 24268
rect 31294 24256 31300 24268
rect 31076 24228 31300 24256
rect 31076 24216 31082 24228
rect 31294 24216 31300 24228
rect 31352 24216 31358 24268
rect 32125 24259 32183 24265
rect 32125 24225 32137 24259
rect 32171 24256 32183 24259
rect 32306 24256 32312 24268
rect 32171 24228 32312 24256
rect 32171 24225 32183 24228
rect 32125 24219 32183 24225
rect 32306 24216 32312 24228
rect 32364 24216 32370 24268
rect 32416 24265 32444 24296
rect 32401 24259 32459 24265
rect 32401 24225 32413 24259
rect 32447 24225 32459 24259
rect 32401 24219 32459 24225
rect 34606 24216 34612 24268
rect 34664 24256 34670 24268
rect 37734 24256 37740 24268
rect 34664 24228 37740 24256
rect 34664 24216 34670 24228
rect 37734 24216 37740 24228
rect 37792 24216 37798 24268
rect 26513 24191 26571 24197
rect 26513 24157 26525 24191
rect 26559 24157 26571 24191
rect 26513 24151 26571 24157
rect 27433 24191 27491 24197
rect 27433 24157 27445 24191
rect 27479 24157 27491 24191
rect 38286 24188 38292 24200
rect 27433 24151 27491 24157
rect 30944 24160 31984 24188
rect 38247 24160 38292 24188
rect 10229 24123 10287 24129
rect 10229 24089 10241 24123
rect 10275 24120 10287 24123
rect 11054 24120 11060 24132
rect 10275 24092 11060 24120
rect 10275 24089 10287 24092
rect 10229 24083 10287 24089
rect 11054 24080 11060 24092
rect 11112 24080 11118 24132
rect 11238 24080 11244 24132
rect 11296 24120 11302 24132
rect 11977 24123 12035 24129
rect 11977 24120 11989 24123
rect 11296 24092 11989 24120
rect 11296 24080 11302 24092
rect 11977 24089 11989 24092
rect 12023 24089 12035 24123
rect 11977 24083 12035 24089
rect 12066 24080 12072 24132
rect 12124 24120 12130 24132
rect 13633 24123 13691 24129
rect 12124 24092 12169 24120
rect 12124 24080 12130 24092
rect 13633 24089 13645 24123
rect 13679 24120 13691 24123
rect 15102 24120 15108 24132
rect 13679 24092 15108 24120
rect 13679 24089 13691 24092
rect 13633 24083 13691 24089
rect 15102 24080 15108 24092
rect 15160 24120 15166 24132
rect 15160 24092 15976 24120
rect 15160 24080 15166 24092
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 5534 24052 5540 24064
rect 1627 24024 5540 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 5534 24012 5540 24024
rect 5592 24012 5598 24064
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 10594 24052 10600 24064
rect 8435 24024 10600 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 13814 24012 13820 24064
rect 13872 24052 13878 24064
rect 14369 24055 14427 24061
rect 14369 24052 14381 24055
rect 13872 24024 14381 24052
rect 13872 24012 13878 24024
rect 14369 24021 14381 24024
rect 14415 24021 14427 24055
rect 14369 24015 14427 24021
rect 15289 24055 15347 24061
rect 15289 24021 15301 24055
rect 15335 24052 15347 24055
rect 15838 24052 15844 24064
rect 15335 24024 15844 24052
rect 15335 24021 15347 24024
rect 15289 24015 15347 24021
rect 15838 24012 15844 24024
rect 15896 24012 15902 24064
rect 15948 24052 15976 24092
rect 16022 24080 16028 24132
rect 16080 24120 16086 24132
rect 16945 24123 17003 24129
rect 16080 24092 16125 24120
rect 16080 24080 16086 24092
rect 16945 24089 16957 24123
rect 16991 24120 17003 24123
rect 17034 24120 17040 24132
rect 16991 24092 17040 24120
rect 16991 24089 17003 24092
rect 16945 24083 17003 24089
rect 17034 24080 17040 24092
rect 17092 24080 17098 24132
rect 17681 24123 17739 24129
rect 17681 24089 17693 24123
rect 17727 24120 17739 24123
rect 18230 24120 18236 24132
rect 17727 24092 18236 24120
rect 17727 24089 17739 24092
rect 17681 24083 17739 24089
rect 18230 24080 18236 24092
rect 18288 24080 18294 24132
rect 18414 24080 18420 24132
rect 18472 24120 18478 24132
rect 19610 24120 19616 24132
rect 18472 24092 19616 24120
rect 18472 24080 18478 24092
rect 19610 24080 19616 24092
rect 19668 24080 19674 24132
rect 20714 24120 20720 24132
rect 20548 24092 20720 24120
rect 18506 24052 18512 24064
rect 15948 24024 18512 24052
rect 18506 24012 18512 24024
rect 18564 24052 18570 24064
rect 18874 24052 18880 24064
rect 18564 24024 18880 24052
rect 18564 24012 18570 24024
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24052 19947 24055
rect 20548 24052 20576 24092
rect 20714 24080 20720 24092
rect 20772 24080 20778 24132
rect 21174 24080 21180 24132
rect 21232 24120 21238 24132
rect 23014 24120 23020 24132
rect 21232 24092 21277 24120
rect 22975 24092 23020 24120
rect 21232 24080 21238 24092
rect 23014 24080 23020 24092
rect 23072 24080 23078 24132
rect 23109 24123 23167 24129
rect 23109 24089 23121 24123
rect 23155 24089 23167 24123
rect 23109 24083 23167 24089
rect 19935 24024 20576 24052
rect 23124 24052 23152 24083
rect 23842 24080 23848 24132
rect 23900 24080 23906 24132
rect 24029 24123 24087 24129
rect 24029 24089 24041 24123
rect 24075 24120 24087 24123
rect 24118 24120 24124 24132
rect 24075 24092 24124 24120
rect 24075 24089 24087 24092
rect 24029 24083 24087 24089
rect 24118 24080 24124 24092
rect 24176 24080 24182 24132
rect 27448 24064 27476 24151
rect 27982 24080 27988 24132
rect 28040 24120 28046 24132
rect 28158 24123 28216 24129
rect 28158 24120 28170 24123
rect 28040 24092 28170 24120
rect 28040 24080 28046 24092
rect 28158 24089 28170 24092
rect 28204 24089 28216 24123
rect 28158 24083 28216 24089
rect 28254 24123 28312 24129
rect 28254 24089 28266 24123
rect 28300 24089 28312 24123
rect 28254 24083 28312 24089
rect 30101 24123 30159 24129
rect 30101 24089 30113 24123
rect 30147 24120 30159 24123
rect 30944 24120 30972 24160
rect 30147 24092 30972 24120
rect 30147 24089 30159 24092
rect 30101 24083 30159 24089
rect 25317 24055 25375 24061
rect 25317 24052 25329 24055
rect 23124 24024 25329 24052
rect 19935 24021 19947 24024
rect 19889 24015 19947 24021
rect 25317 24021 25329 24024
rect 25363 24021 25375 24055
rect 25317 24015 25375 24021
rect 25406 24012 25412 24064
rect 25464 24052 25470 24064
rect 27430 24052 27436 24064
rect 25464 24024 27436 24052
rect 25464 24012 25470 24024
rect 27430 24012 27436 24024
rect 27488 24012 27494 24064
rect 27525 24055 27583 24061
rect 27525 24021 27537 24055
rect 27571 24052 27583 24055
rect 28276 24052 28304 24083
rect 27571 24024 28304 24052
rect 31956 24052 31984 24160
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 32214 24080 32220 24132
rect 32272 24120 32278 24132
rect 32272 24092 32317 24120
rect 32272 24080 32278 24092
rect 34054 24052 34060 24064
rect 31956 24024 34060 24052
rect 27571 24021 27583 24024
rect 27525 24015 27583 24021
rect 34054 24012 34060 24024
rect 34112 24012 34118 24064
rect 38102 24052 38108 24064
rect 38063 24024 38108 24052
rect 38102 24012 38108 24024
rect 38160 24012 38166 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1670 23808 1676 23860
rect 1728 23848 1734 23860
rect 1765 23851 1823 23857
rect 1765 23848 1777 23851
rect 1728 23820 1777 23848
rect 1728 23808 1734 23820
rect 1765 23817 1777 23820
rect 1811 23817 1823 23851
rect 2406 23848 2412 23860
rect 2367 23820 2412 23848
rect 1765 23811 1823 23817
rect 2406 23808 2412 23820
rect 2464 23808 2470 23860
rect 10318 23848 10324 23860
rect 10279 23820 10324 23848
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 14458 23848 14464 23860
rect 10980 23820 14464 23848
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23681 2007 23715
rect 2590 23712 2596 23724
rect 2551 23684 2596 23712
rect 1949 23675 2007 23681
rect 1964 23644 1992 23675
rect 2590 23672 2596 23684
rect 2648 23672 2654 23724
rect 10502 23712 10508 23724
rect 10463 23684 10508 23712
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10980 23721 11008 23820
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 18230 23848 18236 23860
rect 14568 23820 18092 23848
rect 18191 23820 18236 23848
rect 11054 23740 11060 23792
rect 11112 23780 11118 23792
rect 13814 23780 13820 23792
rect 11112 23752 11157 23780
rect 11256 23752 12664 23780
rect 13775 23752 13820 23780
rect 11112 23740 11118 23752
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 6454 23644 6460 23656
rect 1964 23616 6460 23644
rect 6454 23604 6460 23616
rect 6512 23604 6518 23656
rect 9950 23604 9956 23656
rect 10008 23644 10014 23656
rect 11256 23644 11284 23752
rect 11606 23672 11612 23724
rect 11664 23712 11670 23724
rect 11793 23715 11851 23721
rect 11793 23712 11805 23715
rect 11664 23684 11805 23712
rect 11664 23672 11670 23684
rect 11793 23681 11805 23684
rect 11839 23681 11851 23715
rect 11793 23675 11851 23681
rect 12529 23715 12587 23721
rect 12529 23681 12541 23715
rect 12575 23681 12587 23715
rect 12529 23675 12587 23681
rect 10008 23616 11284 23644
rect 10008 23604 10014 23616
rect 10778 23536 10784 23588
rect 10836 23576 10842 23588
rect 12544 23576 12572 23675
rect 12636 23644 12664 23752
rect 13814 23740 13820 23752
rect 13872 23740 13878 23792
rect 14568 23653 14596 23820
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 15381 23783 15439 23789
rect 15381 23780 15393 23783
rect 14700 23752 15393 23780
rect 14700 23740 14706 23752
rect 15381 23749 15393 23752
rect 15427 23749 15439 23783
rect 15381 23743 15439 23749
rect 16301 23783 16359 23789
rect 16301 23749 16313 23783
rect 16347 23780 16359 23783
rect 17770 23780 17776 23792
rect 16347 23752 17776 23780
rect 16347 23749 16359 23752
rect 16301 23743 16359 23749
rect 17770 23740 17776 23752
rect 17828 23740 17834 23792
rect 18064 23780 18092 23820
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 19886 23848 19892 23860
rect 18432 23820 19892 23848
rect 18432 23780 18460 23820
rect 19886 23808 19892 23820
rect 19944 23808 19950 23860
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 28442 23848 28448 23860
rect 23348 23820 28448 23848
rect 23348 23808 23354 23820
rect 28442 23808 28448 23820
rect 28500 23808 28506 23860
rect 30282 23808 30288 23860
rect 30340 23848 30346 23860
rect 30377 23851 30435 23857
rect 30377 23848 30389 23851
rect 30340 23820 30389 23848
rect 30340 23808 30346 23820
rect 30377 23817 30389 23820
rect 30423 23817 30435 23851
rect 30377 23811 30435 23817
rect 31665 23851 31723 23857
rect 31665 23817 31677 23851
rect 31711 23848 31723 23851
rect 32214 23848 32220 23860
rect 31711 23820 32220 23848
rect 31711 23817 31723 23820
rect 31665 23811 31723 23817
rect 32214 23808 32220 23820
rect 32272 23808 32278 23860
rect 33689 23851 33747 23857
rect 33689 23817 33701 23851
rect 33735 23848 33747 23851
rect 34790 23848 34796 23860
rect 33735 23820 34796 23848
rect 33735 23817 33747 23820
rect 33689 23811 33747 23817
rect 34790 23808 34796 23820
rect 34848 23808 34854 23860
rect 37829 23851 37887 23857
rect 37829 23817 37841 23851
rect 37875 23848 37887 23851
rect 38010 23848 38016 23860
rect 37875 23820 38016 23848
rect 37875 23817 37887 23820
rect 37829 23811 37887 23817
rect 38010 23808 38016 23820
rect 38068 23808 38074 23860
rect 18874 23780 18880 23792
rect 18064 23752 18460 23780
rect 18835 23752 18880 23780
rect 18874 23740 18880 23752
rect 18932 23740 18938 23792
rect 18969 23783 19027 23789
rect 18969 23749 18981 23783
rect 19015 23780 19027 23783
rect 19518 23780 19524 23792
rect 19015 23752 19524 23780
rect 19015 23749 19027 23752
rect 18969 23743 19027 23749
rect 19518 23740 19524 23752
rect 19576 23740 19582 23792
rect 20342 23783 20400 23789
rect 20342 23749 20354 23783
rect 20388 23780 20400 23783
rect 20714 23780 20720 23792
rect 20388 23752 20720 23780
rect 20388 23749 20400 23752
rect 20342 23743 20400 23749
rect 20714 23740 20720 23752
rect 20772 23740 20778 23792
rect 21910 23740 21916 23792
rect 21968 23780 21974 23792
rect 22086 23783 22144 23789
rect 22086 23780 22098 23783
rect 21968 23752 22098 23780
rect 21968 23740 21974 23752
rect 22086 23749 22098 23752
rect 22132 23749 22144 23783
rect 22086 23743 22144 23749
rect 22198 23783 22256 23789
rect 22198 23749 22210 23783
rect 22244 23780 22256 23783
rect 22370 23780 22376 23792
rect 22244 23752 22376 23780
rect 22244 23749 22256 23752
rect 22198 23743 22256 23749
rect 22370 23740 22376 23752
rect 22428 23740 22434 23792
rect 24302 23780 24308 23792
rect 24263 23752 24308 23780
rect 24302 23740 24308 23752
rect 24360 23740 24366 23792
rect 26513 23783 26571 23789
rect 26513 23749 26525 23783
rect 26559 23780 26571 23783
rect 27341 23783 27399 23789
rect 27341 23780 27353 23783
rect 26559 23752 27353 23780
rect 26559 23749 26571 23752
rect 26513 23743 26571 23749
rect 27341 23749 27353 23752
rect 27387 23749 27399 23783
rect 28902 23780 28908 23792
rect 28863 23752 28908 23780
rect 27341 23743 27399 23749
rect 28902 23740 28908 23752
rect 28960 23740 28966 23792
rect 30558 23740 30564 23792
rect 30616 23780 30622 23792
rect 31478 23780 31484 23792
rect 30616 23752 31484 23780
rect 30616 23740 30622 23752
rect 31478 23740 31484 23752
rect 31536 23780 31542 23792
rect 32585 23783 32643 23789
rect 32585 23780 32597 23783
rect 31536 23752 32597 23780
rect 31536 23740 31542 23752
rect 32585 23749 32597 23752
rect 32631 23749 32643 23783
rect 32585 23743 32643 23749
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16592 23684 16865 23712
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 12636 23616 13737 23644
rect 13725 23613 13737 23616
rect 13771 23613 13783 23647
rect 13725 23607 13783 23613
rect 14553 23647 14611 23653
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 15289 23647 15347 23653
rect 15289 23613 15301 23647
rect 15335 23644 15347 23647
rect 15930 23644 15936 23656
rect 15335 23616 15936 23644
rect 15335 23613 15347 23616
rect 15289 23607 15347 23613
rect 15930 23604 15936 23616
rect 15988 23604 15994 23656
rect 10836 23548 12572 23576
rect 12713 23579 12771 23585
rect 10836 23536 10842 23548
rect 12713 23545 12725 23579
rect 12759 23576 12771 23579
rect 16482 23576 16488 23588
rect 12759 23548 16488 23576
rect 12759 23545 12771 23548
rect 12713 23539 12771 23545
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12066 23508 12072 23520
rect 11931 23480 12072 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12066 23468 12072 23480
rect 12124 23508 12130 23520
rect 12894 23508 12900 23520
rect 12124 23480 12900 23508
rect 12124 23468 12130 23480
rect 12894 23468 12900 23480
rect 12952 23468 12958 23520
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 16592 23508 16620 23684
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17034 23672 17040 23724
rect 17092 23712 17098 23724
rect 17402 23712 17408 23724
rect 17092 23684 17408 23712
rect 17092 23672 17098 23684
rect 17402 23672 17408 23684
rect 17460 23712 17466 23724
rect 17497 23715 17555 23721
rect 17497 23712 17509 23715
rect 17460 23684 17509 23712
rect 17460 23672 17466 23684
rect 17497 23681 17509 23684
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23712 18199 23715
rect 18414 23712 18420 23724
rect 18187 23684 18420 23712
rect 18187 23681 18199 23684
rect 18141 23675 18199 23681
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 23569 23715 23627 23721
rect 23569 23712 23581 23715
rect 23216 23684 23581 23712
rect 23216 23656 23244 23684
rect 23569 23681 23581 23684
rect 23615 23681 23627 23715
rect 24210 23712 24216 23724
rect 24171 23684 24216 23712
rect 23569 23675 23627 23681
rect 24210 23672 24216 23684
rect 24268 23672 24274 23724
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 20257 23647 20315 23653
rect 20257 23613 20269 23647
rect 20303 23644 20315 23647
rect 20530 23644 20536 23656
rect 20303 23616 20536 23644
rect 20303 23613 20315 23616
rect 20257 23607 20315 23613
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 20714 23644 20720 23656
rect 20675 23616 20720 23644
rect 20714 23604 20720 23616
rect 20772 23604 20778 23656
rect 21726 23604 21732 23656
rect 21784 23644 21790 23656
rect 22373 23647 22431 23653
rect 22373 23644 22385 23647
rect 21784 23616 22385 23644
rect 21784 23604 21790 23616
rect 22373 23613 22385 23616
rect 22419 23613 22431 23647
rect 22373 23607 22431 23613
rect 23198 23604 23204 23656
rect 23256 23604 23262 23656
rect 24872 23644 24900 23675
rect 25222 23672 25228 23724
rect 25280 23712 25286 23724
rect 25501 23715 25559 23721
rect 25501 23712 25513 23715
rect 25280 23684 25513 23712
rect 25280 23672 25286 23684
rect 25501 23681 25513 23684
rect 25547 23712 25559 23715
rect 25682 23712 25688 23724
rect 25547 23684 25688 23712
rect 25547 23681 25559 23684
rect 25501 23675 25559 23681
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23681 26479 23715
rect 26421 23675 26479 23681
rect 24946 23644 24952 23656
rect 24872 23616 24952 23644
rect 24946 23604 24952 23616
rect 25004 23644 25010 23656
rect 25590 23644 25596 23656
rect 25004 23616 25596 23644
rect 25004 23604 25010 23616
rect 25590 23604 25596 23616
rect 25648 23604 25654 23656
rect 19429 23579 19487 23585
rect 19429 23545 19441 23579
rect 19475 23576 19487 23579
rect 22002 23576 22008 23588
rect 19475 23548 22008 23576
rect 19475 23545 19487 23548
rect 19429 23539 19487 23545
rect 22002 23536 22008 23548
rect 22060 23536 22066 23588
rect 26436 23576 26464 23675
rect 29822 23672 29828 23724
rect 29880 23712 29886 23724
rect 30282 23712 30288 23724
rect 29880 23684 30288 23712
rect 29880 23672 29886 23684
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 30929 23715 30987 23721
rect 30929 23681 30941 23715
rect 30975 23681 30987 23715
rect 30929 23675 30987 23681
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23712 31631 23715
rect 31846 23712 31852 23724
rect 31619 23684 31852 23712
rect 31619 23681 31631 23684
rect 31573 23675 31631 23681
rect 26878 23604 26884 23656
rect 26936 23644 26942 23656
rect 27249 23647 27307 23653
rect 27249 23644 27261 23647
rect 26936 23616 27261 23644
rect 26936 23604 26942 23616
rect 27249 23613 27261 23616
rect 27295 23613 27307 23647
rect 27522 23644 27528 23656
rect 27483 23616 27528 23644
rect 27249 23607 27307 23613
rect 27522 23604 27528 23616
rect 27580 23644 27586 23656
rect 28166 23644 28172 23656
rect 27580 23616 28172 23644
rect 27580 23604 27586 23616
rect 28166 23604 28172 23616
rect 28224 23604 28230 23656
rect 28810 23644 28816 23656
rect 28771 23616 28816 23644
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 29086 23644 29092 23656
rect 29047 23616 29092 23644
rect 29086 23604 29092 23616
rect 29144 23604 29150 23656
rect 30742 23576 30748 23588
rect 26436 23548 30748 23576
rect 30742 23536 30748 23548
rect 30800 23536 30806 23588
rect 30944 23576 30972 23675
rect 31846 23672 31852 23684
rect 31904 23672 31910 23724
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23681 32551 23715
rect 33870 23712 33876 23724
rect 33831 23684 33876 23712
rect 32493 23675 32551 23681
rect 32508 23644 32536 23675
rect 33870 23672 33876 23684
rect 33928 23672 33934 23724
rect 37918 23672 37924 23724
rect 37976 23712 37982 23724
rect 38013 23715 38071 23721
rect 38013 23712 38025 23715
rect 37976 23684 38025 23712
rect 37976 23672 37982 23684
rect 38013 23681 38025 23684
rect 38059 23681 38071 23715
rect 38013 23675 38071 23681
rect 34514 23644 34520 23656
rect 32508 23616 34520 23644
rect 34514 23604 34520 23616
rect 34572 23604 34578 23656
rect 32858 23576 32864 23588
rect 30944 23548 32864 23576
rect 32858 23536 32864 23548
rect 32916 23536 32922 23588
rect 13044 23480 16620 23508
rect 13044 23468 13050 23480
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 16945 23511 17003 23517
rect 16945 23508 16957 23511
rect 16908 23480 16957 23508
rect 16908 23468 16914 23480
rect 16945 23477 16957 23480
rect 16991 23477 17003 23511
rect 16945 23471 17003 23477
rect 17494 23468 17500 23520
rect 17552 23508 17558 23520
rect 17589 23511 17647 23517
rect 17589 23508 17601 23511
rect 17552 23480 17601 23508
rect 17552 23468 17558 23480
rect 17589 23477 17601 23480
rect 17635 23477 17647 23511
rect 23658 23508 23664 23520
rect 23619 23480 23664 23508
rect 17589 23471 17647 23477
rect 23658 23468 23664 23480
rect 23716 23468 23722 23520
rect 24946 23508 24952 23520
rect 24907 23480 24952 23508
rect 24946 23468 24952 23480
rect 25004 23468 25010 23520
rect 25222 23468 25228 23520
rect 25280 23508 25286 23520
rect 25593 23511 25651 23517
rect 25593 23508 25605 23511
rect 25280 23480 25605 23508
rect 25280 23468 25286 23480
rect 25593 23477 25605 23480
rect 25639 23477 25651 23511
rect 25593 23471 25651 23477
rect 27430 23468 27436 23520
rect 27488 23508 27494 23520
rect 30466 23508 30472 23520
rect 27488 23480 30472 23508
rect 27488 23468 27494 23480
rect 30466 23468 30472 23480
rect 30524 23468 30530 23520
rect 31018 23508 31024 23520
rect 30979 23480 31024 23508
rect 31018 23468 31024 23480
rect 31076 23468 31082 23520
rect 31846 23468 31852 23520
rect 31904 23508 31910 23520
rect 32674 23508 32680 23520
rect 31904 23480 32680 23508
rect 31904 23468 31910 23480
rect 32674 23468 32680 23480
rect 32732 23468 32738 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 4062 23264 4068 23316
rect 4120 23304 4126 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 4120 23276 9137 23304
rect 4120 23264 4126 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 10689 23307 10747 23313
rect 10689 23304 10701 23307
rect 10192 23276 10701 23304
rect 10192 23264 10198 23276
rect 10689 23273 10701 23276
rect 10735 23304 10747 23307
rect 11238 23304 11244 23316
rect 10735 23276 11244 23304
rect 10735 23273 10747 23276
rect 10689 23267 10747 23273
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 13633 23307 13691 23313
rect 13633 23273 13645 23307
rect 13679 23304 13691 23307
rect 13906 23304 13912 23316
rect 13679 23276 13912 23304
rect 13679 23273 13691 23276
rect 13633 23267 13691 23273
rect 13906 23264 13912 23276
rect 13964 23264 13970 23316
rect 15194 23264 15200 23316
rect 15252 23304 15258 23316
rect 15654 23304 15660 23316
rect 15252 23276 15660 23304
rect 15252 23264 15258 23276
rect 15654 23264 15660 23276
rect 15712 23304 15718 23316
rect 22462 23304 22468 23316
rect 15712 23276 22468 23304
rect 15712 23264 15718 23276
rect 22462 23264 22468 23276
rect 22520 23304 22526 23316
rect 23290 23304 23296 23316
rect 22520 23276 23296 23304
rect 22520 23264 22526 23276
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23934 23304 23940 23316
rect 23895 23276 23940 23304
rect 23934 23264 23940 23276
rect 23992 23264 23998 23316
rect 25498 23264 25504 23316
rect 25556 23304 25562 23316
rect 27798 23304 27804 23316
rect 25556 23276 27660 23304
rect 27759 23276 27804 23304
rect 25556 23264 25562 23276
rect 10778 23196 10784 23248
rect 10836 23236 10842 23248
rect 14090 23236 14096 23248
rect 10836 23208 14096 23236
rect 10836 23196 10842 23208
rect 14090 23196 14096 23208
rect 14148 23196 14154 23248
rect 24026 23236 24032 23248
rect 14384 23208 24032 23236
rect 14384 23177 14412 23208
rect 24026 23196 24032 23208
rect 24084 23196 24090 23248
rect 25774 23236 25780 23248
rect 24688 23208 25780 23236
rect 7285 23171 7343 23177
rect 7285 23137 7297 23171
rect 7331 23168 7343 23171
rect 14369 23171 14427 23177
rect 14369 23168 14381 23171
rect 7331 23140 14381 23168
rect 7331 23137 7343 23140
rect 7285 23131 7343 23137
rect 14369 23137 14381 23140
rect 14415 23137 14427 23171
rect 14642 23168 14648 23180
rect 14603 23140 14648 23168
rect 14369 23131 14427 23137
rect 14642 23128 14648 23140
rect 14700 23128 14706 23180
rect 15841 23171 15899 23177
rect 15841 23137 15853 23171
rect 15887 23168 15899 23171
rect 15930 23168 15936 23180
rect 15887 23140 15936 23168
rect 15887 23137 15899 23140
rect 15841 23131 15899 23137
rect 15930 23128 15936 23140
rect 15988 23128 15994 23180
rect 17126 23128 17132 23180
rect 17184 23168 17190 23180
rect 18417 23171 18475 23177
rect 18417 23168 18429 23171
rect 17184 23140 18429 23168
rect 17184 23128 17190 23140
rect 18417 23137 18429 23140
rect 18463 23168 18475 23171
rect 22922 23168 22928 23180
rect 18463 23140 22928 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 22922 23128 22928 23140
rect 22980 23128 22986 23180
rect 24688 23177 24716 23208
rect 25774 23196 25780 23208
rect 25832 23196 25838 23248
rect 27632 23236 27660 23276
rect 27798 23264 27804 23276
rect 27856 23264 27862 23316
rect 28445 23307 28503 23313
rect 28445 23273 28457 23307
rect 28491 23304 28503 23307
rect 28902 23304 28908 23316
rect 28491 23276 28908 23304
rect 28491 23273 28503 23276
rect 28445 23267 28503 23273
rect 28902 23264 28908 23276
rect 28960 23264 28966 23316
rect 31570 23304 31576 23316
rect 29012 23276 31576 23304
rect 29012 23236 29040 23276
rect 31570 23264 31576 23276
rect 31628 23264 31634 23316
rect 31662 23264 31668 23316
rect 31720 23304 31726 23316
rect 33042 23304 33048 23316
rect 31720 23276 33048 23304
rect 31720 23264 31726 23276
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 33226 23236 33232 23248
rect 27632 23208 29040 23236
rect 29104 23208 33232 23236
rect 24673 23171 24731 23177
rect 24673 23137 24685 23171
rect 24719 23137 24731 23171
rect 24673 23131 24731 23137
rect 26234 23128 26240 23180
rect 26292 23168 26298 23180
rect 29104 23168 29132 23208
rect 33226 23196 33232 23208
rect 33284 23196 33290 23248
rect 26292 23140 29132 23168
rect 29825 23171 29883 23177
rect 26292 23128 26298 23140
rect 5534 23060 5540 23112
rect 5592 23100 5598 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 5592 23072 7205 23100
rect 5592 23060 5598 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7834 23100 7840 23112
rect 7795 23072 7840 23100
rect 7193 23063 7251 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 8904 23072 9321 23100
rect 8904 23060 8910 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 10597 23103 10655 23109
rect 10597 23100 10609 23103
rect 9309 23063 9367 23069
rect 9646 23072 10609 23100
rect 934 22992 940 23044
rect 992 23032 998 23044
rect 9646 23032 9674 23072
rect 10597 23069 10609 23072
rect 10643 23100 10655 23103
rect 10778 23100 10784 23112
rect 10643 23072 10784 23100
rect 10643 23069 10655 23072
rect 10597 23063 10655 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11241 23103 11299 23109
rect 11241 23069 11253 23103
rect 11287 23100 11299 23103
rect 11790 23100 11796 23112
rect 11287 23072 11796 23100
rect 11287 23069 11299 23072
rect 11241 23063 11299 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23100 13599 23103
rect 14090 23100 14096 23112
rect 13587 23072 14096 23100
rect 13587 23069 13599 23072
rect 13541 23063 13599 23069
rect 14090 23060 14096 23072
rect 14148 23060 14154 23112
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23100 19487 23103
rect 20254 23100 20260 23112
rect 19475 23072 20260 23100
rect 19475 23069 19487 23072
rect 19429 23063 19487 23069
rect 20254 23060 20260 23072
rect 20312 23100 20318 23112
rect 20438 23100 20444 23112
rect 20312 23072 20444 23100
rect 20312 23060 20318 23072
rect 20438 23060 20444 23072
rect 20496 23060 20502 23112
rect 20990 23100 20996 23112
rect 20951 23072 20996 23100
rect 20990 23060 20996 23072
rect 21048 23060 21054 23112
rect 21634 23100 21640 23112
rect 21595 23072 21640 23100
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 23658 23100 23664 23112
rect 21775 23072 22094 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 992 23004 9674 23032
rect 992 22992 998 23004
rect 11698 22992 11704 23044
rect 11756 23032 11762 23044
rect 11977 23035 12035 23041
rect 11977 23032 11989 23035
rect 11756 23004 11989 23032
rect 11756 22992 11762 23004
rect 11977 23001 11989 23004
rect 12023 23001 12035 23035
rect 11977 22995 12035 23001
rect 12069 23035 12127 23041
rect 12069 23001 12081 23035
rect 12115 23001 12127 23035
rect 12069 22995 12127 23001
rect 12989 23035 13047 23041
rect 12989 23001 13001 23035
rect 13035 23001 13047 23035
rect 12989 22995 13047 23001
rect 7742 22924 7748 22976
rect 7800 22964 7806 22976
rect 7929 22967 7987 22973
rect 7929 22964 7941 22967
rect 7800 22936 7941 22964
rect 7800 22924 7806 22936
rect 7929 22933 7941 22936
rect 7975 22933 7987 22967
rect 7929 22927 7987 22933
rect 11333 22967 11391 22973
rect 11333 22933 11345 22967
rect 11379 22964 11391 22967
rect 12084 22964 12112 22995
rect 11379 22936 12112 22964
rect 13004 22964 13032 22995
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 14516 23004 14561 23032
rect 14516 22992 14522 23004
rect 15930 22992 15936 23044
rect 15988 23032 15994 23044
rect 16853 23035 16911 23041
rect 15988 23004 16033 23032
rect 15988 22992 15994 23004
rect 16853 23001 16865 23035
rect 16899 23001 16911 23035
rect 17402 23032 17408 23044
rect 17363 23004 17408 23032
rect 16853 22995 16911 23001
rect 16574 22964 16580 22976
rect 13004 22936 16580 22964
rect 11379 22933 11391 22936
rect 11333 22927 11391 22933
rect 16574 22924 16580 22936
rect 16632 22964 16638 22976
rect 16868 22964 16896 22995
rect 17402 22992 17408 23004
rect 17460 22992 17466 23044
rect 17494 22992 17500 23044
rect 17552 23032 17558 23044
rect 19518 23032 19524 23044
rect 17552 23004 17597 23032
rect 19479 23004 19524 23032
rect 17552 22992 17558 23004
rect 19518 22992 19524 23004
rect 19576 22992 19582 23044
rect 22066 23032 22094 23072
rect 23216 23072 23664 23100
rect 22370 23032 22376 23044
rect 22066 23004 22376 23032
rect 22370 22992 22376 23004
rect 22428 22992 22434 23044
rect 22465 23035 22523 23041
rect 22465 23001 22477 23035
rect 22511 23032 22523 23035
rect 23216 23032 23244 23072
rect 23658 23060 23664 23072
rect 23716 23060 23722 23112
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23100 23903 23103
rect 24486 23100 24492 23112
rect 23891 23072 24492 23100
rect 23891 23069 23903 23072
rect 23845 23063 23903 23069
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 26142 23100 26148 23112
rect 26103 23072 26148 23100
rect 26142 23060 26148 23072
rect 26200 23060 26206 23112
rect 27062 23100 27068 23112
rect 27023 23072 27068 23100
rect 27062 23060 27068 23072
rect 27120 23060 27126 23112
rect 27706 23100 27712 23112
rect 27667 23072 27712 23100
rect 27706 23060 27712 23072
rect 27764 23060 27770 23112
rect 28350 23100 28356 23112
rect 28311 23072 28356 23100
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 29012 23109 29040 23140
rect 29825 23137 29837 23171
rect 29871 23168 29883 23171
rect 33778 23168 33784 23180
rect 29871 23140 33784 23168
rect 29871 23137 29883 23140
rect 29825 23131 29883 23137
rect 33778 23128 33784 23140
rect 33836 23128 33842 23180
rect 28997 23103 29055 23109
rect 28997 23069 29009 23103
rect 29043 23069 29055 23103
rect 28997 23063 29055 23069
rect 29086 23060 29092 23112
rect 29144 23100 29150 23112
rect 29362 23100 29368 23112
rect 29144 23072 29368 23100
rect 29144 23060 29150 23072
rect 29362 23060 29368 23072
rect 29420 23060 29426 23112
rect 31202 23060 31208 23112
rect 31260 23100 31266 23112
rect 31297 23103 31355 23109
rect 31297 23100 31309 23103
rect 31260 23072 31309 23100
rect 31260 23060 31266 23072
rect 31297 23069 31309 23072
rect 31343 23069 31355 23103
rect 31297 23063 31355 23069
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23100 35311 23103
rect 35342 23100 35348 23112
rect 35299 23072 35348 23100
rect 35299 23069 35311 23072
rect 35253 23063 35311 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 22511 23004 23244 23032
rect 22511 23001 22523 23004
rect 22465 22995 22523 23001
rect 24762 22992 24768 23044
rect 24820 23032 24826 23044
rect 25685 23035 25743 23041
rect 24820 23004 24865 23032
rect 24820 22992 24826 23004
rect 25685 23001 25697 23035
rect 25731 23032 25743 23035
rect 26050 23032 26056 23044
rect 25731 23004 26056 23032
rect 25731 23001 25743 23004
rect 25685 22995 25743 23001
rect 16632 22936 16896 22964
rect 21085 22967 21143 22973
rect 16632 22924 16638 22936
rect 21085 22933 21097 22967
rect 21131 22964 21143 22967
rect 21910 22964 21916 22976
rect 21131 22936 21916 22964
rect 21131 22933 21143 22936
rect 21085 22927 21143 22933
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 25406 22924 25412 22976
rect 25464 22964 25470 22976
rect 25700 22964 25728 22995
rect 26050 22992 26056 23004
rect 26108 22992 26114 23044
rect 26694 22992 26700 23044
rect 26752 23032 26758 23044
rect 29822 23032 29828 23044
rect 26752 23004 27476 23032
rect 26752 22992 26758 23004
rect 26234 22964 26240 22976
rect 25464 22936 25728 22964
rect 26195 22936 26240 22964
rect 25464 22924 25470 22936
rect 26234 22924 26240 22936
rect 26292 22924 26298 22976
rect 27157 22967 27215 22973
rect 27157 22933 27169 22967
rect 27203 22964 27215 22967
rect 27338 22964 27344 22976
rect 27203 22936 27344 22964
rect 27203 22933 27215 22936
rect 27157 22927 27215 22933
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 27448 22964 27476 23004
rect 28368 23004 29828 23032
rect 28368 22964 28396 23004
rect 29822 22992 29828 23004
rect 29880 22992 29886 23044
rect 29917 23035 29975 23041
rect 29917 23001 29929 23035
rect 29963 23001 29975 23035
rect 29917 22995 29975 23001
rect 30837 23035 30895 23041
rect 30837 23001 30849 23035
rect 30883 23032 30895 23035
rect 30926 23032 30932 23044
rect 30883 23004 30932 23032
rect 30883 23001 30895 23004
rect 30837 22995 30895 23001
rect 27448 22936 28396 22964
rect 28534 22924 28540 22976
rect 28592 22964 28598 22976
rect 29089 22967 29147 22973
rect 29089 22964 29101 22967
rect 28592 22936 29101 22964
rect 28592 22924 28598 22936
rect 29089 22933 29101 22936
rect 29135 22933 29147 22967
rect 29932 22964 29960 22995
rect 30926 22992 30932 23004
rect 30984 22992 30990 23044
rect 32030 23032 32036 23044
rect 31991 23004 32036 23032
rect 32030 22992 32036 23004
rect 32088 22992 32094 23044
rect 32125 23035 32183 23041
rect 32125 23001 32137 23035
rect 32171 23001 32183 23035
rect 33042 23032 33048 23044
rect 33003 23004 33048 23032
rect 32125 22995 32183 23001
rect 31389 22967 31447 22973
rect 31389 22964 31401 22967
rect 29932 22936 31401 22964
rect 29089 22927 29147 22933
rect 31389 22933 31401 22936
rect 31435 22933 31447 22967
rect 32140 22964 32168 22995
rect 33042 22992 33048 23004
rect 33100 22992 33106 23044
rect 33962 22964 33968 22976
rect 32140 22936 33968 22964
rect 31389 22927 31447 22933
rect 33962 22924 33968 22936
rect 34020 22924 34026 22976
rect 35069 22967 35127 22973
rect 35069 22933 35081 22967
rect 35115 22964 35127 22967
rect 38010 22964 38016 22976
rect 35115 22936 38016 22964
rect 35115 22933 35127 22936
rect 35069 22927 35127 22933
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 13722 22760 13728 22772
rect 12406 22732 13728 22760
rect 7742 22692 7748 22704
rect 7703 22664 7748 22692
rect 7742 22652 7748 22664
rect 7800 22652 7806 22704
rect 10226 22692 10232 22704
rect 10187 22664 10232 22692
rect 10226 22652 10232 22664
rect 10284 22652 10290 22704
rect 10594 22652 10600 22704
rect 10652 22692 10658 22704
rect 11149 22695 11207 22701
rect 10652 22664 11008 22692
rect 10652 22652 10658 22664
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 7561 22559 7619 22565
rect 7561 22525 7573 22559
rect 7607 22556 7619 22559
rect 8386 22556 8392 22568
rect 7607 22528 8392 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 8386 22516 8392 22528
rect 8444 22516 8450 22568
rect 9398 22556 9404 22568
rect 9359 22528 9404 22556
rect 9398 22516 9404 22528
rect 9456 22516 9462 22568
rect 10134 22556 10140 22568
rect 10095 22528 10140 22556
rect 10134 22516 10140 22528
rect 10192 22516 10198 22568
rect 10980 22556 11008 22664
rect 11149 22661 11161 22695
rect 11195 22692 11207 22695
rect 11238 22692 11244 22704
rect 11195 22664 11244 22692
rect 11195 22661 11207 22664
rect 11149 22655 11207 22661
rect 11238 22652 11244 22664
rect 11296 22652 11302 22704
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22624 12127 22627
rect 12406 22624 12434 22732
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 14936 22732 15792 22760
rect 13354 22692 13360 22704
rect 13315 22664 13360 22692
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 12115 22596 12434 22624
rect 12529 22627 12587 22633
rect 12115 22593 12127 22596
rect 12069 22587 12127 22593
rect 12529 22593 12541 22627
rect 12575 22624 12587 22627
rect 12986 22624 12992 22636
rect 12575 22596 12992 22624
rect 12575 22593 12587 22596
rect 12529 22587 12587 22593
rect 12986 22584 12992 22596
rect 13044 22584 13050 22636
rect 14936 22624 14964 22732
rect 15102 22692 15108 22704
rect 15063 22664 15108 22692
rect 15102 22652 15108 22664
rect 15160 22652 15166 22704
rect 15197 22695 15255 22701
rect 15197 22661 15209 22695
rect 15243 22692 15255 22695
rect 15654 22692 15660 22704
rect 15243 22664 15660 22692
rect 15243 22661 15255 22664
rect 15197 22655 15255 22661
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 15764 22692 15792 22732
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 19613 22763 19671 22769
rect 19613 22760 19625 22763
rect 19484 22732 19625 22760
rect 19484 22720 19490 22732
rect 19613 22729 19625 22732
rect 19659 22729 19671 22763
rect 19613 22723 19671 22729
rect 19978 22720 19984 22772
rect 20036 22760 20042 22772
rect 20257 22763 20315 22769
rect 20257 22760 20269 22763
rect 20036 22732 20269 22760
rect 20036 22720 20042 22732
rect 20257 22729 20269 22732
rect 20303 22729 20315 22763
rect 20257 22723 20315 22729
rect 24486 22720 24492 22772
rect 24544 22760 24550 22772
rect 29270 22760 29276 22772
rect 24544 22732 29276 22760
rect 24544 22720 24550 22732
rect 29270 22720 29276 22732
rect 29328 22720 29334 22772
rect 29638 22720 29644 22772
rect 29696 22760 29702 22772
rect 29914 22760 29920 22772
rect 29696 22732 29920 22760
rect 29696 22720 29702 22732
rect 29914 22720 29920 22732
rect 29972 22760 29978 22772
rect 31662 22760 31668 22772
rect 29972 22732 31668 22760
rect 29972 22720 29978 22732
rect 31662 22720 31668 22732
rect 31720 22720 31726 22772
rect 37918 22760 37924 22772
rect 32324 22732 37924 22760
rect 20622 22692 20628 22704
rect 15764 22664 20628 22692
rect 20622 22652 20628 22664
rect 20680 22652 20686 22704
rect 22465 22695 22523 22701
rect 22465 22661 22477 22695
rect 22511 22692 22523 22695
rect 23474 22692 23480 22704
rect 22511 22664 23480 22692
rect 22511 22661 22523 22664
rect 22465 22655 22523 22661
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 24213 22695 24271 22701
rect 24213 22661 24225 22695
rect 24259 22692 24271 22695
rect 24946 22692 24952 22704
rect 24259 22664 24952 22692
rect 24259 22661 24271 22664
rect 24213 22655 24271 22661
rect 24946 22652 24952 22664
rect 25004 22652 25010 22704
rect 25130 22652 25136 22704
rect 25188 22692 25194 22704
rect 27338 22692 27344 22704
rect 25188 22664 26280 22692
rect 27299 22664 27344 22692
rect 25188 22652 25194 22664
rect 17218 22624 17224 22636
rect 14200 22596 14964 22624
rect 17179 22596 17224 22624
rect 13265 22559 13323 22565
rect 13265 22556 13277 22559
rect 10980 22528 13277 22556
rect 13265 22525 13277 22528
rect 13311 22556 13323 22559
rect 14200 22556 14228 22596
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 18322 22624 18328 22636
rect 18283 22596 18328 22624
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 19518 22624 19524 22636
rect 19479 22596 19524 22624
rect 19518 22584 19524 22596
rect 19576 22584 19582 22636
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22624 20223 22627
rect 21358 22624 21364 22636
rect 20211 22596 21364 22624
rect 20211 22593 20223 22596
rect 20165 22587 20223 22593
rect 21358 22584 21364 22596
rect 21416 22584 21422 22636
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 26252 22633 26280 22664
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 28534 22692 28540 22704
rect 28495 22664 28540 22692
rect 28534 22652 28540 22664
rect 28592 22652 28598 22704
rect 29457 22695 29515 22701
rect 29457 22661 29469 22695
rect 29503 22692 29515 22695
rect 29546 22692 29552 22704
rect 29503 22664 29552 22692
rect 29503 22661 29515 22664
rect 29457 22655 29515 22661
rect 29546 22652 29552 22664
rect 29604 22692 29610 22704
rect 29822 22692 29828 22704
rect 29604 22664 29828 22692
rect 29604 22652 29610 22664
rect 29822 22652 29828 22664
rect 29880 22652 29886 22704
rect 30193 22695 30251 22701
rect 30193 22661 30205 22695
rect 30239 22692 30251 22695
rect 31018 22692 31024 22704
rect 30239 22664 31024 22692
rect 30239 22661 30251 22664
rect 30193 22655 30251 22661
rect 31018 22652 31024 22664
rect 31076 22652 31082 22704
rect 31113 22695 31171 22701
rect 31113 22661 31125 22695
rect 31159 22692 31171 22695
rect 32214 22692 32220 22704
rect 31159 22664 32220 22692
rect 31159 22661 31171 22664
rect 31113 22655 31171 22661
rect 32214 22652 32220 22664
rect 32272 22652 32278 22704
rect 32324 22633 32352 22732
rect 37918 22720 37924 22732
rect 37976 22720 37982 22772
rect 38102 22692 38108 22704
rect 32968 22664 38108 22692
rect 32968 22633 32996 22664
rect 38102 22652 38108 22664
rect 38160 22652 38166 22704
rect 25593 22627 25651 22633
rect 25593 22624 25605 22627
rect 25556 22596 25605 22624
rect 25556 22584 25562 22596
rect 25593 22593 25605 22596
rect 25639 22593 25651 22627
rect 25593 22587 25651 22593
rect 26237 22627 26295 22633
rect 26237 22593 26249 22627
rect 26283 22593 26295 22627
rect 26237 22587 26295 22593
rect 31573 22627 31631 22633
rect 31573 22593 31585 22627
rect 31619 22593 31631 22627
rect 31573 22587 31631 22593
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 32953 22627 33011 22633
rect 32953 22593 32965 22627
rect 32999 22593 33011 22627
rect 32953 22587 33011 22593
rect 34885 22627 34943 22633
rect 34885 22593 34897 22627
rect 34931 22624 34943 22627
rect 35342 22624 35348 22636
rect 34931 22596 35348 22624
rect 34931 22593 34943 22596
rect 34885 22587 34943 22593
rect 13311 22528 14228 22556
rect 14277 22559 14335 22565
rect 13311 22525 13323 22528
rect 13265 22519 13323 22525
rect 14277 22525 14289 22559
rect 14323 22556 14335 22559
rect 15194 22556 15200 22568
rect 14323 22528 15200 22556
rect 14323 22525 14335 22528
rect 14277 22519 14335 22525
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 16117 22559 16175 22565
rect 16117 22525 16129 22559
rect 16163 22556 16175 22559
rect 21266 22556 21272 22568
rect 16163 22528 21272 22556
rect 16163 22525 16175 22528
rect 16117 22519 16175 22525
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 22370 22556 22376 22568
rect 22331 22528 22376 22556
rect 22370 22516 22376 22528
rect 22428 22516 22434 22568
rect 22554 22516 22560 22568
rect 22612 22556 22618 22568
rect 22649 22559 22707 22565
rect 22649 22556 22661 22559
rect 22612 22528 22661 22556
rect 22612 22516 22618 22528
rect 22649 22525 22661 22528
rect 22695 22525 22707 22559
rect 22649 22519 22707 22525
rect 24121 22559 24179 22565
rect 24121 22525 24133 22559
rect 24167 22556 24179 22559
rect 25038 22556 25044 22568
rect 24167 22528 25044 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 25038 22516 25044 22528
rect 25096 22516 25102 22568
rect 25133 22559 25191 22565
rect 25133 22525 25145 22559
rect 25179 22525 25191 22559
rect 27246 22556 27252 22568
rect 27207 22528 27252 22556
rect 25133 22519 25191 22525
rect 7834 22448 7840 22500
rect 7892 22488 7898 22500
rect 21174 22488 21180 22500
rect 7892 22460 21180 22488
rect 7892 22448 7898 22460
rect 21174 22448 21180 22460
rect 21232 22448 21238 22500
rect 22094 22488 22100 22500
rect 21284 22460 22100 22488
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 5534 22420 5540 22432
rect 1627 22392 5540 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 10318 22380 10324 22432
rect 10376 22420 10382 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 10376 22392 11897 22420
rect 10376 22380 10382 22392
rect 11885 22389 11897 22392
rect 11931 22389 11943 22423
rect 11885 22383 11943 22389
rect 12158 22380 12164 22432
rect 12216 22420 12222 22432
rect 12621 22423 12679 22429
rect 12621 22420 12633 22423
rect 12216 22392 12633 22420
rect 12216 22380 12222 22392
rect 12621 22389 12633 22392
rect 12667 22389 12679 22423
rect 12621 22383 12679 22389
rect 17313 22423 17371 22429
rect 17313 22389 17325 22423
rect 17359 22420 17371 22423
rect 17862 22420 17868 22432
rect 17359 22392 17868 22420
rect 17359 22389 17371 22392
rect 17313 22383 17371 22389
rect 17862 22380 17868 22392
rect 17920 22380 17926 22432
rect 18138 22380 18144 22432
rect 18196 22420 18202 22432
rect 18417 22423 18475 22429
rect 18417 22420 18429 22423
rect 18196 22392 18429 22420
rect 18196 22380 18202 22392
rect 18417 22389 18429 22392
rect 18463 22389 18475 22423
rect 18417 22383 18475 22389
rect 19058 22380 19064 22432
rect 19116 22420 19122 22432
rect 21284 22420 21312 22460
rect 22094 22448 22100 22460
rect 22152 22448 22158 22500
rect 25148 22488 25176 22519
rect 27246 22516 27252 22528
rect 27304 22516 27310 22568
rect 27430 22516 27436 22568
rect 27488 22556 27494 22568
rect 27525 22559 27583 22565
rect 27525 22556 27537 22559
rect 27488 22528 27537 22556
rect 27488 22516 27494 22528
rect 27525 22525 27537 22528
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 28445 22559 28503 22565
rect 28445 22525 28457 22559
rect 28491 22525 28503 22559
rect 28445 22519 28503 22525
rect 30101 22559 30159 22565
rect 30101 22525 30113 22559
rect 30147 22525 30159 22559
rect 30101 22519 30159 22525
rect 28460 22488 28488 22519
rect 29914 22488 29920 22500
rect 25148 22460 28396 22488
rect 28460 22460 29920 22488
rect 19116 22392 21312 22420
rect 19116 22380 19122 22392
rect 25130 22380 25136 22432
rect 25188 22420 25194 22432
rect 25685 22423 25743 22429
rect 25685 22420 25697 22423
rect 25188 22392 25697 22420
rect 25188 22380 25194 22392
rect 25685 22389 25697 22392
rect 25731 22389 25743 22423
rect 26326 22420 26332 22432
rect 26287 22392 26332 22420
rect 25685 22383 25743 22389
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 28368 22420 28396 22460
rect 29914 22448 29920 22460
rect 29972 22488 29978 22500
rect 30116 22488 30144 22519
rect 30742 22516 30748 22568
rect 30800 22556 30806 22568
rect 31478 22556 31484 22568
rect 30800 22528 31484 22556
rect 30800 22516 30806 22528
rect 31478 22516 31484 22528
rect 31536 22556 31542 22568
rect 31588 22556 31616 22587
rect 35342 22584 35348 22596
rect 35400 22584 35406 22636
rect 38010 22624 38016 22636
rect 37971 22596 38016 22624
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 31536 22528 31616 22556
rect 31536 22516 31542 22528
rect 31662 22516 31668 22568
rect 31720 22556 31726 22568
rect 34606 22556 34612 22568
rect 31720 22528 34612 22556
rect 31720 22516 31726 22528
rect 34606 22516 34612 22528
rect 34664 22516 34670 22568
rect 29972 22460 30144 22488
rect 29972 22448 29978 22460
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 33045 22491 33103 22497
rect 33045 22488 33057 22491
rect 30432 22460 33057 22488
rect 30432 22448 30438 22460
rect 33045 22457 33057 22460
rect 33091 22457 33103 22491
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 33045 22451 33103 22457
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 30742 22420 30748 22432
rect 28368 22392 30748 22420
rect 30742 22380 30748 22392
rect 30800 22380 30806 22432
rect 30926 22380 30932 22432
rect 30984 22420 30990 22432
rect 31665 22423 31723 22429
rect 31665 22420 31677 22423
rect 30984 22392 31677 22420
rect 30984 22380 30990 22392
rect 31665 22389 31677 22392
rect 31711 22389 31723 22423
rect 31665 22383 31723 22389
rect 32306 22380 32312 22432
rect 32364 22420 32370 22432
rect 32401 22423 32459 22429
rect 32401 22420 32413 22423
rect 32364 22392 32413 22420
rect 32364 22380 32370 22392
rect 32401 22389 32413 22392
rect 32447 22389 32459 22423
rect 32401 22383 32459 22389
rect 33134 22380 33140 22432
rect 33192 22420 33198 22432
rect 34977 22423 35035 22429
rect 34977 22420 34989 22423
rect 33192 22392 34989 22420
rect 33192 22380 33198 22392
rect 34977 22389 34989 22392
rect 35023 22389 35035 22423
rect 34977 22383 35035 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 8386 22216 8392 22228
rect 8299 22188 8392 22216
rect 8386 22176 8392 22188
rect 8444 22216 8450 22228
rect 17402 22216 17408 22228
rect 8444 22188 17408 22216
rect 8444 22176 8450 22188
rect 17402 22176 17408 22188
rect 17460 22216 17466 22228
rect 18230 22216 18236 22228
rect 17460 22188 18236 22216
rect 17460 22176 17466 22188
rect 18230 22176 18236 22188
rect 18288 22176 18294 22228
rect 18322 22176 18328 22228
rect 18380 22216 18386 22228
rect 20254 22216 20260 22228
rect 18380 22188 20260 22216
rect 18380 22176 18386 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 21100 22188 23612 22216
rect 1946 22108 1952 22160
rect 2004 22148 2010 22160
rect 8202 22148 8208 22160
rect 2004 22120 8208 22148
rect 2004 22108 2010 22120
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 11698 22108 11704 22160
rect 11756 22148 11762 22160
rect 12342 22148 12348 22160
rect 11756 22120 12348 22148
rect 11756 22108 11762 22120
rect 12342 22108 12348 22120
rect 12400 22108 12406 22160
rect 12894 22148 12900 22160
rect 12728 22120 12900 22148
rect 7469 22083 7527 22089
rect 1596 22052 2774 22080
rect 1596 22021 1624 22052
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 21981 1639 22015
rect 1581 21975 1639 21981
rect 1762 21876 1768 21888
rect 1723 21848 1768 21876
rect 1762 21836 1768 21848
rect 1820 21836 1826 21888
rect 2746 21876 2774 22052
rect 7469 22049 7481 22083
rect 7515 22080 7527 22083
rect 9950 22080 9956 22092
rect 7515 22052 9956 22080
rect 7515 22049 7527 22052
rect 7469 22043 7527 22049
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 12728 22089 12756 22120
rect 12894 22108 12900 22120
rect 12952 22148 12958 22160
rect 16942 22148 16948 22160
rect 12952 22120 16948 22148
rect 12952 22108 12958 22120
rect 16942 22108 16948 22120
rect 17000 22108 17006 22160
rect 17696 22120 20392 22148
rect 12713 22083 12771 22089
rect 10192 22052 10237 22080
rect 10192 22040 10198 22052
rect 12713 22049 12725 22083
rect 12759 22049 12771 22083
rect 12713 22043 12771 22049
rect 13814 22040 13820 22092
rect 13872 22080 13878 22092
rect 14458 22080 14464 22092
rect 13872 22052 14464 22080
rect 13872 22040 13878 22052
rect 14458 22040 14464 22052
rect 14516 22040 14522 22092
rect 15105 22083 15163 22089
rect 15105 22049 15117 22083
rect 15151 22080 15163 22083
rect 15194 22080 15200 22092
rect 15151 22052 15200 22080
rect 15151 22049 15163 22052
rect 15105 22043 15163 22049
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15749 22083 15807 22089
rect 15749 22049 15761 22083
rect 15795 22080 15807 22083
rect 15795 22052 16988 22080
rect 15795 22049 15807 22052
rect 15749 22043 15807 22049
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 5592 21984 7389 22012
rect 5592 21972 5598 21984
rect 7377 21981 7389 21984
rect 7423 21981 7435 22015
rect 7377 21975 7435 21981
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 22012 8355 22015
rect 8478 22012 8484 22024
rect 8343 21984 8484 22012
rect 8343 21981 8355 21984
rect 8297 21975 8355 21981
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 12986 21972 12992 22024
rect 13044 22012 13050 22024
rect 13446 22012 13452 22024
rect 13044 21984 13452 22012
rect 13044 21972 13050 21984
rect 13446 21972 13452 21984
rect 13504 22012 13510 22024
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 13504 21984 13553 22012
rect 13504 21972 13510 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 10134 21904 10140 21956
rect 10192 21944 10198 21956
rect 10229 21947 10287 21953
rect 10229 21944 10241 21947
rect 10192 21916 10241 21944
rect 10192 21904 10198 21916
rect 10229 21913 10241 21916
rect 10275 21913 10287 21947
rect 11146 21944 11152 21956
rect 11107 21916 11152 21944
rect 10229 21907 10287 21913
rect 11146 21904 11152 21916
rect 11204 21904 11210 21956
rect 11698 21944 11704 21956
rect 11659 21916 11704 21944
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 11790 21904 11796 21956
rect 11848 21944 11854 21956
rect 11848 21916 11893 21944
rect 11848 21904 11854 21916
rect 13078 21904 13084 21956
rect 13136 21944 13142 21956
rect 14384 21944 14412 21975
rect 13136 21916 14412 21944
rect 15197 21947 15255 21953
rect 13136 21904 13142 21916
rect 15197 21913 15209 21947
rect 15243 21913 15255 21947
rect 16298 21944 16304 21956
rect 16259 21916 16304 21944
rect 15197 21907 15255 21913
rect 10318 21876 10324 21888
rect 2746 21848 10324 21876
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 13633 21879 13691 21885
rect 13633 21845 13645 21879
rect 13679 21876 13691 21879
rect 13814 21876 13820 21888
rect 13679 21848 13820 21876
rect 13679 21845 13691 21848
rect 13633 21839 13691 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14461 21879 14519 21885
rect 14461 21845 14473 21879
rect 14507 21876 14519 21879
rect 15212 21876 15240 21907
rect 16298 21904 16304 21916
rect 16356 21904 16362 21956
rect 16393 21947 16451 21953
rect 16393 21913 16405 21947
rect 16439 21944 16451 21947
rect 16758 21944 16764 21956
rect 16439 21916 16764 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 16960 21953 16988 22052
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 17696 22080 17724 22120
rect 17368 22052 17724 22080
rect 18785 22083 18843 22089
rect 17368 22040 17374 22052
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 19886 22080 19892 22092
rect 18831 22052 19892 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 20364 22080 20392 22120
rect 20441 22083 20499 22089
rect 20441 22080 20453 22083
rect 20364 22052 20453 22080
rect 20441 22049 20453 22052
rect 20487 22080 20499 22083
rect 21100 22080 21128 22188
rect 21174 22108 21180 22160
rect 21232 22148 21238 22160
rect 23474 22148 23480 22160
rect 21232 22120 23480 22148
rect 21232 22108 21238 22120
rect 23474 22108 23480 22120
rect 23532 22108 23538 22160
rect 23584 22148 23612 22188
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 33134 22216 33140 22228
rect 23808 22188 33140 22216
rect 23808 22176 23814 22188
rect 33134 22176 33140 22188
rect 33192 22176 33198 22228
rect 27246 22148 27252 22160
rect 23584 22120 27252 22148
rect 27246 22108 27252 22120
rect 27304 22108 27310 22160
rect 29638 22148 29644 22160
rect 27908 22120 29644 22148
rect 23566 22080 23572 22092
rect 20487 22052 21128 22080
rect 23527 22052 23572 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 25958 22080 25964 22092
rect 25919 22052 25964 22080
rect 25958 22040 25964 22052
rect 26016 22040 26022 22092
rect 26050 22040 26056 22092
rect 26108 22080 26114 22092
rect 27908 22089 27936 22120
rect 29638 22108 29644 22120
rect 29696 22108 29702 22160
rect 32306 22108 32312 22160
rect 32364 22108 32370 22160
rect 38105 22151 38163 22157
rect 38105 22117 38117 22151
rect 38151 22117 38163 22151
rect 38105 22111 38163 22117
rect 27893 22083 27951 22089
rect 26108 22052 27844 22080
rect 26108 22040 26114 22052
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19705 22015 19763 22021
rect 19705 22012 19717 22015
rect 19484 21984 19717 22012
rect 19484 21972 19490 21984
rect 19705 21981 19717 21984
rect 19751 21981 19763 22015
rect 19705 21975 19763 21981
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 22012 22707 22015
rect 22738 22012 22744 22024
rect 22695 21984 22744 22012
rect 22695 21981 22707 21984
rect 22649 21975 22707 21981
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 23477 22015 23535 22021
rect 23477 21981 23489 22015
rect 23523 22012 23535 22015
rect 23842 22012 23848 22024
rect 23523 21984 23848 22012
rect 23523 21981 23535 21984
rect 23477 21975 23535 21981
rect 23842 21972 23848 21984
rect 23900 21972 23906 22024
rect 27816 22012 27844 22052
rect 27893 22049 27905 22083
rect 27939 22049 27951 22083
rect 27893 22043 27951 22049
rect 28442 22040 28448 22092
rect 28500 22080 28506 22092
rect 30374 22080 30380 22092
rect 28500 22052 30380 22080
rect 28500 22040 28506 22052
rect 30374 22040 30380 22052
rect 30432 22040 30438 22092
rect 30837 22083 30895 22089
rect 30837 22049 30849 22083
rect 30883 22080 30895 22083
rect 32324 22080 32352 22108
rect 33778 22080 33784 22092
rect 30883 22052 32352 22080
rect 33739 22052 33784 22080
rect 30883 22049 30895 22052
rect 30837 22043 30895 22049
rect 33778 22040 33784 22052
rect 33836 22040 33842 22092
rect 34514 22040 34520 22092
rect 34572 22080 34578 22092
rect 38120 22080 38148 22111
rect 34572 22052 38148 22080
rect 34572 22040 34578 22052
rect 27816 21984 28304 22012
rect 16945 21947 17003 21953
rect 16945 21913 16957 21947
rect 16991 21944 17003 21947
rect 17402 21944 17408 21956
rect 16991 21916 17408 21944
rect 16991 21913 17003 21916
rect 16945 21907 17003 21913
rect 17402 21904 17408 21916
rect 17460 21904 17466 21956
rect 17773 21947 17831 21953
rect 17773 21913 17785 21947
rect 17819 21913 17831 21947
rect 17773 21907 17831 21913
rect 14507 21848 15240 21876
rect 17788 21876 17816 21907
rect 17862 21904 17868 21956
rect 17920 21944 17926 21956
rect 19797 21947 19855 21953
rect 17920 21916 17965 21944
rect 17920 21904 17926 21916
rect 19797 21913 19809 21947
rect 19843 21944 19855 21947
rect 20533 21947 20591 21953
rect 20533 21944 20545 21947
rect 19843 21916 20545 21944
rect 19843 21913 19855 21916
rect 19797 21907 19855 21913
rect 20533 21913 20545 21916
rect 20579 21913 20591 21947
rect 20533 21907 20591 21913
rect 21085 21947 21143 21953
rect 21085 21913 21097 21947
rect 21131 21944 21143 21947
rect 21266 21944 21272 21956
rect 21131 21916 21272 21944
rect 21131 21913 21143 21916
rect 21085 21907 21143 21913
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 25130 21944 25136 21956
rect 25091 21916 25136 21944
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 25222 21904 25228 21956
rect 25280 21944 25286 21956
rect 25280 21916 25325 21944
rect 25280 21904 25286 21916
rect 25498 21904 25504 21956
rect 25556 21944 25562 21956
rect 26326 21944 26332 21956
rect 25556 21916 26332 21944
rect 25556 21904 25562 21916
rect 26326 21904 26332 21916
rect 26384 21904 26390 21956
rect 26878 21944 26884 21956
rect 26839 21916 26884 21944
rect 26878 21904 26884 21916
rect 26936 21904 26942 21956
rect 26973 21947 27031 21953
rect 26973 21913 26985 21947
rect 27019 21944 27031 21947
rect 27522 21944 27528 21956
rect 27019 21916 27528 21944
rect 27019 21913 27031 21916
rect 26973 21907 27031 21913
rect 27522 21904 27528 21916
rect 27580 21904 27586 21956
rect 28276 21944 28304 21984
rect 31754 21972 31760 22024
rect 31812 22012 31818 22024
rect 32214 22012 32220 22024
rect 31812 21984 32220 22012
rect 31812 21972 31818 21984
rect 32214 21972 32220 21984
rect 32272 21972 32278 22024
rect 32309 22015 32367 22021
rect 32309 21981 32321 22015
rect 32355 22012 32367 22015
rect 32766 22012 32772 22024
rect 32355 21984 32772 22012
rect 32355 21981 32367 21984
rect 32309 21975 32367 21981
rect 32766 21972 32772 21984
rect 32824 21972 32830 22024
rect 33045 22015 33103 22021
rect 33045 21981 33057 22015
rect 33091 22012 33103 22015
rect 33689 22015 33747 22021
rect 33091 21984 33640 22012
rect 33091 21981 33103 21984
rect 33045 21975 33103 21981
rect 28442 21944 28448 21956
rect 28276 21916 28448 21944
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 28537 21947 28595 21953
rect 28537 21913 28549 21947
rect 28583 21944 28595 21947
rect 28902 21944 28908 21956
rect 28583 21916 28908 21944
rect 28583 21913 28595 21916
rect 28537 21907 28595 21913
rect 28902 21904 28908 21916
rect 28960 21904 28966 21956
rect 29089 21947 29147 21953
rect 29089 21913 29101 21947
rect 29135 21944 29147 21947
rect 29638 21944 29644 21956
rect 29135 21916 29644 21944
rect 29135 21913 29147 21916
rect 29089 21907 29147 21913
rect 29638 21904 29644 21916
rect 29696 21904 29702 21956
rect 30926 21904 30932 21956
rect 30984 21944 30990 21956
rect 31849 21947 31907 21953
rect 31849 21944 31861 21947
rect 30984 21916 31029 21944
rect 31726 21916 31861 21944
rect 30984 21904 30990 21916
rect 22278 21876 22284 21888
rect 17788 21848 22284 21876
rect 14507 21845 14519 21848
rect 14461 21839 14519 21845
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 22741 21879 22799 21885
rect 22741 21845 22753 21879
rect 22787 21876 22799 21879
rect 22922 21876 22928 21888
rect 22787 21848 22928 21876
rect 22787 21845 22799 21848
rect 22741 21839 22799 21845
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 27982 21836 27988 21888
rect 28040 21876 28046 21888
rect 29733 21879 29791 21885
rect 29733 21876 29745 21879
rect 28040 21848 29745 21876
rect 28040 21836 28046 21848
rect 29733 21845 29745 21848
rect 29779 21845 29791 21879
rect 29733 21839 29791 21845
rect 30006 21836 30012 21888
rect 30064 21876 30070 21888
rect 31726 21876 31754 21916
rect 31849 21913 31861 21916
rect 31895 21913 31907 21947
rect 31849 21907 31907 21913
rect 32490 21904 32496 21956
rect 32548 21944 32554 21956
rect 33137 21947 33195 21953
rect 33137 21944 33149 21947
rect 32548 21916 33149 21944
rect 32548 21904 32554 21916
rect 33137 21913 33149 21916
rect 33183 21913 33195 21947
rect 33137 21907 33195 21913
rect 32398 21876 32404 21888
rect 30064 21848 31754 21876
rect 32359 21848 32404 21876
rect 30064 21836 30070 21848
rect 32398 21836 32404 21848
rect 32456 21836 32462 21888
rect 33612 21876 33640 21984
rect 33689 21981 33701 22015
rect 33735 21981 33747 22015
rect 33689 21975 33747 21981
rect 35161 22015 35219 22021
rect 35161 21981 35173 22015
rect 35207 22012 35219 22015
rect 36354 22012 36360 22024
rect 35207 21984 36360 22012
rect 35207 21981 35219 21984
rect 35161 21975 35219 21981
rect 33704 21944 33732 21975
rect 36354 21972 36360 21984
rect 36412 21972 36418 22024
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 38010 21944 38016 21956
rect 33704 21916 38016 21944
rect 38010 21904 38016 21916
rect 38068 21904 38074 21956
rect 33870 21876 33876 21888
rect 33612 21848 33876 21876
rect 33870 21836 33876 21848
rect 33928 21836 33934 21888
rect 34977 21879 35035 21885
rect 34977 21845 34989 21879
rect 35023 21876 35035 21879
rect 36538 21876 36544 21888
rect 35023 21848 36544 21876
rect 35023 21845 35035 21848
rect 34977 21839 35035 21845
rect 36538 21836 36544 21848
rect 36596 21836 36602 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 11057 21675 11115 21681
rect 11057 21641 11069 21675
rect 11103 21672 11115 21675
rect 11698 21672 11704 21684
rect 11103 21644 11704 21672
rect 11103 21641 11115 21644
rect 11057 21635 11115 21641
rect 11698 21632 11704 21644
rect 11756 21632 11762 21684
rect 11790 21632 11796 21684
rect 11848 21672 11854 21684
rect 12437 21675 12495 21681
rect 12437 21672 12449 21675
rect 11848 21644 12449 21672
rect 11848 21632 11854 21644
rect 12437 21641 12449 21644
rect 12483 21641 12495 21675
rect 12437 21635 12495 21641
rect 15289 21675 15347 21681
rect 15289 21641 15301 21675
rect 15335 21672 15347 21675
rect 16298 21672 16304 21684
rect 15335 21644 16304 21672
rect 15335 21641 15347 21644
rect 15289 21635 15347 21641
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 16390 21632 16396 21684
rect 16448 21672 16454 21684
rect 19794 21672 19800 21684
rect 16448 21644 19800 21672
rect 16448 21632 16454 21644
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 20349 21675 20407 21681
rect 20349 21672 20361 21675
rect 20036 21644 20361 21672
rect 20036 21632 20042 21644
rect 20349 21641 20361 21644
rect 20395 21641 20407 21675
rect 20349 21635 20407 21641
rect 22097 21675 22155 21681
rect 22097 21641 22109 21675
rect 22143 21672 22155 21675
rect 22186 21672 22192 21684
rect 22143 21644 22192 21672
rect 22143 21641 22155 21644
rect 22097 21635 22155 21641
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 27062 21672 27068 21684
rect 22796 21644 27068 21672
rect 22796 21632 22802 21644
rect 27062 21632 27068 21644
rect 27120 21632 27126 21684
rect 27798 21672 27804 21684
rect 27759 21644 27804 21672
rect 27798 21632 27804 21644
rect 27856 21632 27862 21684
rect 33045 21675 33103 21681
rect 33045 21672 33057 21675
rect 28736 21644 33057 21672
rect 10686 21564 10692 21616
rect 10744 21604 10750 21616
rect 11146 21604 11152 21616
rect 10744 21576 11152 21604
rect 10744 21564 10750 21576
rect 11146 21564 11152 21576
rect 11204 21564 11210 21616
rect 12710 21604 12716 21616
rect 11716 21576 12716 21604
rect 11716 21548 11744 21576
rect 12710 21564 12716 21576
rect 12768 21564 12774 21616
rect 13081 21607 13139 21613
rect 13081 21573 13093 21607
rect 13127 21604 13139 21607
rect 13817 21607 13875 21613
rect 13817 21604 13829 21607
rect 13127 21576 13829 21604
rect 13127 21573 13139 21576
rect 13081 21567 13139 21573
rect 13817 21573 13829 21576
rect 13863 21573 13875 21607
rect 13817 21567 13875 21573
rect 14369 21607 14427 21613
rect 14369 21573 14381 21607
rect 14415 21604 14427 21607
rect 14642 21604 14648 21616
rect 14415 21576 14648 21604
rect 14415 21573 14427 21576
rect 14369 21567 14427 21573
rect 14642 21564 14648 21576
rect 14700 21564 14706 21616
rect 16025 21607 16083 21613
rect 16025 21573 16037 21607
rect 16071 21604 16083 21607
rect 16666 21604 16672 21616
rect 16071 21576 16672 21604
rect 16071 21573 16083 21576
rect 16025 21567 16083 21573
rect 16666 21564 16672 21576
rect 16724 21564 16730 21616
rect 17218 21604 17224 21616
rect 17179 21576 17224 21604
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 19061 21607 19119 21613
rect 19061 21573 19073 21607
rect 19107 21604 19119 21607
rect 19334 21604 19340 21616
rect 19107 21576 19340 21604
rect 19107 21573 19119 21576
rect 19061 21567 19119 21573
rect 19334 21564 19340 21576
rect 19392 21564 19398 21616
rect 21266 21604 21272 21616
rect 20180 21576 21272 21604
rect 10318 21536 10324 21548
rect 10279 21508 10324 21536
rect 10318 21496 10324 21508
rect 10376 21496 10382 21548
rect 10502 21496 10508 21548
rect 10560 21536 10566 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10560 21508 10977 21536
rect 10560 21496 10566 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 11698 21536 11704 21548
rect 11659 21508 11704 21536
rect 10965 21499 11023 21505
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21536 12403 21539
rect 12526 21536 12532 21548
rect 12391 21508 12532 21536
rect 12391 21505 12403 21508
rect 12345 21499 12403 21505
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21536 13047 21539
rect 13035 21508 13124 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13096 21480 13124 21508
rect 15930 21496 15936 21548
rect 15988 21536 15994 21548
rect 18325 21539 18383 21545
rect 15988 21508 16033 21536
rect 15988 21496 15994 21508
rect 18325 21505 18337 21539
rect 18371 21536 18383 21539
rect 18598 21536 18604 21548
rect 18371 21508 18604 21536
rect 18371 21505 18383 21508
rect 18325 21499 18383 21505
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21536 19027 21539
rect 19242 21536 19248 21548
rect 19015 21508 19248 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 19610 21536 19616 21548
rect 19571 21508 19616 21536
rect 19610 21496 19616 21508
rect 19668 21496 19674 21548
rect 20180 21536 20208 21576
rect 21266 21564 21272 21576
rect 21324 21564 21330 21616
rect 23566 21604 23572 21616
rect 22664 21576 23572 21604
rect 19720 21508 20208 21536
rect 20257 21539 20315 21545
rect 13078 21428 13084 21480
rect 13136 21428 13142 21480
rect 13725 21471 13783 21477
rect 13725 21468 13737 21471
rect 13188 21440 13737 21468
rect 10778 21360 10784 21412
rect 10836 21400 10842 21412
rect 11238 21400 11244 21412
rect 10836 21372 11244 21400
rect 10836 21360 10842 21372
rect 11238 21360 11244 21372
rect 11296 21400 11302 21412
rect 11296 21372 11913 21400
rect 11296 21360 11302 21372
rect 11790 21332 11796 21344
rect 11751 21304 11796 21332
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 11885 21332 11913 21372
rect 12066 21360 12072 21412
rect 12124 21400 12130 21412
rect 13188 21400 13216 21440
rect 13725 21437 13737 21440
rect 13771 21468 13783 21471
rect 14458 21468 14464 21480
rect 13771 21440 14464 21468
rect 13771 21437 13783 21440
rect 13725 21431 13783 21437
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 15838 21468 15844 21480
rect 15252 21440 15844 21468
rect 15252 21428 15258 21440
rect 15838 21428 15844 21440
rect 15896 21468 15902 21480
rect 17129 21471 17187 21477
rect 17129 21468 17141 21471
rect 15896 21440 17141 21468
rect 15896 21428 15902 21440
rect 17129 21437 17141 21440
rect 17175 21437 17187 21471
rect 17129 21431 17187 21437
rect 17402 21428 17408 21480
rect 17460 21468 17466 21480
rect 19720 21468 19748 21508
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20530 21536 20536 21548
rect 20303 21508 20536 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 20898 21536 20904 21548
rect 20859 21508 20904 21536
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 21818 21536 21824 21548
rect 21232 21508 21824 21536
rect 21232 21496 21238 21508
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22002 21536 22008 21548
rect 21963 21508 22008 21536
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22664 21545 22692 21576
rect 23566 21564 23572 21576
rect 23624 21564 23630 21616
rect 23661 21607 23719 21613
rect 23661 21573 23673 21607
rect 23707 21604 23719 21607
rect 23934 21604 23940 21616
rect 23707 21576 23940 21604
rect 23707 21573 23719 21576
rect 23661 21567 23719 21573
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 25225 21607 25283 21613
rect 25225 21573 25237 21607
rect 25271 21604 25283 21607
rect 25498 21604 25504 21616
rect 25271 21576 25504 21604
rect 25271 21573 25283 21576
rect 25225 21567 25283 21573
rect 25498 21564 25504 21576
rect 25556 21564 25562 21616
rect 28530 21607 28588 21613
rect 28530 21573 28542 21607
rect 28576 21604 28588 21607
rect 28736 21604 28764 21644
rect 33045 21641 33057 21644
rect 33091 21641 33103 21675
rect 33045 21635 33103 21641
rect 28576 21576 28764 21604
rect 28576 21573 28588 21576
rect 28530 21567 28588 21573
rect 28902 21564 28908 21616
rect 28960 21604 28966 21616
rect 29641 21607 29699 21613
rect 29641 21604 29653 21607
rect 28960 21576 29653 21604
rect 28960 21564 28966 21576
rect 29641 21573 29653 21576
rect 29687 21573 29699 21607
rect 29641 21567 29699 21573
rect 30098 21564 30104 21616
rect 30156 21604 30162 21616
rect 30745 21607 30803 21613
rect 30745 21604 30757 21607
rect 30156 21576 30757 21604
rect 30156 21564 30162 21576
rect 30745 21573 30757 21576
rect 30791 21573 30803 21607
rect 30745 21567 30803 21573
rect 30837 21607 30895 21613
rect 30837 21573 30849 21607
rect 30883 21604 30895 21607
rect 32398 21604 32404 21616
rect 30883 21576 32404 21604
rect 30883 21573 30895 21576
rect 30837 21567 30895 21573
rect 32398 21564 32404 21576
rect 32456 21564 32462 21616
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 27614 21536 27620 21548
rect 27575 21508 27620 21536
rect 22649 21499 22707 21505
rect 27614 21496 27620 21508
rect 27672 21496 27678 21548
rect 29546 21536 29552 21548
rect 29507 21508 29552 21536
rect 29546 21496 29552 21508
rect 29604 21496 29610 21548
rect 30558 21536 30564 21548
rect 29656 21508 30564 21536
rect 17460 21440 19748 21468
rect 17460 21428 17466 21440
rect 19886 21428 19892 21480
rect 19944 21468 19950 21480
rect 23569 21471 23627 21477
rect 19944 21440 23520 21468
rect 19944 21428 19950 21440
rect 12124 21372 13216 21400
rect 17681 21403 17739 21409
rect 12124 21360 12130 21372
rect 17681 21369 17693 21403
rect 17727 21400 17739 21403
rect 23492 21400 23520 21440
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 23750 21468 23756 21480
rect 23615 21440 23756 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 23750 21428 23756 21440
rect 23808 21428 23814 21480
rect 24118 21428 24124 21480
rect 24176 21468 24182 21480
rect 25130 21468 25136 21480
rect 24176 21440 24221 21468
rect 25091 21440 25136 21468
rect 24176 21428 24182 21440
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 25958 21468 25964 21480
rect 25919 21440 25964 21468
rect 25958 21428 25964 21440
rect 26016 21428 26022 21480
rect 28258 21428 28264 21480
rect 28316 21468 28322 21480
rect 28446 21471 28504 21477
rect 28316 21456 28396 21468
rect 28446 21456 28458 21471
rect 28316 21440 28458 21456
rect 28316 21428 28322 21440
rect 28368 21437 28458 21440
rect 28492 21437 28504 21471
rect 28368 21431 28504 21437
rect 28368 21428 28488 21431
rect 28626 21428 28632 21480
rect 28684 21456 28690 21480
rect 29656 21468 29684 21508
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 31846 21536 31852 21548
rect 31404 21508 31852 21536
rect 31021 21471 31079 21477
rect 31021 21468 31033 21471
rect 28736 21456 29684 21468
rect 28684 21440 29684 21456
rect 29840 21440 31033 21468
rect 28684 21428 28764 21440
rect 24854 21400 24860 21412
rect 17727 21372 23428 21400
rect 23492 21372 24860 21400
rect 17727 21369 17739 21372
rect 17681 21363 17739 21369
rect 17126 21332 17132 21344
rect 11885 21304 17132 21332
rect 17126 21292 17132 21304
rect 17184 21292 17190 21344
rect 18417 21335 18475 21341
rect 18417 21301 18429 21335
rect 18463 21332 18475 21335
rect 18874 21332 18880 21344
rect 18463 21304 18880 21332
rect 18463 21301 18475 21304
rect 18417 21295 18475 21301
rect 18874 21292 18880 21304
rect 18932 21292 18938 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19705 21335 19763 21341
rect 19705 21332 19717 21335
rect 19484 21304 19717 21332
rect 19484 21292 19490 21304
rect 19705 21301 19717 21304
rect 19751 21301 19763 21335
rect 19705 21295 19763 21301
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 20898 21332 20904 21344
rect 19852 21304 20904 21332
rect 19852 21292 19858 21304
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 20993 21335 21051 21341
rect 20993 21301 21005 21335
rect 21039 21332 21051 21335
rect 22186 21332 22192 21344
rect 21039 21304 22192 21332
rect 21039 21301 21051 21304
rect 20993 21295 21051 21301
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 22278 21292 22284 21344
rect 22336 21332 22342 21344
rect 22741 21335 22799 21341
rect 22741 21332 22753 21335
rect 22336 21304 22753 21332
rect 22336 21292 22342 21304
rect 22741 21301 22753 21304
rect 22787 21301 22799 21335
rect 23400 21332 23428 21372
rect 24854 21360 24860 21372
rect 24912 21360 24918 21412
rect 28997 21403 29055 21409
rect 28997 21369 29009 21403
rect 29043 21369 29055 21403
rect 28997 21363 29055 21369
rect 27430 21332 27436 21344
rect 23400 21304 27436 21332
rect 22741 21295 22799 21301
rect 27430 21292 27436 21304
rect 27488 21292 27494 21344
rect 28626 21292 28632 21344
rect 28684 21332 28690 21344
rect 29012 21332 29040 21363
rect 29638 21360 29644 21412
rect 29696 21400 29702 21412
rect 29840 21400 29868 21440
rect 31021 21437 31033 21440
rect 31067 21468 31079 21471
rect 31404 21468 31432 21508
rect 31846 21496 31852 21508
rect 31904 21496 31910 21548
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 32272 21508 32321 21536
rect 32272 21496 32278 21508
rect 32309 21505 32321 21508
rect 32355 21536 32367 21539
rect 32582 21536 32588 21548
rect 32355 21508 32588 21536
rect 32355 21505 32367 21508
rect 32309 21499 32367 21505
rect 32582 21496 32588 21508
rect 32640 21496 32646 21548
rect 32950 21536 32956 21548
rect 32911 21508 32956 21536
rect 32950 21496 32956 21508
rect 33008 21496 33014 21548
rect 33594 21536 33600 21548
rect 33555 21508 33600 21536
rect 33594 21496 33600 21508
rect 33652 21496 33658 21548
rect 34241 21539 34299 21545
rect 34241 21505 34253 21539
rect 34287 21536 34299 21539
rect 36354 21536 36360 21548
rect 34287 21508 36360 21536
rect 34287 21505 34299 21508
rect 34241 21499 34299 21505
rect 36354 21496 36360 21508
rect 36412 21496 36418 21548
rect 33689 21471 33747 21477
rect 33689 21468 33701 21471
rect 31067 21440 31432 21468
rect 31496 21440 33701 21468
rect 31067 21437 31079 21440
rect 31021 21431 31079 21437
rect 29696 21372 29868 21400
rect 29696 21360 29702 21372
rect 29914 21360 29920 21412
rect 29972 21400 29978 21412
rect 31496 21400 31524 21440
rect 33689 21437 33701 21440
rect 33735 21437 33747 21471
rect 33689 21431 33747 21437
rect 29972 21372 31524 21400
rect 29972 21360 29978 21372
rect 28684 21304 29040 21332
rect 28684 21292 28690 21304
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 32401 21335 32459 21341
rect 32401 21332 32413 21335
rect 30432 21304 32413 21332
rect 30432 21292 30438 21304
rect 32401 21301 32413 21304
rect 32447 21301 32459 21335
rect 32401 21295 32459 21301
rect 32490 21292 32496 21344
rect 32548 21332 32554 21344
rect 33410 21332 33416 21344
rect 32548 21304 33416 21332
rect 32548 21292 32554 21304
rect 33410 21292 33416 21304
rect 33468 21292 33474 21344
rect 34330 21332 34336 21344
rect 34291 21304 34336 21332
rect 34330 21292 34336 21304
rect 34388 21292 34394 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 10134 21088 10140 21140
rect 10192 21128 10198 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 10192 21100 13645 21128
rect 10192 21088 10198 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13633 21091 13691 21097
rect 14553 21131 14611 21137
rect 14553 21097 14565 21131
rect 14599 21128 14611 21131
rect 15378 21128 15384 21140
rect 14599 21100 15384 21128
rect 14599 21097 14611 21100
rect 14553 21091 14611 21097
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 17034 21128 17040 21140
rect 15764 21100 17040 21128
rect 12526 21020 12532 21072
rect 12584 21060 12590 21072
rect 12894 21060 12900 21072
rect 12584 21032 12900 21060
rect 12584 21020 12590 21032
rect 12894 21020 12900 21032
rect 12952 21020 12958 21072
rect 13446 21020 13452 21072
rect 13504 21060 13510 21072
rect 15764 21060 15792 21100
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 23934 21128 23940 21140
rect 17184 21100 23796 21128
rect 23895 21100 23940 21128
rect 17184 21088 17190 21100
rect 23768 21060 23796 21100
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 24673 21131 24731 21137
rect 24673 21097 24685 21131
rect 24719 21128 24731 21131
rect 24762 21128 24768 21140
rect 24719 21100 24768 21128
rect 24719 21097 24731 21100
rect 24673 21091 24731 21097
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 24946 21088 24952 21140
rect 25004 21128 25010 21140
rect 26142 21128 26148 21140
rect 25004 21100 26148 21128
rect 25004 21088 25010 21100
rect 26142 21088 26148 21100
rect 26200 21088 26206 21140
rect 27614 21088 27620 21140
rect 27672 21128 27678 21140
rect 37274 21128 37280 21140
rect 27672 21100 37280 21128
rect 27672 21088 27678 21100
rect 37274 21088 37280 21100
rect 37332 21088 37338 21140
rect 37918 21088 37924 21140
rect 37976 21128 37982 21140
rect 38105 21131 38163 21137
rect 38105 21128 38117 21131
rect 37976 21100 38117 21128
rect 37976 21088 37982 21100
rect 38105 21097 38117 21100
rect 38151 21097 38163 21131
rect 38105 21091 38163 21097
rect 24118 21060 24124 21072
rect 13504 21032 15792 21060
rect 15856 21032 22048 21060
rect 23768 21032 24124 21060
rect 13504 21020 13510 21032
rect 13630 20992 13636 21004
rect 12406 20964 13636 20992
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 6822 20924 6828 20936
rect 1627 20896 6828 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20924 12127 20927
rect 12406 20924 12434 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 15856 21001 15884 21032
rect 15841 20995 15899 21001
rect 15841 20992 15853 20995
rect 13740 20964 15853 20992
rect 12115 20896 12434 20924
rect 12115 20893 12127 20896
rect 12069 20887 12127 20893
rect 13446 20884 13452 20936
rect 13504 20924 13510 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13504 20896 13553 20924
rect 13504 20884 13510 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 10686 20816 10692 20868
rect 10744 20856 10750 20868
rect 10744 20828 12434 20856
rect 10744 20816 10750 20828
rect 1762 20788 1768 20800
rect 1723 20760 1768 20788
rect 1762 20748 1768 20760
rect 1820 20748 1826 20800
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 10502 20788 10508 20800
rect 4120 20760 10508 20788
rect 4120 20748 4126 20760
rect 10502 20748 10508 20760
rect 10560 20748 10566 20800
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 12161 20791 12219 20797
rect 12161 20788 12173 20791
rect 11204 20760 12173 20788
rect 11204 20748 11210 20760
rect 12161 20757 12173 20760
rect 12207 20757 12219 20791
rect 12406 20788 12434 20828
rect 13740 20788 13768 20964
rect 15841 20961 15853 20964
rect 15887 20961 15899 20995
rect 15841 20955 15899 20961
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 18046 20992 18052 21004
rect 17451 20964 18052 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 21818 20992 21824 21004
rect 18340 20964 21824 20992
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 14384 20896 14473 20924
rect 12406 20760 13768 20788
rect 12161 20751 12219 20757
rect 14090 20748 14096 20800
rect 14148 20788 14154 20800
rect 14384 20788 14412 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14734 20884 14740 20936
rect 14792 20924 14798 20936
rect 15105 20927 15163 20933
rect 15105 20924 15117 20927
rect 14792 20896 15117 20924
rect 14792 20884 14798 20896
rect 15105 20893 15117 20896
rect 15151 20893 15163 20927
rect 15105 20887 15163 20893
rect 15930 20816 15936 20868
rect 15988 20856 15994 20868
rect 16853 20859 16911 20865
rect 15988 20828 16033 20856
rect 15988 20816 15994 20828
rect 16853 20825 16865 20859
rect 16899 20856 16911 20859
rect 16899 20828 17448 20856
rect 16899 20825 16911 20828
rect 16853 20819 16911 20825
rect 14148 20760 14412 20788
rect 15197 20791 15255 20797
rect 14148 20748 14154 20760
rect 15197 20757 15209 20791
rect 15243 20788 15255 20791
rect 17034 20788 17040 20800
rect 15243 20760 17040 20788
rect 15243 20757 15255 20760
rect 15197 20751 15255 20757
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17420 20788 17448 20828
rect 17494 20816 17500 20868
rect 17552 20856 17558 20868
rect 17552 20828 17597 20856
rect 17552 20816 17558 20828
rect 17678 20816 17684 20868
rect 17736 20856 17742 20868
rect 18340 20856 18368 20964
rect 21818 20952 21824 20964
rect 21876 20952 21882 21004
rect 22020 20992 22048 21032
rect 24118 21020 24124 21032
rect 24176 21020 24182 21072
rect 27522 21020 27528 21072
rect 27580 21060 27586 21072
rect 29825 21063 29883 21069
rect 29825 21060 29837 21063
rect 27580 21032 29837 21060
rect 27580 21020 27586 21032
rect 29825 21029 29837 21032
rect 29871 21029 29883 21063
rect 30834 21060 30840 21072
rect 29825 21023 29883 21029
rect 30300 21032 30840 21060
rect 24302 20992 24308 21004
rect 22020 20964 24308 20992
rect 24302 20952 24308 20964
rect 24360 20952 24366 21004
rect 25130 20952 25136 21004
rect 25188 20992 25194 21004
rect 25501 20995 25559 21001
rect 25501 20992 25513 20995
rect 25188 20964 25513 20992
rect 25188 20952 25194 20964
rect 25501 20961 25513 20964
rect 25547 20961 25559 20995
rect 25501 20955 25559 20961
rect 25685 20995 25743 21001
rect 25685 20961 25697 20995
rect 25731 20992 25743 20995
rect 26234 20992 26240 21004
rect 25731 20964 26240 20992
rect 25731 20961 25743 20964
rect 25685 20955 25743 20961
rect 26234 20952 26240 20964
rect 26292 20952 26298 21004
rect 27982 20992 27988 21004
rect 27943 20964 27988 20992
rect 27982 20952 27988 20964
rect 28040 20952 28046 21004
rect 28258 20992 28264 21004
rect 28219 20964 28264 20992
rect 28258 20952 28264 20964
rect 28316 20992 28322 21004
rect 30190 20992 30196 21004
rect 28316 20964 30196 20992
rect 28316 20952 28322 20964
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20924 21511 20927
rect 21542 20924 21548 20936
rect 21499 20896 21548 20924
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20924 23903 20927
rect 23934 20924 23940 20936
rect 23891 20896 23940 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 23934 20884 23940 20896
rect 23992 20884 23998 20936
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20924 24639 20927
rect 24946 20924 24952 20936
rect 24627 20896 24952 20924
rect 24627 20893 24639 20896
rect 24581 20887 24639 20893
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 29178 20884 29184 20936
rect 29236 20924 29242 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29236 20896 29745 20924
rect 29236 20884 29242 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 17736 20828 18368 20856
rect 18417 20859 18475 20865
rect 17736 20816 17742 20828
rect 18417 20825 18429 20859
rect 18463 20825 18475 20859
rect 19886 20856 19892 20868
rect 19847 20828 19892 20856
rect 18417 20819 18475 20825
rect 17586 20788 17592 20800
rect 17420 20760 17592 20788
rect 17586 20748 17592 20760
rect 17644 20788 17650 20800
rect 18432 20788 18460 20819
rect 19886 20816 19892 20828
rect 19944 20816 19950 20868
rect 19978 20816 19984 20868
rect 20036 20856 20042 20868
rect 20036 20828 20081 20856
rect 20036 20816 20042 20828
rect 20806 20816 20812 20868
rect 20864 20856 20870 20868
rect 20901 20859 20959 20865
rect 20901 20856 20913 20859
rect 20864 20828 20913 20856
rect 20864 20816 20870 20828
rect 20901 20825 20913 20828
rect 20947 20856 20959 20859
rect 21082 20856 21088 20868
rect 20947 20828 21088 20856
rect 20947 20825 20959 20828
rect 20901 20819 20959 20825
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 21910 20816 21916 20868
rect 21968 20856 21974 20868
rect 22189 20859 22247 20865
rect 22189 20856 22201 20859
rect 21968 20828 22201 20856
rect 21968 20816 21974 20828
rect 22189 20825 22201 20828
rect 22235 20825 22247 20859
rect 22189 20819 22247 20825
rect 22278 20816 22284 20868
rect 22336 20856 22342 20868
rect 23201 20859 23259 20865
rect 22336 20828 22381 20856
rect 22336 20816 22342 20828
rect 23201 20825 23213 20859
rect 23247 20856 23259 20859
rect 23290 20856 23296 20868
rect 23247 20828 23296 20856
rect 23247 20825 23259 20828
rect 23201 20819 23259 20825
rect 23290 20816 23296 20828
rect 23348 20816 23354 20868
rect 27341 20859 27399 20865
rect 27341 20825 27353 20859
rect 27387 20825 27399 20859
rect 27341 20819 27399 20825
rect 17644 20760 18460 20788
rect 17644 20748 17650 20760
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 19150 20788 19156 20800
rect 18656 20760 19156 20788
rect 18656 20748 18662 20760
rect 19150 20748 19156 20760
rect 19208 20748 19214 20800
rect 19610 20748 19616 20800
rect 19668 20788 19674 20800
rect 20530 20788 20536 20800
rect 19668 20760 20536 20788
rect 19668 20748 19674 20760
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 21542 20788 21548 20800
rect 21503 20760 21548 20788
rect 21542 20748 21548 20760
rect 21600 20748 21606 20800
rect 21634 20748 21640 20800
rect 21692 20788 21698 20800
rect 25498 20788 25504 20800
rect 21692 20760 25504 20788
rect 21692 20748 21698 20760
rect 25498 20748 25504 20760
rect 25556 20748 25562 20800
rect 25682 20748 25688 20800
rect 25740 20788 25746 20800
rect 26326 20788 26332 20800
rect 25740 20760 26332 20788
rect 25740 20748 25746 20760
rect 26326 20748 26332 20760
rect 26384 20748 26390 20800
rect 27356 20788 27384 20819
rect 28074 20816 28080 20868
rect 28132 20856 28138 20868
rect 28132 20828 28177 20856
rect 28132 20816 28138 20828
rect 28626 20816 28632 20868
rect 28684 20856 28690 20868
rect 30006 20856 30012 20868
rect 28684 20828 30012 20856
rect 28684 20816 28690 20828
rect 30006 20816 30012 20828
rect 30064 20816 30070 20868
rect 30300 20788 30328 21032
rect 30834 21020 30840 21032
rect 30892 21020 30898 21072
rect 31021 21063 31079 21069
rect 31021 21029 31033 21063
rect 31067 21060 31079 21063
rect 31110 21060 31116 21072
rect 31067 21032 31116 21060
rect 31067 21029 31079 21032
rect 31021 21023 31079 21029
rect 31110 21020 31116 21032
rect 31168 21020 31174 21072
rect 31938 21020 31944 21072
rect 31996 21060 32002 21072
rect 35434 21060 35440 21072
rect 31996 21032 35440 21060
rect 31996 21020 32002 21032
rect 35434 21020 35440 21032
rect 35492 21020 35498 21072
rect 30469 20995 30527 21001
rect 30469 20961 30481 20995
rect 30515 20992 30527 20995
rect 30926 20992 30932 21004
rect 30515 20964 30932 20992
rect 30515 20961 30527 20964
rect 30469 20955 30527 20961
rect 30926 20952 30932 20964
rect 30984 20992 30990 21004
rect 31849 20995 31907 21001
rect 31849 20992 31861 20995
rect 30984 20964 31861 20992
rect 30984 20952 30990 20964
rect 31849 20961 31861 20964
rect 31895 20992 31907 20995
rect 34330 20992 34336 21004
rect 31895 20964 34336 20992
rect 31895 20961 31907 20964
rect 31849 20955 31907 20961
rect 34330 20952 34336 20964
rect 34388 20952 34394 21004
rect 32766 20884 32772 20936
rect 32824 20924 32830 20936
rect 32953 20927 33011 20933
rect 32953 20924 32965 20927
rect 32824 20896 32965 20924
rect 32824 20884 32830 20896
rect 32953 20893 32965 20896
rect 32999 20893 33011 20927
rect 32953 20887 33011 20893
rect 33226 20884 33232 20936
rect 33284 20924 33290 20936
rect 33597 20927 33655 20933
rect 33597 20924 33609 20927
rect 33284 20896 33609 20924
rect 33284 20884 33290 20896
rect 33597 20893 33609 20896
rect 33643 20893 33655 20927
rect 38286 20924 38292 20936
rect 38247 20896 38292 20924
rect 33597 20887 33655 20893
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 30561 20859 30619 20865
rect 30561 20825 30573 20859
rect 30607 20825 30619 20859
rect 30561 20819 30619 20825
rect 27356 20760 30328 20788
rect 30576 20788 30604 20819
rect 31938 20816 31944 20868
rect 31996 20856 32002 20868
rect 31996 20828 32041 20856
rect 31996 20816 32002 20828
rect 32214 20816 32220 20868
rect 32272 20856 32278 20868
rect 32490 20856 32496 20868
rect 32272 20828 32496 20856
rect 32272 20816 32278 20828
rect 32490 20816 32496 20828
rect 32548 20816 32554 20868
rect 33689 20859 33747 20865
rect 33689 20856 33701 20859
rect 32692 20828 33701 20856
rect 32692 20788 32720 20828
rect 33689 20825 33701 20828
rect 33735 20825 33747 20859
rect 33689 20819 33747 20825
rect 33870 20816 33876 20868
rect 33928 20856 33934 20868
rect 35894 20856 35900 20868
rect 33928 20828 35900 20856
rect 33928 20816 33934 20828
rect 35894 20816 35900 20828
rect 35952 20816 35958 20868
rect 33042 20788 33048 20800
rect 30576 20760 32720 20788
rect 33003 20760 33048 20788
rect 33042 20748 33048 20760
rect 33100 20748 33106 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6822 20584 6828 20596
rect 6783 20556 6828 20584
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 13725 20587 13783 20593
rect 13725 20584 13737 20587
rect 12860 20556 13737 20584
rect 12860 20544 12866 20556
rect 13725 20553 13737 20556
rect 13771 20553 13783 20587
rect 16209 20587 16267 20593
rect 13725 20547 13783 20553
rect 14384 20556 16160 20584
rect 13078 20516 13084 20528
rect 12406 20488 13084 20516
rect 1854 20408 1860 20460
rect 1912 20448 1918 20460
rect 1949 20451 2007 20457
rect 1949 20448 1961 20451
rect 1912 20420 1961 20448
rect 1912 20408 1918 20420
rect 1949 20417 1961 20420
rect 1995 20417 2007 20451
rect 1949 20411 2007 20417
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20448 7067 20451
rect 7558 20448 7564 20460
rect 7055 20420 7564 20448
rect 7055 20417 7067 20420
rect 7009 20411 7067 20417
rect 7558 20408 7564 20420
rect 7616 20408 7622 20460
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20448 12219 20451
rect 12406 20448 12434 20488
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 13262 20476 13268 20528
rect 13320 20516 13326 20528
rect 14384 20516 14412 20556
rect 13320 20488 14412 20516
rect 14461 20519 14519 20525
rect 13320 20476 13326 20488
rect 14461 20485 14473 20519
rect 14507 20516 14519 20519
rect 15286 20516 15292 20528
rect 14507 20488 15292 20516
rect 14507 20485 14519 20488
rect 14461 20479 14519 20485
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 16132 20516 16160 20556
rect 16209 20553 16221 20587
rect 16255 20584 16267 20587
rect 17218 20584 17224 20596
rect 16255 20556 17224 20584
rect 16255 20553 16267 20556
rect 16209 20547 16267 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20349 20587 20407 20593
rect 20349 20584 20361 20587
rect 20036 20556 20361 20584
rect 20036 20544 20042 20556
rect 20349 20553 20361 20556
rect 20395 20553 20407 20587
rect 20349 20547 20407 20553
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 21600 20556 24164 20584
rect 21600 20544 21606 20556
rect 16758 20516 16764 20528
rect 16132 20488 16764 20516
rect 16758 20476 16764 20488
rect 16816 20476 16822 20528
rect 17034 20516 17040 20528
rect 16995 20488 17040 20516
rect 17034 20476 17040 20488
rect 17092 20476 17098 20528
rect 18874 20516 18880 20528
rect 18835 20488 18880 20516
rect 18874 20476 18880 20488
rect 18932 20476 18938 20528
rect 22186 20516 22192 20528
rect 22147 20488 22192 20516
rect 22186 20476 22192 20488
rect 22244 20476 22250 20528
rect 22278 20476 22284 20528
rect 22336 20516 22342 20528
rect 22554 20516 22560 20528
rect 22336 20488 22560 20516
rect 22336 20476 22342 20488
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 23750 20476 23756 20528
rect 23808 20516 23814 20528
rect 24136 20525 24164 20556
rect 24210 20544 24216 20596
rect 24268 20584 24274 20596
rect 25406 20584 25412 20596
rect 24268 20556 25412 20584
rect 24268 20544 24274 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 25498 20544 25504 20596
rect 25556 20584 25562 20596
rect 29454 20584 29460 20596
rect 25556 20556 29460 20584
rect 25556 20544 25562 20556
rect 29454 20544 29460 20556
rect 29512 20544 29518 20596
rect 29730 20544 29736 20596
rect 29788 20584 29794 20596
rect 30006 20584 30012 20596
rect 29788 20556 30012 20584
rect 29788 20544 29794 20556
rect 30006 20544 30012 20556
rect 30064 20544 30070 20596
rect 30926 20544 30932 20596
rect 30984 20584 30990 20596
rect 31294 20584 31300 20596
rect 30984 20556 31300 20584
rect 30984 20544 30990 20556
rect 31294 20544 31300 20556
rect 31352 20544 31358 20596
rect 31570 20544 31576 20596
rect 31628 20584 31634 20596
rect 31628 20556 34836 20584
rect 31628 20544 31634 20556
rect 24029 20519 24087 20525
rect 24029 20516 24041 20519
rect 23808 20488 24041 20516
rect 23808 20476 23814 20488
rect 24029 20485 24041 20488
rect 24075 20485 24087 20519
rect 24029 20479 24087 20485
rect 24121 20519 24179 20525
rect 24121 20485 24133 20519
rect 24167 20485 24179 20519
rect 24121 20479 24179 20485
rect 24394 20476 24400 20528
rect 24452 20516 24458 20528
rect 25222 20516 25228 20528
rect 24452 20488 25228 20516
rect 24452 20476 24458 20488
rect 25222 20476 25228 20488
rect 25280 20476 25286 20528
rect 27338 20516 27344 20528
rect 27299 20488 27344 20516
rect 27338 20476 27344 20488
rect 27396 20476 27402 20528
rect 28905 20519 28963 20525
rect 28905 20485 28917 20519
rect 28951 20516 28963 20519
rect 30374 20516 30380 20528
rect 28951 20488 30380 20516
rect 28951 20485 28963 20488
rect 28905 20479 28963 20485
rect 30374 20476 30380 20488
rect 30432 20476 30438 20528
rect 30745 20519 30803 20525
rect 30745 20485 30757 20519
rect 30791 20516 30803 20519
rect 32398 20516 32404 20528
rect 30791 20488 31984 20516
rect 32359 20488 32404 20516
rect 30791 20485 30803 20488
rect 30745 20479 30803 20485
rect 12207 20420 12434 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12952 20420 13001 20448
rect 12952 20408 12958 20420
rect 12989 20417 13001 20420
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 13633 20451 13691 20457
rect 13633 20448 13645 20451
rect 13412 20420 13645 20448
rect 13412 20408 13418 20420
rect 13633 20417 13645 20420
rect 13679 20417 13691 20451
rect 16114 20448 16120 20460
rect 16075 20420 16120 20448
rect 13633 20411 13691 20417
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 19628 20420 20269 20448
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 14550 20380 14556 20392
rect 14415 20352 14556 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 14550 20340 14556 20352
rect 14608 20380 14614 20392
rect 14826 20380 14832 20392
rect 14608 20352 14832 20380
rect 14608 20340 14614 20352
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 15194 20380 15200 20392
rect 15155 20352 15200 20380
rect 15194 20340 15200 20352
rect 15252 20340 15258 20392
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20349 17003 20383
rect 17862 20380 17868 20392
rect 17823 20352 17868 20380
rect 16945 20343 17003 20349
rect 6638 20272 6644 20324
rect 6696 20312 6702 20324
rect 13081 20315 13139 20321
rect 13081 20312 13093 20315
rect 6696 20284 13093 20312
rect 6696 20272 6702 20284
rect 13081 20281 13093 20284
rect 13127 20281 13139 20315
rect 16960 20312 16988 20343
rect 17862 20340 17868 20352
rect 17920 20340 17926 20392
rect 18230 20340 18236 20392
rect 18288 20380 18294 20392
rect 18785 20383 18843 20389
rect 18785 20380 18797 20383
rect 18288 20352 18797 20380
rect 18288 20340 18294 20352
rect 18785 20349 18797 20352
rect 18831 20349 18843 20383
rect 18785 20343 18843 20349
rect 13081 20275 13139 20281
rect 14384 20284 16988 20312
rect 1762 20244 1768 20256
rect 1723 20216 1768 20244
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 11698 20204 11704 20256
rect 11756 20244 11762 20256
rect 12253 20247 12311 20253
rect 12253 20244 12265 20247
rect 11756 20216 12265 20244
rect 11756 20204 11762 20216
rect 12253 20213 12265 20216
rect 12299 20213 12311 20247
rect 12253 20207 12311 20213
rect 12342 20204 12348 20256
rect 12400 20244 12406 20256
rect 14384 20244 14412 20284
rect 12400 20216 14412 20244
rect 12400 20204 12406 20216
rect 14458 20204 14464 20256
rect 14516 20244 14522 20256
rect 16390 20244 16396 20256
rect 14516 20216 16396 20244
rect 14516 20204 14522 20216
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 17770 20244 17776 20256
rect 16816 20216 17776 20244
rect 16816 20204 16822 20216
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 19628 20244 19656 20420
rect 20257 20417 20269 20420
rect 20303 20417 20315 20451
rect 20898 20448 20904 20460
rect 20859 20420 20904 20448
rect 20257 20411 20315 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20380 19855 20383
rect 20070 20380 20076 20392
rect 19843 20352 20076 20380
rect 19843 20349 19855 20352
rect 19797 20343 19855 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20380 22155 20383
rect 22370 20380 22376 20392
rect 22143 20352 22376 20380
rect 22143 20349 22155 20352
rect 22097 20343 22155 20349
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 23109 20383 23167 20389
rect 23109 20380 23121 20383
rect 22612 20352 23121 20380
rect 22612 20340 22618 20352
rect 23109 20349 23121 20352
rect 23155 20380 23167 20383
rect 24210 20380 24216 20392
rect 23155 20352 24216 20380
rect 23155 20349 23167 20352
rect 23109 20343 23167 20349
rect 24210 20340 24216 20352
rect 24268 20340 24274 20392
rect 24302 20340 24308 20392
rect 24360 20380 24366 20392
rect 24360 20352 24405 20380
rect 24360 20340 24366 20352
rect 20088 20312 20116 20340
rect 22278 20312 22284 20324
rect 20088 20284 22284 20312
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 22830 20272 22836 20324
rect 22888 20312 22894 20324
rect 25516 20312 25544 20411
rect 25774 20408 25780 20460
rect 25832 20448 25838 20460
rect 26145 20451 26203 20457
rect 26145 20448 26157 20451
rect 25832 20420 26157 20448
rect 25832 20408 25838 20420
rect 26145 20417 26157 20420
rect 26191 20448 26203 20451
rect 26878 20448 26884 20460
rect 26191 20420 26884 20448
rect 26191 20417 26203 20420
rect 26145 20411 26203 20417
rect 26878 20408 26884 20420
rect 26936 20448 26942 20460
rect 27062 20448 27068 20460
rect 26936 20420 27068 20448
rect 26936 20408 26942 20420
rect 27062 20408 27068 20420
rect 27120 20408 27126 20460
rect 27249 20383 27307 20389
rect 27249 20349 27261 20383
rect 27295 20349 27307 20383
rect 27614 20380 27620 20392
rect 27575 20352 27620 20380
rect 27249 20343 27307 20349
rect 22888 20284 25544 20312
rect 22888 20272 22894 20284
rect 18288 20216 19656 20244
rect 20993 20247 21051 20253
rect 18288 20204 18294 20216
rect 20993 20213 21005 20247
rect 21039 20244 21051 20247
rect 21450 20244 21456 20256
rect 21039 20216 21456 20244
rect 21039 20213 21051 20216
rect 20993 20207 21051 20213
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 23014 20204 23020 20256
rect 23072 20244 23078 20256
rect 25593 20247 25651 20253
rect 25593 20244 25605 20247
rect 23072 20216 25605 20244
rect 23072 20204 23078 20216
rect 25593 20213 25605 20216
rect 25639 20213 25651 20247
rect 26234 20244 26240 20256
rect 26195 20216 26240 20244
rect 25593 20207 25651 20213
rect 26234 20204 26240 20216
rect 26292 20204 26298 20256
rect 27264 20244 27292 20343
rect 27614 20340 27620 20352
rect 27672 20380 27678 20392
rect 27890 20380 27896 20392
rect 27672 20352 27896 20380
rect 27672 20340 27678 20352
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 28810 20380 28816 20392
rect 28771 20352 28816 20380
rect 28810 20340 28816 20352
rect 28868 20340 28874 20392
rect 28994 20340 29000 20392
rect 29052 20380 29058 20392
rect 29089 20383 29147 20389
rect 29089 20380 29101 20383
rect 29052 20352 29101 20380
rect 29052 20340 29058 20352
rect 29089 20349 29101 20352
rect 29135 20349 29147 20383
rect 29089 20343 29147 20349
rect 29454 20340 29460 20392
rect 29512 20380 29518 20392
rect 30374 20380 30380 20392
rect 29512 20352 30380 20380
rect 29512 20340 29518 20352
rect 30374 20340 30380 20352
rect 30432 20340 30438 20392
rect 30653 20383 30711 20389
rect 30653 20349 30665 20383
rect 30699 20349 30711 20383
rect 30653 20343 30711 20349
rect 31297 20383 31355 20389
rect 31297 20349 31309 20383
rect 31343 20349 31355 20383
rect 31956 20380 31984 20488
rect 32398 20476 32404 20488
rect 32456 20476 32462 20528
rect 32493 20519 32551 20525
rect 32493 20485 32505 20519
rect 32539 20516 32551 20519
rect 33410 20516 33416 20528
rect 32539 20488 33416 20516
rect 32539 20485 32551 20488
rect 32493 20479 32551 20485
rect 33410 20476 33416 20488
rect 33468 20476 33474 20528
rect 33597 20519 33655 20525
rect 33597 20485 33609 20519
rect 33643 20516 33655 20519
rect 34054 20516 34060 20528
rect 33643 20488 34060 20516
rect 33643 20485 33655 20488
rect 33597 20479 33655 20485
rect 34054 20476 34060 20488
rect 34112 20476 34118 20528
rect 33505 20451 33563 20457
rect 33505 20417 33517 20451
rect 33551 20448 33563 20451
rect 33686 20448 33692 20460
rect 33551 20420 33692 20448
rect 33551 20417 33563 20420
rect 33505 20411 33563 20417
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 34146 20448 34152 20460
rect 34107 20420 34152 20448
rect 34146 20408 34152 20420
rect 34204 20408 34210 20460
rect 34808 20457 34836 20556
rect 34793 20451 34851 20457
rect 34793 20417 34805 20451
rect 34839 20417 34851 20451
rect 34793 20411 34851 20417
rect 34241 20383 34299 20389
rect 34241 20380 34253 20383
rect 31956 20368 32168 20380
rect 32324 20368 34253 20380
rect 31956 20352 34253 20368
rect 31297 20343 31355 20349
rect 27430 20272 27436 20324
rect 27488 20312 27494 20324
rect 30558 20312 30564 20324
rect 27488 20284 30564 20312
rect 27488 20272 27494 20284
rect 30558 20272 30564 20284
rect 30616 20272 30622 20324
rect 30668 20312 30696 20343
rect 31018 20312 31024 20324
rect 30668 20284 31024 20312
rect 31018 20272 31024 20284
rect 31076 20272 31082 20324
rect 29914 20244 29920 20256
rect 27264 20216 29920 20244
rect 29914 20204 29920 20216
rect 29972 20204 29978 20256
rect 30190 20204 30196 20256
rect 30248 20244 30254 20256
rect 31312 20244 31340 20343
rect 32140 20340 32352 20352
rect 34241 20349 34253 20352
rect 34287 20349 34299 20383
rect 34241 20343 34299 20349
rect 32950 20312 32956 20324
rect 32911 20284 32956 20312
rect 32950 20272 32956 20284
rect 33008 20272 33014 20324
rect 30248 20216 31340 20244
rect 30248 20204 30254 20216
rect 32122 20204 32128 20256
rect 32180 20244 32186 20256
rect 34885 20247 34943 20253
rect 34885 20244 34897 20247
rect 32180 20216 34897 20244
rect 32180 20204 32186 20216
rect 34885 20213 34897 20216
rect 34931 20213 34943 20247
rect 34885 20207 34943 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 15562 20040 15568 20052
rect 7984 20012 15568 20040
rect 7984 20000 7990 20012
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 15988 20012 16129 20040
rect 15988 20000 15994 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 16117 20003 16175 20009
rect 17405 20043 17463 20049
rect 17405 20009 17417 20043
rect 17451 20040 17463 20043
rect 17494 20040 17500 20052
rect 17451 20012 17500 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 17770 20000 17776 20052
rect 17828 20040 17834 20052
rect 23658 20040 23664 20052
rect 17828 20012 23664 20040
rect 17828 20000 17834 20012
rect 23658 20000 23664 20012
rect 23716 20040 23722 20052
rect 23716 20012 24992 20040
rect 23716 20000 23722 20012
rect 6178 19932 6184 19984
rect 6236 19972 6242 19984
rect 13170 19972 13176 19984
rect 6236 19944 13176 19972
rect 6236 19932 6242 19944
rect 13170 19932 13176 19944
rect 13228 19932 13234 19984
rect 15838 19932 15844 19984
rect 15896 19972 15902 19984
rect 20073 19975 20131 19981
rect 20073 19972 20085 19975
rect 15896 19944 20085 19972
rect 15896 19932 15902 19944
rect 20073 19941 20085 19944
rect 20119 19972 20131 19975
rect 20162 19972 20168 19984
rect 20119 19944 20168 19972
rect 20119 19941 20131 19944
rect 20073 19935 20131 19941
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 20622 19932 20628 19984
rect 20680 19932 20686 19984
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 24026 19972 24032 19984
rect 22152 19944 24032 19972
rect 22152 19932 22158 19944
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19904 1915 19907
rect 11606 19904 11612 19916
rect 1903 19876 11612 19904
rect 1903 19873 1915 19876
rect 1857 19867 1915 19873
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 12253 19907 12311 19913
rect 12253 19873 12265 19907
rect 12299 19904 12311 19907
rect 12342 19904 12348 19916
rect 12299 19876 12348 19904
rect 12299 19873 12311 19876
rect 12253 19867 12311 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20640 19904 20668 19932
rect 19567 19876 20668 19904
rect 21361 19907 21419 19913
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 21361 19873 21373 19907
rect 21407 19904 21419 19907
rect 21910 19904 21916 19916
rect 21407 19876 21916 19904
rect 21407 19873 21419 19876
rect 21361 19867 21419 19873
rect 21910 19864 21916 19876
rect 21968 19904 21974 19916
rect 23216 19913 23244 19944
rect 24026 19932 24032 19944
rect 24084 19932 24090 19984
rect 22925 19907 22983 19913
rect 22925 19904 22937 19907
rect 21968 19876 22937 19904
rect 21968 19864 21974 19876
rect 22925 19873 22937 19876
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 23201 19907 23259 19913
rect 23201 19873 23213 19907
rect 23247 19873 23259 19907
rect 23201 19867 23259 19873
rect 23750 19864 23756 19916
rect 23808 19904 23814 19916
rect 24964 19913 24992 20012
rect 25130 20000 25136 20052
rect 25188 20040 25194 20052
rect 25866 20040 25872 20052
rect 25188 20012 25872 20040
rect 25188 20000 25194 20012
rect 25866 20000 25872 20012
rect 25924 20000 25930 20052
rect 26142 20000 26148 20052
rect 26200 20040 26206 20052
rect 28350 20040 28356 20052
rect 26200 20012 28356 20040
rect 26200 20000 26206 20012
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 30190 20040 30196 20052
rect 29656 20012 30196 20040
rect 25314 19932 25320 19984
rect 25372 19972 25378 19984
rect 28258 19972 28264 19984
rect 25372 19944 28264 19972
rect 25372 19932 25378 19944
rect 28258 19932 28264 19944
rect 28316 19932 28322 19984
rect 29546 19972 29552 19984
rect 28966 19944 29552 19972
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 23808 19876 24685 19904
rect 23808 19864 23814 19876
rect 24673 19873 24685 19876
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 24949 19907 25007 19913
rect 24949 19873 24961 19907
rect 24995 19873 25007 19907
rect 24949 19867 25007 19873
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 26973 19907 27031 19913
rect 26973 19904 26985 19907
rect 25096 19876 26985 19904
rect 25096 19864 25102 19876
rect 26973 19873 26985 19876
rect 27019 19873 27031 19907
rect 27430 19904 27436 19916
rect 27391 19876 27436 19904
rect 26973 19867 27031 19873
rect 27430 19864 27436 19876
rect 27488 19864 27494 19916
rect 28718 19904 28724 19916
rect 28679 19876 28724 19904
rect 28718 19864 28724 19876
rect 28776 19864 28782 19916
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13630 19836 13636 19848
rect 12943 19808 13636 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 15436 19808 15481 19836
rect 15436 19796 15442 19808
rect 15562 19796 15568 19848
rect 15620 19836 15626 19848
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15620 19808 16037 19836
rect 15620 19796 15626 19808
rect 16025 19805 16037 19808
rect 16071 19805 16083 19839
rect 16666 19836 16672 19848
rect 16627 19808 16672 19836
rect 16025 19799 16083 19805
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 17494 19836 17500 19848
rect 17359 19808 17500 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 20622 19836 20628 19848
rect 20583 19808 20628 19836
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 26142 19836 26148 19848
rect 26103 19808 26148 19836
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 27982 19796 27988 19848
rect 28040 19836 28046 19848
rect 28077 19839 28135 19845
rect 28077 19836 28089 19839
rect 28040 19808 28089 19836
rect 28040 19796 28046 19808
rect 28077 19805 28089 19808
rect 28123 19836 28135 19839
rect 28966 19836 28994 19944
rect 29546 19932 29552 19944
rect 29604 19932 29610 19984
rect 28123 19808 28994 19836
rect 28123 19805 28135 19808
rect 28077 19799 28135 19805
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 11609 19771 11667 19777
rect 11609 19768 11621 19771
rect 11020 19740 11621 19768
rect 11020 19728 11026 19740
rect 11609 19737 11621 19740
rect 11655 19737 11667 19771
rect 11609 19731 11667 19737
rect 11698 19728 11704 19780
rect 11756 19768 11762 19780
rect 15102 19768 15108 19780
rect 11756 19740 11801 19768
rect 12406 19740 15108 19768
rect 11756 19728 11762 19740
rect 8570 19660 8576 19712
rect 8628 19700 8634 19712
rect 12406 19700 12434 19740
rect 15102 19728 15108 19740
rect 15160 19728 15166 19780
rect 15470 19768 15476 19780
rect 15431 19740 15476 19768
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 18049 19771 18107 19777
rect 18049 19768 18061 19771
rect 15580 19740 18061 19768
rect 12986 19700 12992 19712
rect 8628 19672 12434 19700
rect 12947 19672 12992 19700
rect 8628 19660 8634 19672
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 14734 19700 14740 19712
rect 14056 19672 14740 19700
rect 14056 19660 14062 19672
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15010 19660 15016 19712
rect 15068 19700 15074 19712
rect 15580 19700 15608 19740
rect 18049 19737 18061 19740
rect 18095 19737 18107 19771
rect 18049 19731 18107 19737
rect 18138 19728 18144 19780
rect 18196 19768 18202 19780
rect 18693 19771 18751 19777
rect 18196 19740 18241 19768
rect 18196 19728 18202 19740
rect 18693 19737 18705 19771
rect 18739 19768 18751 19771
rect 18874 19768 18880 19780
rect 18739 19740 18880 19768
rect 18739 19737 18751 19740
rect 18693 19731 18751 19737
rect 18874 19728 18880 19740
rect 18932 19728 18938 19780
rect 19613 19771 19671 19777
rect 19613 19737 19625 19771
rect 19659 19737 19671 19771
rect 21450 19768 21456 19780
rect 21411 19740 21456 19768
rect 19613 19731 19671 19737
rect 15068 19672 15608 19700
rect 16761 19703 16819 19709
rect 15068 19660 15074 19672
rect 16761 19669 16773 19703
rect 16807 19700 16819 19703
rect 19334 19700 19340 19712
rect 16807 19672 19340 19700
rect 16807 19669 16819 19672
rect 16761 19663 16819 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 19628 19700 19656 19731
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 22370 19768 22376 19780
rect 22331 19740 22376 19768
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 23014 19728 23020 19780
rect 23072 19768 23078 19780
rect 23072 19740 23117 19768
rect 23072 19728 23078 19740
rect 24210 19728 24216 19780
rect 24268 19768 24274 19780
rect 24742 19771 24800 19777
rect 24742 19768 24754 19771
rect 24268 19740 24754 19768
rect 24268 19728 24274 19740
rect 24742 19737 24754 19740
rect 24788 19737 24800 19771
rect 24742 19731 24800 19737
rect 27065 19771 27123 19777
rect 27065 19737 27077 19771
rect 27111 19768 27123 19771
rect 27111 19740 27292 19768
rect 27111 19737 27123 19740
rect 27065 19731 27123 19737
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 19628 19672 20729 19700
rect 20717 19669 20729 19672
rect 20763 19669 20775 19703
rect 20717 19663 20775 19669
rect 20898 19660 20904 19712
rect 20956 19700 20962 19712
rect 22554 19700 22560 19712
rect 20956 19672 22560 19700
rect 20956 19660 20962 19672
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 23658 19660 23664 19712
rect 23716 19700 23722 19712
rect 26237 19703 26295 19709
rect 26237 19700 26249 19703
rect 23716 19672 26249 19700
rect 23716 19660 23722 19672
rect 26237 19669 26249 19672
rect 26283 19669 26295 19703
rect 27264 19700 27292 19740
rect 27890 19728 27896 19780
rect 27948 19768 27954 19780
rect 29362 19768 29368 19780
rect 27948 19740 29368 19768
rect 27948 19728 27954 19740
rect 29362 19728 29368 19740
rect 29420 19768 29426 19780
rect 29656 19768 29684 20012
rect 30190 20000 30196 20012
rect 30248 20000 30254 20052
rect 30374 20000 30380 20052
rect 30432 20040 30438 20052
rect 30432 20012 31156 20040
rect 30432 20000 30438 20012
rect 31018 19972 31024 19984
rect 29840 19944 31024 19972
rect 29840 19913 29868 19944
rect 31018 19932 31024 19944
rect 31076 19932 31082 19984
rect 31128 19972 31156 20012
rect 31938 20000 31944 20052
rect 31996 20040 32002 20052
rect 33045 20043 33103 20049
rect 33045 20040 33057 20043
rect 31996 20012 33057 20040
rect 31996 20000 32002 20012
rect 33045 20009 33057 20012
rect 33091 20009 33103 20043
rect 33045 20003 33103 20009
rect 33410 20000 33416 20052
rect 33468 20040 33474 20052
rect 34977 20043 35035 20049
rect 34977 20040 34989 20043
rect 33468 20012 34989 20040
rect 33468 20000 33474 20012
rect 34977 20009 34989 20012
rect 35023 20009 35035 20043
rect 34977 20003 35035 20009
rect 38289 19975 38347 19981
rect 38289 19972 38301 19975
rect 31128 19944 38301 19972
rect 38289 19941 38301 19944
rect 38335 19941 38347 19975
rect 38289 19935 38347 19941
rect 29825 19907 29883 19913
rect 29825 19873 29837 19907
rect 29871 19873 29883 19907
rect 29825 19867 29883 19873
rect 29914 19864 29920 19916
rect 29972 19904 29978 19916
rect 33689 19907 33747 19913
rect 33689 19904 33701 19907
rect 29972 19876 33701 19904
rect 29972 19864 29978 19876
rect 33689 19873 33701 19876
rect 33735 19873 33747 19907
rect 33689 19867 33747 19873
rect 34606 19864 34612 19916
rect 34664 19904 34670 19916
rect 38746 19904 38752 19916
rect 34664 19876 38752 19904
rect 34664 19864 34670 19876
rect 38746 19864 38752 19876
rect 38804 19864 38810 19916
rect 30469 19839 30527 19845
rect 30469 19805 30481 19839
rect 30515 19836 30527 19839
rect 30558 19836 30564 19848
rect 30515 19808 30564 19836
rect 30515 19805 30527 19808
rect 30469 19799 30527 19805
rect 30558 19796 30564 19808
rect 30616 19796 30622 19848
rect 31849 19839 31907 19845
rect 31849 19805 31861 19839
rect 31895 19836 31907 19839
rect 31938 19836 31944 19848
rect 31895 19808 31944 19836
rect 31895 19805 31907 19808
rect 31849 19799 31907 19805
rect 31938 19796 31944 19808
rect 31996 19836 32002 19848
rect 32214 19836 32220 19848
rect 31996 19808 32220 19836
rect 31996 19796 32002 19808
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32306 19796 32312 19848
rect 32364 19836 32370 19848
rect 32950 19836 32956 19848
rect 32364 19808 32409 19836
rect 32911 19808 32956 19836
rect 32364 19796 32370 19808
rect 32950 19796 32956 19808
rect 33008 19796 33014 19848
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19836 33655 19839
rect 34146 19836 34152 19848
rect 33643 19808 34152 19836
rect 33643 19805 33655 19808
rect 33597 19799 33655 19805
rect 34146 19796 34152 19808
rect 34204 19796 34210 19848
rect 34790 19796 34796 19848
rect 34848 19836 34854 19848
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 34848 19808 34897 19836
rect 34848 19796 34854 19808
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 29420 19740 29684 19768
rect 29917 19771 29975 19777
rect 29420 19728 29426 19740
rect 29917 19737 29929 19771
rect 29963 19768 29975 19771
rect 31202 19768 31208 19780
rect 29963 19740 30144 19768
rect 31163 19740 31208 19768
rect 29963 19737 29975 19740
rect 29917 19731 29975 19737
rect 28169 19703 28227 19709
rect 28169 19700 28181 19703
rect 27264 19672 28181 19700
rect 26237 19663 26295 19669
rect 28169 19669 28181 19672
rect 28215 19669 28227 19703
rect 28169 19663 28227 19669
rect 28810 19660 28816 19712
rect 28868 19700 28874 19712
rect 29730 19700 29736 19712
rect 28868 19672 29736 19700
rect 28868 19660 28874 19672
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 30116 19700 30144 19740
rect 31202 19728 31208 19740
rect 31260 19728 31266 19780
rect 31294 19728 31300 19780
rect 31352 19768 31358 19780
rect 34422 19768 34428 19780
rect 31352 19740 31397 19768
rect 31496 19740 34428 19768
rect 31352 19728 31358 19740
rect 30190 19700 30196 19712
rect 30116 19672 30196 19700
rect 30190 19660 30196 19672
rect 30248 19660 30254 19712
rect 31386 19660 31392 19712
rect 31444 19700 31450 19712
rect 31496 19700 31524 19740
rect 34422 19728 34428 19740
rect 34480 19728 34486 19780
rect 38102 19768 38108 19780
rect 38063 19740 38108 19768
rect 38102 19728 38108 19740
rect 38160 19728 38166 19780
rect 31444 19672 31524 19700
rect 31444 19660 31450 19672
rect 32398 19660 32404 19712
rect 32456 19700 32462 19712
rect 32456 19672 32501 19700
rect 32456 19660 32462 19672
rect 33318 19660 33324 19712
rect 33376 19700 33382 19712
rect 34698 19700 34704 19712
rect 33376 19672 34704 19700
rect 33376 19660 33382 19672
rect 34698 19660 34704 19672
rect 34756 19660 34762 19712
rect 35342 19660 35348 19712
rect 35400 19700 35406 19712
rect 37642 19700 37648 19712
rect 35400 19672 37648 19700
rect 35400 19660 35406 19672
rect 37642 19660 37648 19672
rect 37700 19660 37706 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 7558 19496 7564 19508
rect 7519 19468 7564 19496
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 8389 19499 8447 19505
rect 8389 19465 8401 19499
rect 8435 19496 8447 19499
rect 8478 19496 8484 19508
rect 8435 19468 8484 19496
rect 8435 19465 8447 19468
rect 8389 19459 8447 19465
rect 8478 19456 8484 19468
rect 8536 19456 8542 19508
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 10962 19496 10968 19508
rect 9171 19468 10968 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 13170 19496 13176 19508
rect 13131 19468 13176 19496
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13817 19499 13875 19505
rect 13817 19496 13829 19499
rect 13320 19468 13829 19496
rect 13320 19456 13326 19468
rect 13817 19465 13829 19468
rect 13863 19465 13875 19499
rect 13817 19459 13875 19465
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 14461 19499 14519 19505
rect 14461 19496 14473 19499
rect 14332 19468 14473 19496
rect 14332 19456 14338 19468
rect 14461 19465 14473 19468
rect 14507 19465 14519 19499
rect 14461 19459 14519 19465
rect 15120 19468 27476 19496
rect 9766 19428 9772 19440
rect 7484 19400 9772 19428
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 1762 19360 1768 19372
rect 1627 19332 1768 19360
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 7484 19369 7512 19400
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 10134 19428 10140 19440
rect 10095 19400 10140 19428
rect 10134 19388 10140 19400
rect 10192 19388 10198 19440
rect 10229 19431 10287 19437
rect 10229 19397 10241 19431
rect 10275 19428 10287 19431
rect 11790 19428 11796 19440
rect 10275 19400 11796 19428
rect 10275 19397 10287 19400
rect 10229 19391 10287 19397
rect 11790 19388 11796 19400
rect 11848 19388 11854 19440
rect 11974 19388 11980 19440
rect 12032 19428 12038 19440
rect 15010 19428 15016 19440
rect 12032 19400 15016 19428
rect 12032 19388 12038 19400
rect 15010 19388 15016 19400
rect 15068 19388 15074 19440
rect 7469 19363 7527 19369
rect 5500 19332 7420 19360
rect 5500 19320 5506 19332
rect 7392 19292 7420 19332
rect 7469 19329 7481 19363
rect 7515 19329 7527 19363
rect 8570 19360 8576 19372
rect 7469 19323 7527 19329
rect 7576 19332 8432 19360
rect 8531 19332 8576 19360
rect 7576 19292 7604 19332
rect 7392 19264 7604 19292
rect 8404 19292 8432 19332
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8680 19332 9045 19360
rect 8680 19292 8708 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12952 19332 13093 19360
rect 12952 19320 12958 19332
rect 13081 19329 13093 19332
rect 13127 19360 13139 19363
rect 13725 19363 13783 19369
rect 13725 19360 13737 19363
rect 13127 19332 13737 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13725 19329 13737 19332
rect 13771 19360 13783 19363
rect 14369 19363 14427 19369
rect 13771 19332 14320 19360
rect 13771 19329 13783 19332
rect 13725 19323 13783 19329
rect 8404 19264 8708 19292
rect 11149 19295 11207 19301
rect 11149 19261 11161 19295
rect 11195 19292 11207 19295
rect 12526 19292 12532 19304
rect 11195 19264 12532 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 14292 19292 14320 19332
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 14734 19360 14740 19372
rect 14415 19332 14740 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15120 19369 15148 19468
rect 17402 19428 17408 19440
rect 17363 19400 17408 19428
rect 17402 19388 17408 19400
rect 17460 19388 17466 19440
rect 18598 19428 18604 19440
rect 18559 19400 18604 19428
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 19334 19388 19340 19440
rect 19392 19428 19398 19440
rect 20165 19431 20223 19437
rect 20165 19428 20177 19431
rect 19392 19400 20177 19428
rect 19392 19388 19398 19400
rect 20165 19397 20177 19400
rect 20211 19397 20223 19431
rect 20165 19391 20223 19397
rect 20346 19388 20352 19440
rect 20404 19428 20410 19440
rect 20898 19428 20904 19440
rect 20404 19400 20904 19428
rect 20404 19388 20410 19400
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 21082 19428 21088 19440
rect 21043 19400 21088 19428
rect 21082 19388 21088 19400
rect 21140 19388 21146 19440
rect 22094 19388 22100 19440
rect 22152 19428 22158 19440
rect 22925 19431 22983 19437
rect 22152 19400 22197 19428
rect 22152 19388 22158 19400
rect 22925 19397 22937 19431
rect 22971 19428 22983 19431
rect 23014 19428 23020 19440
rect 22971 19400 23020 19428
rect 22971 19397 22983 19400
rect 22925 19391 22983 19397
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 23658 19437 23664 19440
rect 23654 19391 23664 19437
rect 23716 19428 23722 19440
rect 23716 19400 23754 19428
rect 23658 19388 23664 19391
rect 23716 19388 23722 19400
rect 23934 19388 23940 19440
rect 23992 19428 23998 19440
rect 25133 19431 25191 19437
rect 25133 19428 25145 19431
rect 23992 19400 25145 19428
rect 23992 19388 23998 19400
rect 25133 19397 25145 19400
rect 25179 19397 25191 19431
rect 25133 19391 25191 19397
rect 25225 19431 25283 19437
rect 25225 19397 25237 19431
rect 25271 19428 25283 19431
rect 26234 19428 26240 19440
rect 25271 19400 26240 19428
rect 25271 19397 25283 19400
rect 25225 19391 25283 19397
rect 26234 19388 26240 19400
rect 26292 19388 26298 19440
rect 27338 19428 27344 19440
rect 27299 19400 27344 19428
rect 27338 19388 27344 19400
rect 27396 19388 27402 19440
rect 27448 19428 27476 19468
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28813 19499 28871 19505
rect 28813 19496 28825 19499
rect 28132 19468 28825 19496
rect 28132 19456 28138 19468
rect 28813 19465 28825 19468
rect 28859 19465 28871 19499
rect 31570 19496 31576 19508
rect 28813 19459 28871 19465
rect 28966 19468 31576 19496
rect 28966 19428 28994 19468
rect 31570 19456 31576 19468
rect 31628 19456 31634 19508
rect 33318 19496 33324 19508
rect 31726 19468 33324 19496
rect 29730 19428 29736 19440
rect 27448 19400 28994 19428
rect 29691 19400 29736 19428
rect 29730 19388 29736 19400
rect 29788 19388 29794 19440
rect 30006 19388 30012 19440
rect 30064 19428 30070 19440
rect 31205 19431 31263 19437
rect 30064 19400 30512 19428
rect 30064 19388 30070 19400
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15194 19320 15200 19372
rect 15252 19360 15258 19372
rect 15252 19332 15297 19360
rect 15252 19320 15258 19332
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 16298 19360 16304 19372
rect 15436 19332 16304 19360
rect 15436 19320 15442 19332
rect 16298 19320 16304 19332
rect 16356 19320 16362 19372
rect 16390 19320 16396 19372
rect 16448 19360 16454 19372
rect 16448 19332 17172 19360
rect 16448 19320 16454 19332
rect 15396 19292 15424 19320
rect 14292 19264 15424 19292
rect 17144 19292 17172 19332
rect 21818 19320 21824 19372
rect 21876 19320 21882 19372
rect 22002 19360 22008 19372
rect 21963 19332 22008 19360
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 22830 19360 22836 19372
rect 22112 19332 22836 19360
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 17144 19264 17325 19292
rect 17313 19261 17325 19264
rect 17359 19261 17371 19295
rect 18506 19292 18512 19304
rect 18467 19264 18512 19292
rect 17313 19255 17371 19261
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19261 19579 19295
rect 20070 19292 20076 19304
rect 20031 19264 20076 19292
rect 19521 19255 19579 19261
rect 6546 19184 6552 19236
rect 6604 19224 6610 19236
rect 17865 19227 17923 19233
rect 6604 19196 17264 19224
rect 6604 19184 6610 19196
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 17236 19156 17264 19196
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 18874 19224 18880 19236
rect 17911 19196 18880 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 18874 19184 18880 19196
rect 18932 19184 18938 19236
rect 19536 19224 19564 19255
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 21836 19292 21864 19320
rect 22112 19292 22140 19332
rect 22830 19320 22836 19332
rect 22888 19320 22894 19372
rect 23382 19320 23388 19372
rect 23440 19320 23446 19372
rect 27062 19360 27068 19372
rect 26160 19332 27068 19360
rect 21836 19264 22140 19292
rect 23400 19292 23428 19320
rect 23569 19295 23627 19301
rect 23569 19292 23581 19295
rect 23400 19264 23581 19292
rect 23569 19261 23581 19264
rect 23615 19261 23627 19295
rect 24118 19292 24124 19304
rect 24079 19264 24124 19292
rect 23569 19255 23627 19261
rect 24118 19252 24124 19264
rect 24176 19252 24182 19304
rect 26160 19301 26188 19332
rect 27062 19320 27068 19332
rect 27120 19320 27126 19372
rect 28442 19360 28448 19372
rect 28092 19332 28448 19360
rect 26145 19295 26203 19301
rect 26145 19261 26157 19295
rect 26191 19261 26203 19295
rect 27246 19292 27252 19304
rect 27207 19264 27252 19292
rect 26145 19255 26203 19261
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 27338 19252 27344 19304
rect 27396 19292 27402 19304
rect 28092 19292 28120 19332
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28534 19320 28540 19372
rect 28592 19360 28598 19372
rect 28721 19363 28779 19369
rect 28721 19360 28733 19363
rect 28592 19332 28733 19360
rect 28592 19320 28598 19332
rect 28721 19329 28733 19332
rect 28767 19329 28779 19363
rect 28721 19323 28779 19329
rect 28902 19320 28908 19372
rect 28960 19360 28966 19372
rect 29454 19360 29460 19372
rect 28960 19332 29460 19360
rect 28960 19320 28966 19332
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 30484 19360 30512 19400
rect 31205 19397 31217 19431
rect 31251 19428 31263 19431
rect 31726 19428 31754 19468
rect 33318 19456 33324 19468
rect 33376 19456 33382 19508
rect 35161 19499 35219 19505
rect 35161 19496 35173 19499
rect 33428 19468 35173 19496
rect 32398 19428 32404 19440
rect 31251 19400 31754 19428
rect 32048 19400 32404 19428
rect 31251 19397 31263 19400
rect 31205 19391 31263 19397
rect 32048 19360 32076 19400
rect 32398 19388 32404 19400
rect 32456 19388 32462 19440
rect 33428 19437 33456 19468
rect 35161 19465 35173 19468
rect 35207 19465 35219 19499
rect 36262 19496 36268 19508
rect 36223 19468 36268 19496
rect 35161 19459 35219 19465
rect 36262 19456 36268 19468
rect 36320 19456 36326 19508
rect 38010 19456 38016 19508
rect 38068 19496 38074 19508
rect 38105 19499 38163 19505
rect 38105 19496 38117 19499
rect 38068 19468 38117 19496
rect 38068 19456 38074 19468
rect 38105 19465 38117 19468
rect 38151 19465 38163 19499
rect 38105 19459 38163 19465
rect 33413 19431 33471 19437
rect 33413 19397 33425 19431
rect 33459 19397 33471 19431
rect 33413 19391 33471 19397
rect 33502 19388 33508 19440
rect 33560 19428 33566 19440
rect 33560 19400 33605 19428
rect 33560 19388 33566 19400
rect 34054 19388 34060 19440
rect 34112 19428 34118 19440
rect 34609 19431 34667 19437
rect 34609 19428 34621 19431
rect 34112 19400 34621 19428
rect 34112 19388 34118 19400
rect 34609 19397 34621 19400
rect 34655 19397 34667 19431
rect 34609 19391 34667 19397
rect 32306 19360 32312 19372
rect 30484 19332 32076 19360
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 34514 19360 34520 19372
rect 34475 19332 34520 19360
rect 34514 19320 34520 19332
rect 34572 19320 34578 19372
rect 36449 19363 36507 19369
rect 36449 19329 36461 19363
rect 36495 19329 36507 19363
rect 38286 19360 38292 19372
rect 38247 19332 38292 19360
rect 36449 19323 36507 19329
rect 27396 19264 28120 19292
rect 28261 19295 28319 19301
rect 27396 19252 27402 19264
rect 28261 19261 28273 19295
rect 28307 19292 28319 19295
rect 28350 19292 28356 19304
rect 28307 19264 28356 19292
rect 28307 19261 28319 19264
rect 28261 19255 28319 19261
rect 28350 19252 28356 19264
rect 28408 19252 28414 19304
rect 29638 19292 29644 19304
rect 28460 19264 28672 19292
rect 29599 19264 29644 19292
rect 20714 19224 20720 19236
rect 19536 19196 20720 19224
rect 20714 19184 20720 19196
rect 20772 19184 20778 19236
rect 28460 19224 28488 19264
rect 22066 19196 28488 19224
rect 28644 19224 28672 19264
rect 29638 19252 29644 19264
rect 29696 19252 29702 19304
rect 30006 19292 30012 19304
rect 29967 19264 30012 19292
rect 30006 19252 30012 19264
rect 30064 19292 30070 19304
rect 30926 19292 30932 19304
rect 30064 19264 30932 19292
rect 30064 19252 30070 19264
rect 30926 19252 30932 19264
rect 30984 19252 30990 19304
rect 33134 19292 33140 19304
rect 31496 19264 33140 19292
rect 31389 19227 31447 19233
rect 31389 19224 31401 19227
rect 28644 19196 31401 19224
rect 22066 19156 22094 19196
rect 31389 19193 31401 19196
rect 31435 19193 31447 19227
rect 31389 19187 31447 19193
rect 17236 19128 22094 19156
rect 24486 19116 24492 19168
rect 24544 19156 24550 19168
rect 26970 19156 26976 19168
rect 24544 19128 26976 19156
rect 24544 19116 24550 19128
rect 26970 19116 26976 19128
rect 27028 19116 27034 19168
rect 27062 19116 27068 19168
rect 27120 19156 27126 19168
rect 28534 19156 28540 19168
rect 27120 19128 28540 19156
rect 27120 19116 27126 19128
rect 28534 19116 28540 19128
rect 28592 19116 28598 19168
rect 28718 19116 28724 19168
rect 28776 19156 28782 19168
rect 30006 19156 30012 19168
rect 28776 19128 30012 19156
rect 28776 19116 28782 19128
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 30650 19116 30656 19168
rect 30708 19156 30714 19168
rect 31496 19156 31524 19264
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 33226 19252 33232 19304
rect 33284 19292 33290 19304
rect 33689 19295 33747 19301
rect 33689 19292 33701 19295
rect 33284 19264 33701 19292
rect 33284 19252 33290 19264
rect 33689 19261 33701 19264
rect 33735 19261 33747 19295
rect 36464 19292 36492 19323
rect 38286 19320 38292 19332
rect 38344 19320 38350 19372
rect 37458 19292 37464 19304
rect 36464 19264 37464 19292
rect 33689 19255 33747 19261
rect 37458 19252 37464 19264
rect 37516 19252 37522 19304
rect 31570 19184 31576 19236
rect 31628 19224 31634 19236
rect 33502 19224 33508 19236
rect 31628 19196 33508 19224
rect 31628 19184 31634 19196
rect 33502 19184 33508 19196
rect 33560 19184 33566 19236
rect 32398 19156 32404 19168
rect 30708 19128 31524 19156
rect 32359 19128 32404 19156
rect 30708 19116 30714 19128
rect 32398 19116 32404 19128
rect 32456 19116 32462 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 8389 18955 8447 18961
rect 8389 18921 8401 18955
rect 8435 18952 8447 18955
rect 10134 18952 10140 18964
rect 8435 18924 10140 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 12618 18952 12624 18964
rect 12579 18924 12624 18952
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 17037 18955 17095 18961
rect 17037 18921 17049 18955
rect 17083 18952 17095 18955
rect 17402 18952 17408 18964
rect 17083 18924 17408 18952
rect 17083 18921 17095 18924
rect 17037 18915 17095 18921
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 18598 18952 18604 18964
rect 18559 18924 18604 18952
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 19518 18952 19524 18964
rect 18708 18924 19524 18952
rect 10152 18816 10180 18912
rect 14642 18844 14648 18896
rect 14700 18884 14706 18896
rect 18708 18884 18736 18924
rect 19518 18912 19524 18924
rect 19576 18952 19582 18964
rect 19886 18952 19892 18964
rect 19576 18924 19892 18952
rect 19576 18912 19582 18924
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 24210 18912 24216 18964
rect 24268 18952 24274 18964
rect 24673 18955 24731 18961
rect 24673 18952 24685 18955
rect 24268 18924 24685 18952
rect 24268 18912 24274 18924
rect 24673 18921 24685 18924
rect 24719 18921 24731 18955
rect 24673 18915 24731 18921
rect 25958 18912 25964 18964
rect 26016 18952 26022 18964
rect 26016 18924 27384 18952
rect 26016 18912 26022 18924
rect 14700 18856 18736 18884
rect 14700 18844 14706 18856
rect 18874 18844 18880 18896
rect 18932 18884 18938 18896
rect 23477 18887 23535 18893
rect 23477 18884 23489 18887
rect 18932 18856 23489 18884
rect 18932 18844 18938 18856
rect 23477 18853 23489 18856
rect 23523 18884 23535 18887
rect 27246 18884 27252 18896
rect 23523 18856 27252 18884
rect 23523 18853 23535 18856
rect 23477 18847 23535 18853
rect 27246 18844 27252 18856
rect 27304 18844 27310 18896
rect 27356 18884 27384 18924
rect 28074 18912 28080 18964
rect 28132 18952 28138 18964
rect 29822 18952 29828 18964
rect 28132 18924 29828 18952
rect 28132 18912 28138 18924
rect 29822 18912 29828 18924
rect 29880 18912 29886 18964
rect 31018 18912 31024 18964
rect 31076 18952 31082 18964
rect 31076 18924 31754 18952
rect 31076 18912 31082 18924
rect 27430 18884 27436 18896
rect 27356 18856 27436 18884
rect 27430 18844 27436 18856
rect 27488 18844 27494 18896
rect 27522 18844 27528 18896
rect 27580 18884 27586 18896
rect 28994 18884 29000 18896
rect 27580 18856 29000 18884
rect 27580 18844 27586 18856
rect 28994 18844 29000 18856
rect 29052 18844 29058 18896
rect 31726 18884 31754 18924
rect 34422 18912 34428 18964
rect 34480 18952 34486 18964
rect 34977 18955 35035 18961
rect 34977 18952 34989 18955
rect 34480 18924 34989 18952
rect 34480 18912 34486 18924
rect 34977 18921 34989 18924
rect 35023 18921 35035 18955
rect 34977 18915 35035 18921
rect 34882 18884 34888 18896
rect 29840 18856 31248 18884
rect 31726 18856 34888 18884
rect 11057 18819 11115 18825
rect 11057 18816 11069 18819
rect 10152 18788 11069 18816
rect 11057 18785 11069 18788
rect 11103 18785 11115 18819
rect 11057 18779 11115 18785
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18816 12127 18819
rect 16574 18816 16580 18828
rect 12115 18788 16580 18816
rect 12115 18785 12127 18788
rect 12069 18779 12127 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 18598 18816 18604 18828
rect 16960 18788 18604 18816
rect 6546 18748 6552 18760
rect 6507 18720 6552 18748
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 8294 18748 8300 18760
rect 8255 18720 8300 18748
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 12529 18751 12587 18757
rect 12529 18748 12541 18751
rect 12406 18720 12541 18748
rect 11146 18680 11152 18692
rect 11107 18652 11152 18680
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 11238 18640 11244 18692
rect 11296 18680 11302 18692
rect 12406 18680 12434 18720
rect 12529 18717 12541 18720
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18748 13231 18751
rect 15562 18748 15568 18760
rect 13219 18720 15568 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16114 18748 16120 18760
rect 15979 18720 16120 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16114 18708 16120 18720
rect 16172 18748 16178 18760
rect 16960 18757 16988 18788
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 19334 18776 19340 18828
rect 19392 18776 19398 18828
rect 19521 18819 19579 18825
rect 19521 18785 19533 18819
rect 19567 18816 19579 18819
rect 22925 18819 22983 18825
rect 22925 18816 22937 18819
rect 19567 18788 22937 18816
rect 19567 18785 19579 18788
rect 19521 18779 19579 18785
rect 22925 18785 22937 18788
rect 22971 18816 22983 18819
rect 23198 18816 23204 18828
rect 22971 18788 23204 18816
rect 22971 18785 22983 18788
rect 22925 18779 22983 18785
rect 23198 18776 23204 18788
rect 23256 18776 23262 18828
rect 29840 18825 29868 18856
rect 29825 18819 29883 18825
rect 29825 18785 29837 18819
rect 29871 18785 29883 18819
rect 29825 18779 29883 18785
rect 30469 18819 30527 18825
rect 30469 18785 30481 18819
rect 30515 18816 30527 18819
rect 31110 18816 31116 18828
rect 30515 18788 31116 18816
rect 30515 18785 30527 18788
rect 30469 18779 30527 18785
rect 31110 18776 31116 18788
rect 31168 18776 31174 18828
rect 31220 18816 31248 18856
rect 34882 18844 34888 18856
rect 34940 18844 34946 18896
rect 31662 18816 31668 18828
rect 31220 18788 31668 18816
rect 31662 18776 31668 18788
rect 31720 18816 31726 18828
rect 32769 18819 32827 18825
rect 32769 18816 32781 18819
rect 31720 18788 32781 18816
rect 31720 18776 31726 18788
rect 32769 18785 32781 18788
rect 32815 18785 32827 18819
rect 33134 18816 33140 18828
rect 33095 18788 33140 18816
rect 32769 18779 32827 18785
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 35894 18776 35900 18828
rect 35952 18816 35958 18828
rect 38562 18816 38568 18828
rect 35952 18788 38568 18816
rect 35952 18776 35958 18788
rect 38562 18776 38568 18788
rect 38620 18776 38626 18828
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16172 18720 16957 18748
rect 16172 18708 16178 18720
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18104 18720 18521 18748
rect 18104 18708 18110 18720
rect 18509 18717 18521 18720
rect 18555 18748 18567 18751
rect 19058 18748 19064 18760
rect 18555 18720 19064 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 11296 18652 12434 18680
rect 19352 18680 19380 18776
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18748 21603 18751
rect 21634 18748 21640 18760
rect 21591 18720 21640 18748
rect 21591 18717 21603 18720
rect 21545 18711 21603 18717
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 19352 18652 19625 18680
rect 11296 18640 11302 18652
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 19613 18643 19671 18649
rect 19886 18640 19892 18692
rect 19944 18680 19950 18692
rect 20165 18683 20223 18689
rect 20165 18680 20177 18683
rect 19944 18652 20177 18680
rect 19944 18640 19950 18652
rect 20165 18649 20177 18652
rect 20211 18649 20223 18683
rect 20640 18680 20668 18711
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 22066 18720 22201 18748
rect 22066 18680 22094 18720
rect 22189 18717 22201 18720
rect 22235 18748 22247 18751
rect 22278 18748 22284 18760
rect 22235 18720 22284 18748
rect 22235 18717 22247 18720
rect 22189 18711 22247 18717
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 24486 18708 24492 18760
rect 24544 18748 24550 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24544 18720 24593 18748
rect 24544 18708 24550 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 28258 18708 28264 18760
rect 28316 18748 28322 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28316 18720 28825 18748
rect 28316 18708 28322 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 34698 18708 34704 18760
rect 34756 18748 34762 18760
rect 34885 18751 34943 18757
rect 34885 18748 34897 18751
rect 34756 18720 34897 18748
rect 34756 18708 34762 18720
rect 34885 18717 34897 18720
rect 34931 18748 34943 18751
rect 38838 18748 38844 18760
rect 34931 18720 38844 18748
rect 34931 18717 34943 18720
rect 34885 18711 34943 18717
rect 38838 18708 38844 18720
rect 38896 18708 38902 18760
rect 20165 18643 20223 18649
rect 20272 18652 22094 18680
rect 6641 18615 6699 18621
rect 6641 18581 6653 18615
rect 6687 18612 6699 18615
rect 8570 18612 8576 18624
rect 6687 18584 8576 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 9732 18584 13277 18612
rect 9732 18572 9738 18584
rect 13265 18581 13277 18584
rect 13311 18581 13323 18615
rect 16022 18612 16028 18624
rect 15983 18584 16028 18612
rect 13265 18575 13323 18581
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 20272 18612 20300 18652
rect 23014 18640 23020 18692
rect 23072 18680 23078 18692
rect 25774 18680 25780 18692
rect 23072 18652 23117 18680
rect 25735 18652 25780 18680
rect 23072 18640 23078 18652
rect 25774 18640 25780 18652
rect 25832 18640 25838 18692
rect 25869 18683 25927 18689
rect 25869 18649 25881 18683
rect 25915 18649 25927 18683
rect 25869 18643 25927 18649
rect 20714 18612 20720 18624
rect 16172 18584 20300 18612
rect 20675 18584 20720 18612
rect 16172 18572 16178 18584
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 21637 18615 21695 18621
rect 21637 18581 21649 18615
rect 21683 18612 21695 18615
rect 21910 18612 21916 18624
rect 21683 18584 21916 18612
rect 21683 18581 21695 18584
rect 21637 18575 21695 18581
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 22281 18615 22339 18621
rect 22281 18581 22293 18615
rect 22327 18612 22339 18615
rect 22830 18612 22836 18624
rect 22327 18584 22836 18612
rect 22327 18581 22339 18584
rect 22281 18575 22339 18581
rect 22830 18572 22836 18584
rect 22888 18572 22894 18624
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 25682 18612 25688 18624
rect 23716 18584 25688 18612
rect 23716 18572 23722 18584
rect 25682 18572 25688 18584
rect 25740 18572 25746 18624
rect 25884 18612 25912 18643
rect 26694 18640 26700 18692
rect 26752 18680 26758 18692
rect 26789 18683 26847 18689
rect 26789 18680 26801 18683
rect 26752 18652 26801 18680
rect 26752 18640 26758 18652
rect 26789 18649 26801 18652
rect 26835 18649 26847 18683
rect 27338 18680 27344 18692
rect 27299 18652 27344 18680
rect 26789 18643 26847 18649
rect 27338 18640 27344 18652
rect 27396 18640 27402 18692
rect 27430 18640 27436 18692
rect 27488 18680 27494 18692
rect 27488 18652 27533 18680
rect 27488 18640 27494 18652
rect 27614 18640 27620 18692
rect 27672 18680 27678 18692
rect 27982 18680 27988 18692
rect 27672 18652 27988 18680
rect 27672 18640 27678 18652
rect 27982 18640 27988 18652
rect 28040 18680 28046 18692
rect 28353 18683 28411 18689
rect 28353 18680 28365 18683
rect 28040 18652 28365 18680
rect 28040 18640 28046 18652
rect 28353 18649 28365 18652
rect 28399 18649 28411 18683
rect 28353 18643 28411 18649
rect 28534 18640 28540 18692
rect 28592 18680 28598 18692
rect 28592 18652 29868 18680
rect 28592 18640 28598 18652
rect 27890 18612 27896 18624
rect 25884 18584 27896 18612
rect 27890 18572 27896 18584
rect 27948 18572 27954 18624
rect 28718 18572 28724 18624
rect 28776 18612 28782 18624
rect 28905 18615 28963 18621
rect 28905 18612 28917 18615
rect 28776 18584 28917 18612
rect 28776 18572 28782 18584
rect 28905 18581 28917 18584
rect 28951 18581 28963 18615
rect 29840 18612 29868 18652
rect 29914 18640 29920 18692
rect 29972 18680 29978 18692
rect 29972 18652 30017 18680
rect 29972 18640 29978 18652
rect 30650 18640 30656 18692
rect 30708 18680 30714 18692
rect 31018 18680 31024 18692
rect 30708 18652 31024 18680
rect 30708 18640 30714 18652
rect 31018 18640 31024 18652
rect 31076 18640 31082 18692
rect 31113 18683 31171 18689
rect 31113 18649 31125 18683
rect 31159 18649 31171 18683
rect 31113 18643 31171 18649
rect 31665 18683 31723 18689
rect 31665 18649 31677 18683
rect 31711 18680 31723 18683
rect 32030 18680 32036 18692
rect 31711 18652 32036 18680
rect 31711 18649 31723 18652
rect 31665 18643 31723 18649
rect 30926 18612 30932 18624
rect 29840 18584 30932 18612
rect 28905 18575 28963 18581
rect 30926 18572 30932 18584
rect 30984 18572 30990 18624
rect 31128 18612 31156 18643
rect 32030 18640 32036 18652
rect 32088 18640 32094 18692
rect 32861 18683 32919 18689
rect 32861 18649 32873 18683
rect 32907 18680 32919 18683
rect 34054 18680 34060 18692
rect 32907 18652 34060 18680
rect 32907 18649 32919 18652
rect 32861 18643 32919 18649
rect 34054 18640 34060 18652
rect 34112 18640 34118 18692
rect 32306 18612 32312 18624
rect 31128 18584 32312 18612
rect 32306 18572 32312 18584
rect 32364 18572 32370 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 8294 18408 8300 18420
rect 1627 18380 8300 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 11572 18380 13277 18408
rect 11572 18368 11578 18380
rect 13265 18377 13277 18380
rect 13311 18377 13323 18411
rect 15654 18408 15660 18420
rect 15615 18380 15660 18408
rect 13265 18371 13323 18377
rect 15654 18368 15660 18380
rect 15712 18368 15718 18420
rect 23658 18408 23664 18420
rect 15751 18380 23664 18408
rect 6730 18340 6736 18352
rect 6691 18312 6736 18340
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 12158 18340 12164 18352
rect 12119 18312 12164 18340
rect 12158 18300 12164 18312
rect 12216 18300 12222 18352
rect 12710 18340 12716 18352
rect 12671 18312 12716 18340
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 13906 18340 13912 18352
rect 12952 18312 13912 18340
rect 12952 18300 12958 18312
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 15102 18300 15108 18352
rect 15160 18340 15166 18352
rect 15751 18340 15779 18380
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 25958 18408 25964 18420
rect 23860 18380 25964 18408
rect 18046 18340 18052 18352
rect 15160 18312 15779 18340
rect 18007 18312 18052 18340
rect 15160 18300 15166 18312
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 18138 18300 18144 18352
rect 18196 18340 18202 18352
rect 18196 18312 18828 18340
rect 18196 18300 18202 18312
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 9033 18275 9091 18281
rect 9033 18272 9045 18275
rect 8076 18244 9045 18272
rect 8076 18232 8082 18244
rect 9033 18241 9045 18244
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18272 17279 18275
rect 17586 18272 17592 18284
rect 17267 18244 17592 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 6086 18164 6092 18216
rect 6144 18204 6150 18216
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6144 18176 6653 18204
rect 6144 18164 6150 18176
rect 6641 18173 6653 18176
rect 6687 18173 6699 18207
rect 7650 18204 7656 18216
rect 7611 18176 7656 18204
rect 6641 18167 6699 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8938 18164 8944 18216
rect 8996 18204 9002 18216
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 8996 18176 12081 18204
rect 8996 18164 9002 18176
rect 12069 18173 12081 18176
rect 12115 18173 12127 18207
rect 13188 18204 13216 18235
rect 12069 18167 12127 18173
rect 12406 18176 13216 18204
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 12406 18136 12434 18176
rect 15580 18136 15608 18235
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18204 18015 18207
rect 18322 18204 18328 18216
rect 18003 18176 18184 18204
rect 18283 18176 18328 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 11204 18108 12434 18136
rect 12728 18108 15608 18136
rect 18156 18136 18184 18176
rect 18322 18164 18328 18176
rect 18380 18164 18386 18216
rect 18800 18204 18828 18312
rect 19886 18300 19892 18352
rect 19944 18340 19950 18352
rect 20257 18343 20315 18349
rect 20257 18340 20269 18343
rect 19944 18312 20269 18340
rect 19944 18300 19950 18312
rect 20257 18309 20269 18312
rect 20303 18309 20315 18343
rect 20257 18303 20315 18309
rect 20349 18343 20407 18349
rect 20349 18309 20361 18343
rect 20395 18340 20407 18343
rect 21082 18340 21088 18352
rect 20395 18312 21088 18340
rect 20395 18309 20407 18312
rect 20349 18303 20407 18309
rect 21082 18300 21088 18312
rect 21140 18300 21146 18352
rect 23860 18349 23888 18380
rect 25958 18368 25964 18380
rect 26016 18368 26022 18420
rect 28626 18368 28632 18420
rect 28684 18408 28690 18420
rect 28684 18380 28764 18408
rect 28684 18368 28690 18380
rect 23845 18343 23903 18349
rect 23845 18309 23857 18343
rect 23891 18309 23903 18343
rect 23845 18303 23903 18309
rect 23937 18343 23995 18349
rect 23937 18309 23949 18343
rect 23983 18340 23995 18343
rect 25314 18340 25320 18352
rect 23983 18312 25320 18340
rect 23983 18309 23995 18312
rect 23937 18303 23995 18309
rect 25314 18300 25320 18312
rect 25372 18300 25378 18352
rect 26053 18343 26111 18349
rect 26053 18309 26065 18343
rect 26099 18340 26111 18343
rect 26326 18340 26332 18352
rect 26099 18312 26332 18340
rect 26099 18309 26111 18312
rect 26053 18303 26111 18309
rect 26326 18300 26332 18312
rect 26384 18300 26390 18352
rect 27246 18300 27252 18352
rect 27304 18340 27310 18352
rect 28736 18349 28764 18380
rect 28902 18368 28908 18420
rect 28960 18408 28966 18420
rect 30282 18408 30288 18420
rect 28960 18380 30288 18408
rect 28960 18368 28966 18380
rect 30282 18368 30288 18380
rect 30340 18368 30346 18420
rect 30926 18368 30932 18420
rect 30984 18408 30990 18420
rect 33597 18411 33655 18417
rect 30984 18380 32444 18408
rect 30984 18368 30990 18380
rect 27341 18343 27399 18349
rect 27341 18340 27353 18343
rect 27304 18312 27353 18340
rect 27304 18300 27310 18312
rect 27341 18309 27353 18312
rect 27387 18309 27399 18343
rect 27341 18303 27399 18309
rect 28721 18343 28779 18349
rect 28721 18309 28733 18343
rect 28767 18309 28779 18343
rect 28721 18303 28779 18309
rect 28810 18300 28816 18352
rect 28868 18340 28874 18352
rect 29638 18340 29644 18352
rect 28868 18312 29644 18340
rect 28868 18300 28874 18312
rect 29638 18300 29644 18312
rect 29696 18300 29702 18352
rect 32416 18349 32444 18380
rect 33597 18377 33609 18411
rect 33643 18408 33655 18411
rect 33962 18408 33968 18420
rect 33643 18380 33968 18408
rect 33643 18377 33655 18380
rect 33597 18371 33655 18377
rect 33962 18368 33968 18380
rect 34020 18368 34026 18420
rect 34882 18408 34888 18420
rect 34843 18380 34888 18408
rect 34882 18368 34888 18380
rect 34940 18368 34946 18420
rect 31021 18343 31079 18349
rect 31021 18340 31033 18343
rect 29932 18312 31033 18340
rect 19429 18275 19487 18281
rect 19429 18241 19441 18275
rect 19475 18272 19487 18275
rect 20070 18272 20076 18284
rect 19475 18244 20076 18272
rect 19475 18241 19487 18244
rect 19429 18235 19487 18241
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18241 22339 18275
rect 22281 18235 22339 18241
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18272 22983 18275
rect 23658 18272 23664 18284
rect 22971 18244 23664 18272
rect 22971 18241 22983 18244
rect 22925 18235 22983 18241
rect 22296 18204 22324 18235
rect 23658 18232 23664 18244
rect 23716 18232 23722 18284
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18272 27951 18275
rect 28534 18272 28540 18284
rect 27939 18244 28396 18272
rect 28495 18244 28540 18272
rect 27939 18241 27951 18244
rect 27893 18235 27951 18241
rect 23198 18204 23204 18216
rect 18800 18176 22094 18204
rect 22296 18176 23204 18204
rect 20346 18136 20352 18148
rect 18156 18108 20352 18136
rect 11204 18096 11210 18108
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9306 18068 9312 18080
rect 9171 18040 9312 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 10134 18068 10140 18080
rect 9456 18040 10140 18068
rect 9456 18028 9462 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 12728 18068 12756 18108
rect 20346 18096 20352 18108
rect 20404 18096 20410 18148
rect 20809 18139 20867 18145
rect 20809 18105 20821 18139
rect 20855 18105 20867 18139
rect 22066 18136 22094 18176
rect 23198 18164 23204 18176
rect 23256 18164 23262 18216
rect 24762 18204 24768 18216
rect 24723 18176 24768 18204
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 25961 18207 26019 18213
rect 25961 18173 25973 18207
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 27249 18207 27307 18213
rect 27249 18173 27261 18207
rect 27295 18204 27307 18207
rect 28074 18204 28080 18216
rect 27295 18176 28080 18204
rect 27295 18173 27307 18176
rect 27249 18167 27307 18173
rect 25976 18136 26004 18167
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 28368 18204 28396 18244
rect 28534 18232 28540 18244
rect 28592 18232 28598 18284
rect 28276 18176 28856 18204
rect 22066 18108 26004 18136
rect 20809 18099 20867 18105
rect 10652 18040 12756 18068
rect 17313 18071 17371 18077
rect 10652 18028 10658 18040
rect 17313 18037 17325 18071
rect 17359 18068 17371 18071
rect 18322 18068 18328 18080
rect 17359 18040 18328 18068
rect 17359 18037 17371 18040
rect 17313 18031 17371 18037
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19426 18068 19432 18080
rect 18656 18040 19432 18068
rect 18656 18028 18662 18040
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 19521 18071 19579 18077
rect 19521 18037 19533 18071
rect 19567 18068 19579 18071
rect 20070 18068 20076 18080
rect 19567 18040 20076 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20824 18068 20852 18099
rect 20772 18040 20852 18068
rect 20772 18028 20778 18040
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 22373 18071 22431 18077
rect 22373 18068 22385 18071
rect 22244 18040 22385 18068
rect 22244 18028 22250 18040
rect 22373 18037 22385 18040
rect 22419 18037 22431 18071
rect 23014 18068 23020 18080
rect 22975 18040 23020 18068
rect 22373 18031 22431 18037
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 25976 18068 26004 18108
rect 26513 18139 26571 18145
rect 26513 18105 26525 18139
rect 26559 18136 26571 18139
rect 28276 18136 28304 18176
rect 26559 18108 28304 18136
rect 28828 18136 28856 18176
rect 28902 18164 28908 18216
rect 28960 18204 28966 18216
rect 29932 18204 29960 18312
rect 31021 18309 31033 18312
rect 31067 18309 31079 18343
rect 31021 18303 31079 18309
rect 32401 18343 32459 18349
rect 32401 18309 32413 18343
rect 32447 18309 32459 18343
rect 32401 18303 32459 18309
rect 32493 18343 32551 18349
rect 32493 18309 32505 18343
rect 32539 18340 32551 18343
rect 34241 18343 34299 18349
rect 34241 18340 34253 18343
rect 32539 18312 34253 18340
rect 32539 18309 32551 18312
rect 32493 18303 32551 18309
rect 34241 18309 34253 18312
rect 34287 18309 34299 18343
rect 37458 18340 37464 18352
rect 34241 18303 34299 18309
rect 34808 18312 37464 18340
rect 33042 18232 33048 18284
rect 33100 18272 33106 18284
rect 33502 18272 33508 18284
rect 33100 18244 33364 18272
rect 33463 18244 33508 18272
rect 33100 18232 33106 18244
rect 30190 18204 30196 18216
rect 28960 18176 29960 18204
rect 30151 18176 30196 18204
rect 28960 18164 28966 18176
rect 30190 18164 30196 18176
rect 30248 18164 30254 18216
rect 30929 18207 30987 18213
rect 30929 18173 30941 18207
rect 30975 18204 30987 18207
rect 31110 18204 31116 18216
rect 30975 18176 31116 18204
rect 30975 18173 30987 18176
rect 30929 18167 30987 18173
rect 31110 18164 31116 18176
rect 31168 18164 31174 18216
rect 31570 18164 31576 18216
rect 31628 18204 31634 18216
rect 32030 18204 32036 18216
rect 31628 18176 32036 18204
rect 31628 18164 31634 18176
rect 32030 18164 32036 18176
rect 32088 18204 32094 18216
rect 32677 18207 32735 18213
rect 32677 18204 32689 18207
rect 32088 18176 32689 18204
rect 32088 18164 32094 18176
rect 32677 18173 32689 18176
rect 32723 18173 32735 18207
rect 33336 18204 33364 18244
rect 33502 18232 33508 18244
rect 33560 18232 33566 18284
rect 34808 18281 34836 18312
rect 37458 18300 37464 18312
rect 37516 18300 37522 18352
rect 34149 18275 34207 18281
rect 34149 18241 34161 18275
rect 34195 18241 34207 18275
rect 34149 18235 34207 18241
rect 34793 18275 34851 18281
rect 34793 18241 34805 18275
rect 34839 18241 34851 18275
rect 35618 18272 35624 18284
rect 35579 18244 35624 18272
rect 34793 18235 34851 18241
rect 34164 18204 34192 18235
rect 35618 18232 35624 18244
rect 35676 18232 35682 18284
rect 38102 18272 38108 18284
rect 38063 18244 38108 18272
rect 38102 18232 38108 18244
rect 38160 18232 38166 18284
rect 33336 18176 34192 18204
rect 32677 18167 32735 18173
rect 31481 18139 31539 18145
rect 31481 18136 31493 18139
rect 28828 18108 31493 18136
rect 26559 18105 26571 18108
rect 26513 18099 26571 18105
rect 31481 18105 31493 18108
rect 31527 18136 31539 18139
rect 33226 18136 33232 18148
rect 31527 18108 33232 18136
rect 31527 18105 31539 18108
rect 31481 18099 31539 18105
rect 33226 18096 33232 18108
rect 33284 18096 33290 18148
rect 37274 18096 37280 18148
rect 37332 18136 37338 18148
rect 38289 18139 38347 18145
rect 38289 18136 38301 18139
rect 37332 18108 38301 18136
rect 37332 18096 37338 18108
rect 38289 18105 38301 18108
rect 38335 18105 38347 18139
rect 38289 18099 38347 18105
rect 27522 18068 27528 18080
rect 25976 18040 27528 18068
rect 27522 18028 27528 18040
rect 27580 18028 27586 18080
rect 27890 18028 27896 18080
rect 27948 18068 27954 18080
rect 28258 18068 28264 18080
rect 27948 18040 28264 18068
rect 27948 18028 27954 18040
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 28626 18028 28632 18080
rect 28684 18068 28690 18080
rect 32766 18068 32772 18080
rect 28684 18040 32772 18068
rect 28684 18028 28690 18040
rect 32766 18028 32772 18040
rect 32824 18028 32830 18080
rect 35437 18071 35495 18077
rect 35437 18037 35449 18071
rect 35483 18068 35495 18071
rect 37918 18068 37924 18080
rect 35483 18040 37924 18068
rect 35483 18037 35495 18040
rect 35437 18031 35495 18037
rect 37918 18028 37924 18040
rect 37976 18028 37982 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6730 17864 6736 17876
rect 6595 17836 6736 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 15010 17824 15016 17876
rect 15068 17864 15074 17876
rect 16482 17864 16488 17876
rect 15068 17836 16488 17864
rect 15068 17824 15074 17836
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 20806 17864 20812 17876
rect 16632 17836 20812 17864
rect 16632 17824 16638 17836
rect 20806 17824 20812 17836
rect 20864 17824 20870 17876
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21450 17824 21456 17876
rect 21508 17864 21514 17876
rect 21508 17836 32720 17864
rect 21508 17824 21514 17836
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 11698 17796 11704 17808
rect 9456 17768 11704 17796
rect 9456 17756 9462 17768
rect 11698 17756 11704 17768
rect 11756 17756 11762 17808
rect 15102 17796 15108 17808
rect 13188 17768 15108 17796
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 13188 17737 13216 17768
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 15378 17756 15384 17808
rect 15436 17796 15442 17808
rect 25682 17796 25688 17808
rect 15436 17768 25688 17796
rect 15436 17756 15442 17768
rect 25682 17756 25688 17768
rect 25740 17756 25746 17808
rect 25774 17756 25780 17808
rect 25832 17796 25838 17808
rect 26602 17796 26608 17808
rect 25832 17768 26608 17796
rect 25832 17756 25838 17768
rect 26602 17756 26608 17768
rect 26660 17796 26666 17808
rect 27338 17796 27344 17808
rect 26660 17768 26832 17796
rect 27299 17768 27344 17796
rect 26660 17756 26666 17768
rect 9217 17731 9275 17737
rect 9217 17728 9229 17731
rect 8628 17700 9229 17728
rect 8628 17688 8634 17700
rect 9217 17697 9229 17700
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17697 13231 17731
rect 13173 17691 13231 17697
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 16485 17731 16543 17737
rect 16485 17728 16497 17731
rect 14976 17700 16497 17728
rect 14976 17688 14982 17700
rect 16485 17697 16497 17700
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 17497 17731 17555 17737
rect 16632 17700 17448 17728
rect 16632 17688 16638 17700
rect 6457 17663 6515 17669
rect 6457 17629 6469 17663
rect 6503 17660 6515 17663
rect 7101 17663 7159 17669
rect 7101 17660 7113 17663
rect 6503 17632 7113 17660
rect 6503 17629 6515 17632
rect 6457 17623 6515 17629
rect 7101 17629 7113 17632
rect 7147 17660 7159 17663
rect 7742 17660 7748 17672
rect 7147 17632 7748 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17660 8447 17663
rect 8754 17660 8760 17672
rect 8435 17632 8760 17660
rect 8435 17629 8447 17632
rect 8389 17623 8447 17629
rect 8754 17620 8760 17632
rect 8812 17620 8818 17672
rect 10594 17620 10600 17672
rect 10652 17660 10658 17672
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 10652 17632 10793 17660
rect 10652 17620 10658 17632
rect 10781 17629 10793 17632
rect 10827 17629 10839 17663
rect 11422 17660 11428 17672
rect 11383 17632 11428 17660
rect 10781 17623 10839 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15470 17660 15476 17672
rect 15151 17632 15476 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 7837 17595 7895 17601
rect 7837 17561 7849 17595
rect 7883 17592 7895 17595
rect 9030 17592 9036 17604
rect 7883 17564 9036 17592
rect 7883 17561 7895 17564
rect 7837 17555 7895 17561
rect 9030 17552 9036 17564
rect 9088 17552 9094 17604
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 9364 17564 9409 17592
rect 9364 17552 9370 17564
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9732 17564 9873 17592
rect 9732 17552 9738 17564
rect 9861 17561 9873 17564
rect 9907 17592 9919 17595
rect 9907 17564 11652 17592
rect 9907 17561 9919 17564
rect 9861 17555 9919 17561
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 7064 17496 7205 17524
rect 7064 17484 7070 17496
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8260 17496 8493 17524
rect 8260 17484 8266 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 8481 17487 8539 17493
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11514 17524 11520 17536
rect 11475 17496 11520 17524
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11624 17524 11652 17564
rect 11790 17552 11796 17604
rect 11848 17592 11854 17604
rect 12161 17595 12219 17601
rect 12161 17592 12173 17595
rect 11848 17564 12173 17592
rect 11848 17552 11854 17564
rect 12161 17561 12173 17564
rect 12207 17561 12219 17595
rect 12161 17555 12219 17561
rect 12253 17595 12311 17601
rect 12253 17561 12265 17595
rect 12299 17592 12311 17595
rect 12986 17592 12992 17604
rect 12299 17564 12992 17592
rect 12299 17561 12311 17564
rect 12253 17555 12311 17561
rect 12986 17552 12992 17564
rect 13044 17552 13050 17604
rect 14292 17592 14320 17623
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 16114 17660 16120 17672
rect 15795 17632 16120 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 17420 17660 17448 17700
rect 17497 17697 17509 17731
rect 17543 17728 17555 17731
rect 24486 17728 24492 17740
rect 17543 17700 24492 17728
rect 17543 17697 17555 17700
rect 17497 17691 17555 17697
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 24673 17731 24731 17737
rect 24673 17697 24685 17731
rect 24719 17728 24731 17731
rect 26050 17728 26056 17740
rect 24719 17700 26056 17728
rect 24719 17697 24731 17700
rect 24673 17691 24731 17697
rect 26050 17688 26056 17700
rect 26108 17688 26114 17740
rect 26804 17737 26832 17768
rect 27338 17756 27344 17768
rect 27396 17756 27402 17808
rect 32398 17796 32404 17808
rect 27816 17768 32404 17796
rect 26789 17731 26847 17737
rect 26789 17697 26801 17731
rect 26835 17697 26847 17731
rect 26789 17691 26847 17697
rect 27154 17688 27160 17740
rect 27212 17728 27218 17740
rect 27706 17728 27712 17740
rect 27212 17700 27712 17728
rect 27212 17688 27218 17700
rect 27706 17688 27712 17700
rect 27764 17688 27770 17740
rect 18049 17663 18107 17669
rect 18049 17660 18061 17663
rect 17420 17632 18061 17660
rect 18049 17629 18061 17632
rect 18095 17629 18107 17663
rect 18690 17660 18696 17672
rect 18651 17632 18696 17660
rect 18049 17623 18107 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19518 17660 19524 17672
rect 19260 17632 19524 17660
rect 16482 17592 16488 17604
rect 14292 17564 16488 17592
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 16577 17595 16635 17601
rect 16577 17561 16589 17595
rect 16623 17561 16635 17595
rect 16577 17555 16635 17561
rect 13722 17524 13728 17536
rect 11624 17496 13728 17524
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 14366 17524 14372 17536
rect 14327 17496 14372 17524
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 15197 17527 15255 17533
rect 15197 17493 15209 17527
rect 15243 17524 15255 17527
rect 15286 17524 15292 17536
rect 15243 17496 15292 17524
rect 15243 17493 15255 17496
rect 15197 17487 15255 17493
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 15838 17524 15844 17536
rect 15799 17496 15844 17524
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 16592 17524 16620 17555
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 19260 17592 19288 17632
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21542 17660 21548 17672
rect 21039 17632 21548 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17660 23351 17663
rect 23566 17660 23572 17672
rect 23339 17632 23572 17660
rect 23339 17629 23351 17632
rect 23293 17623 23351 17629
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 16908 17564 19288 17592
rect 16908 17552 16914 17564
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 19392 17564 19717 17592
rect 19392 17552 19398 17564
rect 19705 17561 19717 17564
rect 19751 17561 19763 17595
rect 19705 17555 19763 17561
rect 19797 17595 19855 17601
rect 19797 17561 19809 17595
rect 19843 17561 19855 17595
rect 19797 17555 19855 17561
rect 20349 17595 20407 17601
rect 20349 17561 20361 17595
rect 20395 17592 20407 17595
rect 20714 17592 20720 17604
rect 20395 17564 20720 17592
rect 20395 17561 20407 17564
rect 20349 17555 20407 17561
rect 18138 17524 18144 17536
rect 16080 17496 16620 17524
rect 18099 17496 18144 17524
rect 16080 17484 16086 17496
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 18785 17527 18843 17533
rect 18785 17493 18797 17527
rect 18831 17524 18843 17527
rect 19812 17524 19840 17555
rect 20714 17552 20720 17564
rect 20772 17552 20778 17604
rect 20806 17552 20812 17604
rect 20864 17592 20870 17604
rect 21821 17595 21879 17601
rect 21821 17592 21833 17595
rect 20864 17564 21833 17592
rect 20864 17552 20870 17564
rect 21821 17561 21833 17564
rect 21867 17561 21879 17595
rect 21821 17555 21879 17561
rect 21910 17552 21916 17604
rect 21968 17592 21974 17604
rect 22833 17595 22891 17601
rect 21968 17564 22013 17592
rect 21968 17552 21974 17564
rect 22833 17561 22845 17595
rect 22879 17592 22891 17595
rect 24670 17592 24676 17604
rect 22879 17564 24676 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 24670 17552 24676 17564
rect 24728 17552 24734 17604
rect 24765 17595 24823 17601
rect 24765 17561 24777 17595
rect 24811 17592 24823 17595
rect 25590 17592 25596 17604
rect 24811 17564 25596 17592
rect 24811 17561 24823 17564
rect 24765 17555 24823 17561
rect 25590 17552 25596 17564
rect 25648 17552 25654 17604
rect 25682 17552 25688 17604
rect 25740 17592 25746 17604
rect 26881 17595 26939 17601
rect 25740 17564 25785 17592
rect 25740 17552 25746 17564
rect 26881 17561 26893 17595
rect 26927 17592 26939 17595
rect 27816 17592 27844 17768
rect 32398 17756 32404 17768
rect 32456 17756 32462 17808
rect 28258 17688 28264 17740
rect 28316 17728 28322 17740
rect 28629 17731 28687 17737
rect 28629 17728 28641 17731
rect 28316 17700 28641 17728
rect 28316 17688 28322 17700
rect 28629 17697 28641 17700
rect 28675 17697 28687 17731
rect 28629 17691 28687 17697
rect 29730 17688 29736 17740
rect 29788 17728 29794 17740
rect 29788 17700 32628 17728
rect 29788 17688 29794 17700
rect 27893 17663 27951 17669
rect 27893 17629 27905 17663
rect 27939 17660 27951 17663
rect 28442 17660 28448 17672
rect 27939 17632 28448 17660
rect 27939 17629 27951 17632
rect 27893 17623 27951 17629
rect 28442 17620 28448 17632
rect 28500 17620 28506 17672
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 26927 17564 27844 17592
rect 26927 17561 26939 17564
rect 26881 17555 26939 17561
rect 18831 17496 19840 17524
rect 18831 17493 18843 17496
rect 18785 17487 18843 17493
rect 19886 17484 19892 17536
rect 19944 17524 19950 17536
rect 21450 17524 21456 17536
rect 19944 17496 21456 17524
rect 19944 17484 19950 17496
rect 21450 17484 21456 17496
rect 21508 17524 21514 17536
rect 21726 17524 21732 17536
rect 21508 17496 21732 17524
rect 21508 17484 21514 17496
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 23385 17527 23443 17533
rect 23385 17524 23397 17527
rect 22612 17496 23397 17524
rect 22612 17484 22618 17496
rect 23385 17493 23397 17496
rect 23431 17493 23443 17527
rect 23385 17487 23443 17493
rect 23934 17484 23940 17536
rect 23992 17524 23998 17536
rect 27985 17527 28043 17533
rect 27985 17524 27997 17527
rect 23992 17496 27997 17524
rect 23992 17484 23998 17496
rect 27985 17493 27997 17496
rect 28031 17493 28043 17527
rect 28552 17524 28580 17623
rect 30926 17620 30932 17672
rect 30984 17660 30990 17672
rect 30984 17632 31432 17660
rect 30984 17620 30990 17632
rect 30006 17592 30012 17604
rect 29967 17564 30012 17592
rect 30006 17552 30012 17564
rect 30064 17552 30070 17604
rect 30098 17552 30104 17604
rect 30156 17592 30162 17604
rect 30156 17564 30201 17592
rect 30156 17552 30162 17564
rect 30466 17552 30472 17604
rect 30524 17592 30530 17604
rect 31021 17595 31079 17601
rect 31021 17592 31033 17595
rect 30524 17564 31033 17592
rect 30524 17552 30530 17564
rect 31021 17561 31033 17564
rect 31067 17592 31079 17595
rect 31294 17592 31300 17604
rect 31067 17564 31300 17592
rect 31067 17561 31079 17564
rect 31021 17555 31079 17561
rect 31294 17552 31300 17564
rect 31352 17552 31358 17604
rect 31404 17592 31432 17632
rect 31570 17592 31576 17604
rect 31404 17564 31576 17592
rect 31570 17552 31576 17564
rect 31628 17552 31634 17604
rect 31665 17595 31723 17601
rect 31665 17561 31677 17595
rect 31711 17561 31723 17595
rect 31665 17555 31723 17561
rect 31110 17524 31116 17536
rect 28552 17496 31116 17524
rect 27985 17487 28043 17493
rect 31110 17484 31116 17496
rect 31168 17484 31174 17536
rect 31680 17524 31708 17555
rect 31846 17552 31852 17604
rect 31904 17592 31910 17604
rect 32214 17592 32220 17604
rect 31904 17564 32220 17592
rect 31904 17552 31910 17564
rect 32214 17552 32220 17564
rect 32272 17552 32278 17604
rect 32600 17592 32628 17700
rect 32692 17669 32720 17836
rect 32766 17824 32772 17876
rect 32824 17864 32830 17876
rect 32824 17836 32869 17864
rect 32824 17824 32830 17836
rect 32858 17756 32864 17808
rect 32916 17796 32922 17808
rect 34514 17796 34520 17808
rect 32916 17768 34520 17796
rect 32916 17756 32922 17768
rect 34514 17756 34520 17768
rect 34572 17756 34578 17808
rect 33226 17688 33232 17740
rect 33284 17728 33290 17740
rect 33284 17700 34928 17728
rect 33284 17688 33290 17700
rect 32677 17663 32735 17669
rect 32677 17629 32689 17663
rect 32723 17629 32735 17663
rect 33318 17660 33324 17672
rect 33279 17632 33324 17660
rect 32677 17623 32735 17629
rect 33318 17620 33324 17632
rect 33376 17620 33382 17672
rect 33962 17660 33968 17672
rect 33923 17632 33968 17660
rect 33962 17620 33968 17632
rect 34020 17620 34026 17672
rect 34900 17669 34928 17700
rect 34885 17663 34943 17669
rect 34885 17629 34897 17663
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 34977 17663 35035 17669
rect 34977 17629 34989 17663
rect 35023 17660 35035 17663
rect 35713 17663 35771 17669
rect 35713 17660 35725 17663
rect 35023 17632 35725 17660
rect 35023 17629 35035 17632
rect 34977 17623 35035 17629
rect 35713 17629 35725 17632
rect 35759 17629 35771 17663
rect 35713 17623 35771 17629
rect 33413 17595 33471 17601
rect 33413 17592 33425 17595
rect 32600 17564 33425 17592
rect 33413 17561 33425 17564
rect 33459 17561 33471 17595
rect 33413 17555 33471 17561
rect 33042 17524 33048 17536
rect 31680 17496 33048 17524
rect 33042 17484 33048 17496
rect 33100 17484 33106 17536
rect 33134 17484 33140 17536
rect 33192 17524 33198 17536
rect 34057 17527 34115 17533
rect 34057 17524 34069 17527
rect 33192 17496 34069 17524
rect 33192 17484 33198 17496
rect 34057 17493 34069 17496
rect 34103 17493 34115 17527
rect 34057 17487 34115 17493
rect 35529 17527 35587 17533
rect 35529 17493 35541 17527
rect 35575 17524 35587 17527
rect 37182 17524 37188 17536
rect 35575 17496 37188 17524
rect 35575 17493 35587 17496
rect 35529 17487 35587 17493
rect 37182 17484 37188 17496
rect 37240 17484 37246 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 9674 17320 9680 17332
rect 7576 17292 9680 17320
rect 7006 17252 7012 17264
rect 6967 17224 7012 17252
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 7576 17261 7604 17292
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 16850 17320 16856 17332
rect 11756 17292 13492 17320
rect 11756 17280 11762 17292
rect 7561 17255 7619 17261
rect 7561 17221 7573 17255
rect 7607 17221 7619 17255
rect 8110 17252 8116 17264
rect 8071 17224 8116 17252
rect 7561 17215 7619 17221
rect 8110 17212 8116 17224
rect 8168 17212 8174 17264
rect 8202 17212 8208 17264
rect 8260 17252 8266 17264
rect 9125 17255 9183 17261
rect 8260 17224 8305 17252
rect 8260 17212 8266 17224
rect 9125 17221 9137 17255
rect 9171 17252 9183 17255
rect 9766 17252 9772 17264
rect 9171 17224 9772 17252
rect 9171 17221 9183 17224
rect 9125 17215 9183 17221
rect 9766 17212 9772 17224
rect 9824 17252 9830 17264
rect 10502 17252 10508 17264
rect 9824 17224 10508 17252
rect 9824 17212 9830 17224
rect 10502 17212 10508 17224
rect 10560 17212 10566 17264
rect 10870 17212 10876 17264
rect 10928 17252 10934 17264
rect 11885 17255 11943 17261
rect 11885 17252 11897 17255
rect 10928 17224 11897 17252
rect 10928 17212 10934 17224
rect 11885 17221 11897 17224
rect 11931 17221 11943 17255
rect 11885 17215 11943 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 5074 17184 5080 17196
rect 1903 17156 5080 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 5074 17144 5080 17156
rect 5132 17184 5138 17196
rect 5442 17184 5448 17196
rect 5132 17156 5448 17184
rect 5132 17144 5138 17156
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 5810 17184 5816 17196
rect 5771 17156 5816 17184
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 10321 17187 10379 17193
rect 9732 17156 9777 17184
rect 9732 17144 9738 17156
rect 10321 17153 10333 17187
rect 10367 17153 10379 17187
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 10321 17147 10379 17153
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6730 17116 6736 17128
rect 5951 17088 6736 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6730 17076 6736 17088
rect 6788 17116 6794 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6788 17088 6929 17116
rect 6788 17076 6794 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 10336 17116 10364 17147
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 13464 17193 13492 17292
rect 14752 17292 16856 17320
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17153 13507 17187
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 13449 17147 13507 17153
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 11422 17116 11428 17128
rect 10336 17088 11428 17116
rect 6917 17079 6975 17085
rect 11422 17076 11428 17088
rect 11480 17076 11486 17128
rect 11790 17116 11796 17128
rect 11751 17088 11796 17116
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12492 17088 12537 17116
rect 12492 17076 12498 17088
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 14752 17116 14780 17292
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 18046 17320 18052 17332
rect 16991 17292 18052 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 27614 17320 27620 17332
rect 18156 17292 23428 17320
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 15289 17255 15347 17261
rect 15289 17252 15301 17255
rect 15252 17224 15301 17252
rect 15252 17212 15258 17224
rect 15289 17221 15301 17224
rect 15335 17221 15347 17255
rect 18156 17252 18184 17292
rect 18322 17252 18328 17264
rect 15289 17215 15347 17221
rect 16776 17224 18184 17252
rect 18283 17224 18328 17252
rect 12768 17088 14780 17116
rect 12768 17076 12774 17088
rect 14826 17076 14832 17128
rect 14884 17116 14890 17128
rect 15197 17119 15255 17125
rect 15197 17116 15209 17119
rect 14884 17088 15209 17116
rect 14884 17076 14890 17088
rect 15197 17085 15209 17088
rect 15243 17085 15255 17119
rect 15654 17116 15660 17128
rect 15615 17088 15660 17116
rect 15197 17079 15255 17085
rect 15654 17076 15660 17088
rect 15712 17116 15718 17128
rect 16776 17116 16804 17224
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 20070 17212 20076 17264
rect 20128 17252 20134 17264
rect 20128 17224 20392 17252
rect 20128 17212 20134 17224
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 16908 17156 16953 17184
rect 16908 17144 16914 17156
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 17497 17187 17555 17193
rect 17497 17184 17509 17187
rect 17092 17156 17509 17184
rect 17092 17144 17098 17156
rect 17497 17153 17509 17156
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17153 19763 17187
rect 20364 17184 20392 17224
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 20901 17255 20959 17261
rect 20901 17252 20913 17255
rect 20864 17224 20913 17252
rect 20864 17212 20870 17224
rect 20901 17221 20913 17224
rect 20947 17221 20959 17255
rect 20901 17215 20959 17221
rect 21726 17212 21732 17264
rect 21784 17252 21790 17264
rect 22281 17255 22339 17261
rect 22281 17252 22293 17255
rect 21784 17224 22293 17252
rect 21784 17212 21790 17224
rect 22281 17221 22293 17224
rect 22327 17221 22339 17255
rect 22281 17215 22339 17221
rect 22373 17255 22431 17261
rect 22373 17221 22385 17255
rect 22419 17252 22431 17255
rect 23290 17252 23296 17264
rect 22419 17224 23296 17252
rect 22419 17221 22431 17224
rect 22373 17215 22431 17221
rect 23290 17212 23296 17224
rect 23348 17212 23354 17264
rect 20438 17184 20444 17196
rect 20364 17156 20444 17184
rect 19705 17147 19763 17153
rect 15712 17088 16804 17116
rect 18233 17119 18291 17125
rect 15712 17076 15718 17088
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18414 17116 18420 17128
rect 18279 17088 18420 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 18414 17076 18420 17088
rect 18472 17076 18478 17128
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 12250 17048 12256 17060
rect 8260 17020 12256 17048
rect 8260 17008 8266 17020
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 17954 17008 17960 17060
rect 18012 17048 18018 17060
rect 18524 17048 18552 17079
rect 18012 17020 18552 17048
rect 18012 17008 18018 17020
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10410 16980 10416 16992
rect 10371 16952 10416 16980
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 13538 16980 13544 16992
rect 13499 16952 13544 16980
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 14553 16983 14611 16989
rect 14553 16949 14565 16983
rect 14599 16980 14611 16983
rect 15102 16980 15108 16992
rect 14599 16952 15108 16980
rect 14599 16949 14611 16952
rect 14553 16943 14611 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 17862 16980 17868 16992
rect 17635 16952 17868 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 19720 16980 19748 17147
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 20070 17116 20076 17128
rect 20027 17088 20076 17116
rect 20027 17085 20039 17088
rect 19981 17079 20039 17085
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20809 17119 20867 17125
rect 20809 17085 20821 17119
rect 20855 17116 20867 17119
rect 21266 17116 21272 17128
rect 20855 17088 21272 17116
rect 20855 17085 20867 17088
rect 20809 17079 20867 17085
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 23290 17116 23296 17128
rect 23251 17088 23296 17116
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 23400 17116 23428 17292
rect 24872 17292 27620 17320
rect 23934 17252 23940 17264
rect 23895 17224 23940 17252
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 24872 17261 24900 17292
rect 27614 17280 27620 17292
rect 27672 17280 27678 17332
rect 30282 17280 30288 17332
rect 30340 17320 30346 17332
rect 31665 17323 31723 17329
rect 31665 17320 31677 17323
rect 30340 17292 31677 17320
rect 30340 17280 30346 17292
rect 31665 17289 31677 17292
rect 31711 17289 31723 17323
rect 31665 17283 31723 17289
rect 32306 17280 32312 17332
rect 32364 17320 32370 17332
rect 32401 17323 32459 17329
rect 32401 17320 32413 17323
rect 32364 17292 32413 17320
rect 32364 17280 32370 17292
rect 32401 17289 32413 17292
rect 32447 17289 32459 17323
rect 33042 17320 33048 17332
rect 33003 17292 33048 17320
rect 32401 17283 32459 17289
rect 33042 17280 33048 17292
rect 33100 17280 33106 17332
rect 33689 17323 33747 17329
rect 33689 17289 33701 17323
rect 33735 17320 33747 17323
rect 35618 17320 35624 17332
rect 33735 17292 35624 17320
rect 33735 17289 33747 17292
rect 33689 17283 33747 17289
rect 35618 17280 35624 17292
rect 35676 17280 35682 17332
rect 24857 17255 24915 17261
rect 24857 17221 24869 17255
rect 24903 17221 24915 17255
rect 25498 17252 25504 17264
rect 25459 17224 25504 17252
rect 24857 17215 24915 17221
rect 25498 17212 25504 17224
rect 25556 17212 25562 17264
rect 28258 17252 28264 17264
rect 26252 17224 28264 17252
rect 23845 17119 23903 17125
rect 23845 17116 23857 17119
rect 23400 17088 23857 17116
rect 23845 17085 23857 17088
rect 23891 17085 23903 17119
rect 23845 17079 23903 17085
rect 24026 17076 24032 17128
rect 24084 17116 24090 17128
rect 25409 17119 25467 17125
rect 25409 17116 25421 17119
rect 24084 17088 25421 17116
rect 24084 17076 24090 17088
rect 25409 17085 25421 17088
rect 25455 17085 25467 17119
rect 25409 17079 25467 17085
rect 25498 17076 25504 17128
rect 25556 17116 25562 17128
rect 26252 17116 26280 17224
rect 28258 17212 28264 17224
rect 28316 17212 28322 17264
rect 28629 17255 28687 17261
rect 28629 17221 28641 17255
rect 28675 17252 28687 17255
rect 30098 17252 30104 17264
rect 28675 17224 30104 17252
rect 28675 17221 28687 17224
rect 28629 17215 28687 17221
rect 30098 17212 30104 17224
rect 30156 17212 30162 17264
rect 30193 17255 30251 17261
rect 30193 17221 30205 17255
rect 30239 17252 30251 17255
rect 31294 17252 31300 17264
rect 30239 17224 31300 17252
rect 30239 17221 30251 17224
rect 30193 17215 30251 17221
rect 31294 17212 31300 17224
rect 31352 17212 31358 17264
rect 34790 17252 34796 17264
rect 32968 17224 34796 17252
rect 32968 17196 32996 17224
rect 34790 17212 34796 17224
rect 34848 17212 34854 17264
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27798 17184 27804 17196
rect 27203 17156 27804 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 31573 17187 31631 17193
rect 31573 17184 31585 17187
rect 30944 17156 31585 17184
rect 26418 17116 26424 17128
rect 25556 17088 26280 17116
rect 26379 17088 26424 17116
rect 25556 17076 25562 17088
rect 26418 17076 26424 17088
rect 26476 17076 26482 17128
rect 27338 17116 27344 17128
rect 27299 17088 27344 17116
rect 27338 17076 27344 17088
rect 27396 17076 27402 17128
rect 27982 17076 27988 17128
rect 28040 17116 28046 17128
rect 28537 17119 28595 17125
rect 28537 17116 28549 17119
rect 28040 17088 28549 17116
rect 28040 17076 28046 17088
rect 28537 17085 28549 17088
rect 28583 17085 28595 17119
rect 29362 17116 29368 17128
rect 29323 17088 29368 17116
rect 28537 17079 28595 17085
rect 29362 17076 29368 17088
rect 29420 17076 29426 17128
rect 30101 17119 30159 17125
rect 30101 17085 30113 17119
rect 30147 17116 30159 17119
rect 30650 17116 30656 17128
rect 30147 17088 30656 17116
rect 30147 17085 30159 17088
rect 30101 17079 30159 17085
rect 30650 17076 30656 17088
rect 30708 17076 30714 17128
rect 30742 17076 30748 17128
rect 30800 17116 30806 17128
rect 30944 17116 30972 17156
rect 31573 17153 31585 17156
rect 31619 17153 31631 17187
rect 32306 17184 32312 17196
rect 32267 17156 32312 17184
rect 31573 17147 31631 17153
rect 32306 17144 32312 17156
rect 32364 17144 32370 17196
rect 32950 17184 32956 17196
rect 32911 17156 32956 17184
rect 32950 17144 32956 17156
rect 33008 17144 33014 17196
rect 33597 17187 33655 17193
rect 33597 17153 33609 17187
rect 33643 17153 33655 17187
rect 38286 17184 38292 17196
rect 38247 17156 38292 17184
rect 33597 17147 33655 17153
rect 30800 17088 30972 17116
rect 30800 17076 30806 17088
rect 31018 17076 31024 17128
rect 31076 17116 31082 17128
rect 31076 17088 31121 17116
rect 31076 17076 31082 17088
rect 20714 17008 20720 17060
rect 20772 17048 20778 17060
rect 21361 17051 21419 17057
rect 21361 17048 21373 17051
rect 20772 17020 21373 17048
rect 20772 17008 20778 17020
rect 21361 17017 21373 17020
rect 21407 17017 21419 17051
rect 33612 17048 33640 17147
rect 38286 17144 38292 17156
rect 38344 17144 38350 17196
rect 21361 17011 21419 17017
rect 22066 17020 33640 17048
rect 20806 16980 20812 16992
rect 19720 16952 20812 16980
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 21376 16980 21404 17011
rect 22066 16980 22094 17020
rect 21376 16952 22094 16980
rect 24762 16940 24768 16992
rect 24820 16980 24826 16992
rect 26418 16980 26424 16992
rect 24820 16952 26424 16980
rect 24820 16940 24826 16952
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 29362 16940 29368 16992
rect 29420 16980 29426 16992
rect 30650 16980 30656 16992
rect 29420 16952 30656 16980
rect 29420 16940 29426 16952
rect 30650 16940 30656 16952
rect 30708 16940 30714 16992
rect 38102 16980 38108 16992
rect 38063 16952 38108 16980
rect 38102 16940 38108 16952
rect 38160 16940 38166 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 12710 16776 12716 16788
rect 12308 16748 12716 16776
rect 12308 16736 12314 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 16206 16776 16212 16788
rect 13280 16748 16212 16776
rect 9398 16708 9404 16720
rect 5184 16680 9404 16708
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 5184 16572 5212 16680
rect 9398 16668 9404 16680
rect 9456 16668 9462 16720
rect 10962 16668 10968 16720
rect 11020 16708 11026 16720
rect 13280 16708 13308 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 17000 16748 18920 16776
rect 17000 16736 17006 16748
rect 11020 16680 13308 16708
rect 11020 16668 11026 16680
rect 5258 16600 5264 16652
rect 5316 16640 5322 16652
rect 7374 16640 7380 16652
rect 5316 16612 6684 16640
rect 7335 16612 7380 16640
rect 5316 16600 5322 16612
rect 6012 16581 6040 16612
rect 6656 16581 6684 16612
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8294 16640 8300 16652
rect 8251 16612 8300 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 5353 16575 5411 16581
rect 5353 16572 5365 16575
rect 1995 16544 2268 16572
rect 5184 16544 5365 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2240 16516 2268 16544
rect 5353 16541 5365 16544
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 5997 16575 6055 16581
rect 5997 16541 6009 16575
rect 6043 16541 6055 16575
rect 5997 16535 6055 16541
rect 6641 16575 6699 16581
rect 6641 16541 6653 16575
rect 6687 16541 6699 16575
rect 6641 16535 6699 16541
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16572 11023 16575
rect 11422 16572 11428 16584
rect 11011 16544 11428 16572
rect 11011 16541 11023 16544
rect 10965 16535 11023 16541
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 12158 16572 12164 16584
rect 11655 16544 12164 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12897 16575 12955 16581
rect 12308 16544 12353 16572
rect 12308 16532 12314 16544
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 13280 16572 13308 16680
rect 13446 16668 13452 16720
rect 13504 16708 13510 16720
rect 13814 16708 13820 16720
rect 13504 16680 13820 16708
rect 13504 16668 13510 16680
rect 13814 16668 13820 16680
rect 13872 16668 13878 16720
rect 16390 16668 16396 16720
rect 16448 16708 16454 16720
rect 18892 16708 18920 16748
rect 19886 16736 19892 16788
rect 19944 16776 19950 16788
rect 20530 16776 20536 16788
rect 19944 16748 20536 16776
rect 19944 16736 19950 16748
rect 20530 16736 20536 16748
rect 20588 16736 20594 16788
rect 20806 16736 20812 16788
rect 20864 16776 20870 16788
rect 23293 16779 23351 16785
rect 23293 16776 23305 16779
rect 20864 16748 23305 16776
rect 20864 16736 20870 16748
rect 23293 16745 23305 16748
rect 23339 16745 23351 16779
rect 25498 16776 25504 16788
rect 23293 16739 23351 16745
rect 24412 16748 25504 16776
rect 21726 16708 21732 16720
rect 16448 16680 18736 16708
rect 18892 16680 21732 16708
rect 16448 16668 16454 16680
rect 13722 16600 13728 16652
rect 13780 16640 13786 16652
rect 15933 16643 15991 16649
rect 15933 16640 15945 16643
rect 13780 16612 15945 16640
rect 13780 16600 13786 16612
rect 15933 16609 15945 16612
rect 15979 16609 15991 16643
rect 15933 16603 15991 16609
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 18598 16640 18604 16652
rect 16172 16612 17080 16640
rect 16172 16600 16178 16612
rect 12943 16544 13308 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13504 16544 13553 16572
rect 13504 16532 13510 16544
rect 13541 16541 13553 16544
rect 13587 16572 13599 16575
rect 14277 16575 14335 16581
rect 14277 16572 14289 16575
rect 13587 16544 14289 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 14277 16541 14289 16544
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16572 14979 16575
rect 15194 16572 15200 16584
rect 14967 16544 15200 16572
rect 14967 16541 14979 16544
rect 14921 16535 14979 16541
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 17052 16581 17080 16612
rect 18064 16612 18604 16640
rect 18064 16581 18092 16612
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 18708 16640 18736 16680
rect 21726 16668 21732 16680
rect 21784 16668 21790 16720
rect 20073 16643 20131 16649
rect 18708 16612 19334 16640
rect 19306 16584 19334 16612
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 24412 16640 24440 16748
rect 25498 16736 25504 16748
rect 25556 16736 25562 16788
rect 25590 16736 25596 16788
rect 25648 16776 25654 16788
rect 25961 16779 26019 16785
rect 25961 16776 25973 16779
rect 25648 16748 25973 16776
rect 25648 16736 25654 16748
rect 25961 16745 25973 16748
rect 26007 16745 26019 16779
rect 25961 16739 26019 16745
rect 26418 16736 26424 16788
rect 26476 16776 26482 16788
rect 30190 16776 30196 16788
rect 26476 16748 30196 16776
rect 26476 16736 26482 16748
rect 30190 16736 30196 16748
rect 30248 16736 30254 16788
rect 31662 16776 31668 16788
rect 30944 16748 31668 16776
rect 24486 16668 24492 16720
rect 24544 16708 24550 16720
rect 29454 16708 29460 16720
rect 24544 16680 26004 16708
rect 24544 16668 24550 16680
rect 20119 16612 24440 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 25976 16640 26004 16680
rect 27724 16680 29460 16708
rect 27724 16640 27752 16680
rect 29454 16668 29460 16680
rect 29512 16668 29518 16720
rect 24912 16612 25912 16640
rect 25976 16612 27752 16640
rect 24912 16600 24918 16612
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 18564 16544 18705 16572
rect 18564 16532 18570 16544
rect 18693 16541 18705 16544
rect 18739 16541 18751 16575
rect 19306 16544 19340 16584
rect 18693 16535 18751 16541
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 24578 16572 24584 16584
rect 23124 16544 23336 16572
rect 24539 16544 24584 16572
rect 2222 16464 2228 16516
rect 2280 16504 2286 16516
rect 5810 16504 5816 16516
rect 2280 16476 5816 16504
rect 2280 16464 2286 16476
rect 5810 16464 5816 16476
rect 5868 16464 5874 16516
rect 6733 16507 6791 16513
rect 6733 16473 6745 16507
rect 6779 16504 6791 16507
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 6779 16476 7481 16504
rect 6779 16473 6791 16476
rect 6733 16467 6791 16473
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 9214 16504 9220 16516
rect 9175 16476 9220 16504
rect 7469 16467 7527 16473
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16473 9367 16507
rect 10226 16504 10232 16516
rect 10187 16476 10232 16504
rect 9309 16467 9367 16473
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 1765 16439 1823 16445
rect 1765 16436 1777 16439
rect 1544 16408 1777 16436
rect 1544 16396 1550 16408
rect 1765 16405 1777 16408
rect 1811 16405 1823 16439
rect 5442 16436 5448 16448
rect 5403 16408 5448 16436
rect 1765 16399 1823 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6089 16439 6147 16445
rect 6089 16405 6101 16439
rect 6135 16436 6147 16439
rect 6914 16436 6920 16448
rect 6135 16408 6920 16436
rect 6135 16405 6147 16408
rect 6089 16399 6147 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 9030 16396 9036 16448
rect 9088 16436 9094 16448
rect 9324 16436 9352 16467
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10594 16464 10600 16516
rect 10652 16504 10658 16516
rect 15013 16507 15071 16513
rect 15013 16504 15025 16507
rect 10652 16476 15025 16504
rect 10652 16464 10658 16476
rect 15013 16473 15025 16476
rect 15059 16473 15071 16507
rect 15654 16504 15660 16516
rect 15615 16476 15660 16504
rect 15013 16467 15071 16473
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 15749 16507 15807 16513
rect 15749 16473 15761 16507
rect 15795 16473 15807 16507
rect 15749 16467 15807 16473
rect 9088 16408 9352 16436
rect 9088 16396 9094 16408
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11057 16439 11115 16445
rect 11057 16436 11069 16439
rect 11020 16408 11069 16436
rect 11020 16396 11026 16408
rect 11057 16405 11069 16408
rect 11103 16405 11115 16439
rect 11057 16399 11115 16405
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11790 16436 11796 16448
rect 11747 16408 11796 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 12345 16439 12403 16445
rect 12345 16405 12357 16439
rect 12391 16436 12403 16439
rect 12618 16436 12624 16448
rect 12391 16408 12624 16436
rect 12391 16405 12403 16408
rect 12345 16399 12403 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12768 16408 13001 16436
rect 12768 16396 12774 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13354 16436 13360 16448
rect 13136 16408 13360 16436
rect 13136 16396 13142 16408
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13630 16436 13636 16448
rect 13591 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14369 16439 14427 16445
rect 14369 16405 14381 16439
rect 14415 16436 14427 16439
rect 14918 16436 14924 16448
rect 14415 16408 14924 16436
rect 14415 16405 14427 16408
rect 14369 16399 14427 16405
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 15764 16436 15792 16467
rect 17954 16464 17960 16516
rect 18012 16504 18018 16516
rect 19886 16504 19892 16516
rect 18012 16476 19892 16504
rect 18012 16464 18018 16476
rect 19886 16464 19892 16476
rect 19944 16464 19950 16516
rect 20165 16507 20223 16513
rect 20165 16473 20177 16507
rect 20211 16504 20223 16507
rect 20211 16476 20300 16504
rect 20211 16473 20223 16476
rect 20165 16467 20223 16473
rect 20272 16448 20300 16476
rect 20530 16464 20536 16516
rect 20588 16504 20594 16516
rect 21085 16507 21143 16513
rect 21085 16504 21097 16507
rect 20588 16476 21097 16504
rect 20588 16464 20594 16476
rect 21085 16473 21097 16476
rect 21131 16473 21143 16507
rect 21085 16467 21143 16473
rect 21450 16464 21456 16516
rect 21508 16504 21514 16516
rect 21637 16507 21695 16513
rect 21637 16504 21649 16507
rect 21508 16476 21649 16504
rect 21508 16464 21514 16476
rect 21637 16473 21649 16476
rect 21683 16473 21695 16507
rect 21637 16467 21695 16473
rect 21729 16507 21787 16513
rect 21729 16473 21741 16507
rect 21775 16504 21787 16507
rect 22186 16504 22192 16516
rect 21775 16476 22192 16504
rect 21775 16473 21787 16476
rect 21729 16467 21787 16473
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 22649 16507 22707 16513
rect 22649 16473 22661 16507
rect 22695 16504 22707 16507
rect 23014 16504 23020 16516
rect 22695 16476 23020 16504
rect 22695 16473 22707 16476
rect 22649 16467 22707 16473
rect 23014 16464 23020 16476
rect 23072 16464 23078 16516
rect 15160 16408 15792 16436
rect 17129 16439 17187 16445
rect 15160 16396 15166 16408
rect 17129 16405 17141 16439
rect 17175 16436 17187 16439
rect 17310 16436 17316 16448
rect 17175 16408 17316 16436
rect 17175 16405 17187 16408
rect 17129 16399 17187 16405
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 18138 16436 18144 16448
rect 18099 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 18785 16439 18843 16445
rect 18785 16405 18797 16439
rect 18831 16436 18843 16439
rect 19426 16436 19432 16448
rect 18831 16408 19432 16436
rect 18831 16405 18843 16408
rect 18785 16399 18843 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 20254 16396 20260 16448
rect 20312 16396 20318 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 23124 16436 23152 16544
rect 23201 16507 23259 16513
rect 23201 16473 23213 16507
rect 23247 16473 23259 16507
rect 23308 16504 23336 16544
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 23308 16476 24685 16504
rect 23201 16467 23259 16473
rect 24673 16473 24685 16476
rect 24719 16473 24731 16507
rect 25240 16504 25268 16535
rect 25314 16532 25320 16584
rect 25372 16572 25378 16584
rect 25884 16581 25912 16612
rect 27798 16600 27804 16652
rect 27856 16640 27862 16652
rect 27856 16612 28488 16640
rect 27856 16600 27862 16612
rect 28460 16581 28488 16612
rect 28718 16600 28724 16652
rect 28776 16640 28782 16652
rect 30944 16649 30972 16748
rect 31662 16736 31668 16748
rect 31720 16776 31726 16788
rect 34698 16776 34704 16788
rect 31720 16748 34704 16776
rect 31720 16736 31726 16748
rect 34698 16736 34704 16748
rect 34756 16736 34762 16788
rect 31018 16668 31024 16720
rect 31076 16708 31082 16720
rect 32674 16708 32680 16720
rect 31076 16680 32680 16708
rect 31076 16668 31082 16680
rect 32674 16668 32680 16680
rect 32732 16668 32738 16720
rect 37550 16708 37556 16720
rect 33980 16680 37556 16708
rect 30929 16643 30987 16649
rect 28776 16612 29776 16640
rect 28776 16600 28782 16612
rect 25869 16575 25927 16581
rect 25372 16544 25417 16572
rect 25372 16532 25378 16544
rect 25869 16541 25881 16575
rect 25915 16541 25927 16575
rect 25869 16535 25927 16541
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16572 28503 16575
rect 28626 16572 28632 16584
rect 28491 16544 28632 16572
rect 28491 16541 28503 16544
rect 28445 16535 28503 16541
rect 28626 16532 28632 16544
rect 28684 16532 28690 16584
rect 29748 16581 29776 16612
rect 30929 16609 30941 16643
rect 30975 16609 30987 16643
rect 30929 16603 30987 16609
rect 31754 16600 31760 16652
rect 31812 16640 31818 16652
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 31812 16612 32505 16640
rect 31812 16600 31818 16612
rect 32493 16609 32505 16612
rect 32539 16609 32551 16643
rect 32493 16603 32551 16609
rect 33980 16581 34008 16680
rect 37550 16668 37556 16680
rect 37608 16668 37614 16720
rect 38102 16640 38108 16652
rect 34900 16612 38108 16640
rect 34900 16581 34928 16612
rect 38102 16600 38108 16612
rect 38160 16600 38166 16652
rect 29733 16575 29791 16581
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 33965 16575 34023 16581
rect 33965 16541 33977 16575
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 25682 16504 25688 16516
rect 25240 16476 25688 16504
rect 24673 16467 24731 16473
rect 20956 16408 23152 16436
rect 23216 16436 23244 16467
rect 25682 16464 25688 16476
rect 25740 16464 25746 16516
rect 26973 16507 27031 16513
rect 26973 16473 26985 16507
rect 27019 16473 27031 16507
rect 26973 16467 27031 16473
rect 27065 16507 27123 16513
rect 27065 16473 27077 16507
rect 27111 16504 27123 16507
rect 27798 16504 27804 16516
rect 27111 16476 27804 16504
rect 27111 16473 27123 16476
rect 27065 16467 27123 16473
rect 23290 16436 23296 16448
rect 23216 16408 23296 16436
rect 20956 16396 20962 16408
rect 23290 16396 23296 16408
rect 23348 16396 23354 16448
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 25498 16436 25504 16448
rect 23440 16408 25504 16436
rect 23440 16396 23446 16408
rect 25498 16396 25504 16408
rect 25556 16396 25562 16448
rect 26988 16436 27016 16467
rect 27798 16464 27804 16476
rect 27856 16464 27862 16516
rect 27985 16507 28043 16513
rect 27985 16473 27997 16507
rect 28031 16504 28043 16507
rect 28258 16504 28264 16516
rect 28031 16476 28264 16504
rect 28031 16473 28043 16476
rect 27985 16467 28043 16473
rect 28258 16464 28264 16476
rect 28316 16464 28322 16516
rect 28721 16507 28779 16513
rect 28721 16473 28733 16507
rect 28767 16504 28779 16507
rect 28810 16504 28816 16516
rect 28767 16476 28816 16504
rect 28767 16473 28779 16476
rect 28721 16467 28779 16473
rect 28810 16464 28816 16476
rect 28868 16464 28874 16516
rect 29638 16464 29644 16516
rect 29696 16504 29702 16516
rect 29825 16507 29883 16513
rect 29825 16504 29837 16507
rect 29696 16476 29837 16504
rect 29696 16464 29702 16476
rect 29825 16473 29837 16476
rect 29871 16473 29883 16507
rect 29825 16467 29883 16473
rect 30006 16464 30012 16516
rect 30064 16504 30070 16516
rect 30926 16504 30932 16516
rect 30064 16476 30932 16504
rect 30064 16464 30070 16476
rect 30926 16464 30932 16476
rect 30984 16464 30990 16516
rect 31021 16507 31079 16513
rect 31021 16473 31033 16507
rect 31067 16504 31079 16507
rect 31386 16504 31392 16516
rect 31067 16476 31392 16504
rect 31067 16473 31079 16476
rect 31021 16467 31079 16473
rect 31386 16464 31392 16476
rect 31444 16464 31450 16516
rect 31846 16464 31852 16516
rect 31904 16504 31910 16516
rect 31941 16507 31999 16513
rect 31941 16504 31953 16507
rect 31904 16476 31953 16504
rect 31904 16464 31910 16476
rect 31941 16473 31953 16476
rect 31987 16473 31999 16507
rect 31941 16467 31999 16473
rect 32582 16464 32588 16516
rect 32640 16504 32646 16516
rect 33502 16504 33508 16516
rect 32640 16476 32685 16504
rect 33463 16476 33508 16504
rect 32640 16464 32646 16476
rect 33502 16464 33508 16476
rect 33560 16464 33566 16516
rect 34977 16507 35035 16513
rect 34977 16504 34989 16507
rect 33612 16476 34989 16504
rect 27154 16436 27160 16448
rect 26988 16408 27160 16436
rect 27154 16396 27160 16408
rect 27212 16396 27218 16448
rect 27246 16396 27252 16448
rect 27304 16436 27310 16448
rect 33612 16436 33640 16476
rect 34977 16473 34989 16476
rect 35023 16473 35035 16507
rect 34977 16467 35035 16473
rect 34054 16436 34060 16448
rect 27304 16408 33640 16436
rect 34015 16408 34060 16436
rect 27304 16396 27310 16408
rect 34054 16396 34060 16408
rect 34112 16396 34118 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 8478 16232 8484 16244
rect 2746 16204 8484 16232
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 1596 15960 1624 16059
rect 2746 15960 2774 16204
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 13630 16232 13636 16244
rect 10376 16204 13636 16232
rect 10376 16192 10382 16204
rect 13630 16192 13636 16204
rect 13688 16192 13694 16244
rect 14274 16192 14280 16244
rect 14332 16232 14338 16244
rect 15654 16232 15660 16244
rect 14332 16204 15660 16232
rect 14332 16192 14338 16204
rect 15654 16192 15660 16204
rect 15712 16232 15718 16244
rect 24118 16232 24124 16244
rect 15712 16204 23428 16232
rect 24079 16204 24124 16232
rect 15712 16192 15718 16204
rect 6822 16164 6828 16176
rect 6783 16136 6828 16164
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 8386 16164 8392 16176
rect 8347 16136 8392 16164
rect 8386 16124 8392 16136
rect 8444 16124 8450 16176
rect 10226 16164 10232 16176
rect 10187 16136 10232 16164
rect 10226 16124 10232 16136
rect 10284 16124 10290 16176
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 10836 16136 11805 16164
rect 10836 16124 10842 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 11885 16167 11943 16173
rect 11885 16133 11897 16167
rect 11931 16164 11943 16167
rect 12066 16164 12072 16176
rect 11931 16136 12072 16164
rect 11931 16133 11943 16136
rect 11885 16127 11943 16133
rect 12066 16124 12072 16136
rect 12124 16124 12130 16176
rect 12802 16164 12808 16176
rect 12763 16136 12808 16164
rect 12802 16124 12808 16136
rect 12860 16124 12866 16176
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 14369 16167 14427 16173
rect 14369 16164 14381 16167
rect 13596 16136 14381 16164
rect 13596 16124 13602 16136
rect 14369 16133 14381 16136
rect 14415 16133 14427 16167
rect 14369 16127 14427 16133
rect 15856 16136 16712 16164
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 5859 16000 6745 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7009 15991 7067 15997
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 16028 8355 16031
rect 8570 16028 8576 16040
rect 8343 16000 8576 16028
rect 8343 15997 8355 16000
rect 8297 15991 8355 15997
rect 1596 15932 2774 15960
rect 7024 15904 7052 15991
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 10134 16028 10140 16040
rect 8720 16000 8765 16028
rect 10095 16000 10140 16028
rect 8720 15988 8726 16000
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10560 16000 11161 16028
rect 10560 15988 10566 16000
rect 11149 15997 11161 16000
rect 11195 16028 11207 16031
rect 12820 16028 12848 16124
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13449 16099 13507 16105
rect 13449 16096 13461 16099
rect 13044 16068 13461 16096
rect 13044 16056 13050 16068
rect 13449 16065 13461 16068
rect 13495 16096 13507 16099
rect 13630 16096 13636 16108
rect 13495 16068 13636 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14274 16028 14280 16040
rect 11195 16000 12848 16028
rect 14235 16000 14280 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 14550 16028 14556 16040
rect 14511 16000 14556 16028
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 8680 15960 8708 15988
rect 15856 15960 15884 16136
rect 16117 16097 16175 16103
rect 16117 16063 16129 16097
rect 16163 16063 16175 16097
rect 16117 16057 16175 16063
rect 16022 15988 16028 16040
rect 16080 16028 16086 16040
rect 16132 16028 16160 16057
rect 16206 16028 16212 16040
rect 16080 16000 16212 16028
rect 16080 15988 16086 16000
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16684 16028 16712 16136
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 16816 16136 17141 16164
rect 16816 16124 16822 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 17221 16167 17279 16173
rect 17221 16133 17233 16167
rect 17267 16164 17279 16167
rect 17310 16164 17316 16176
rect 17267 16136 17316 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 18138 16124 18144 16176
rect 18196 16164 18202 16176
rect 18877 16167 18935 16173
rect 18877 16164 18889 16167
rect 18196 16136 18889 16164
rect 18196 16124 18202 16136
rect 18877 16133 18889 16136
rect 18923 16133 18935 16167
rect 18877 16127 18935 16133
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 20162 16164 20168 16176
rect 19392 16136 20168 16164
rect 19392 16124 19398 16136
rect 20162 16124 20168 16136
rect 20220 16164 20226 16176
rect 22002 16164 22008 16176
rect 20220 16136 22008 16164
rect 20220 16124 20226 16136
rect 22002 16124 22008 16136
rect 22060 16164 22066 16176
rect 22462 16164 22468 16176
rect 22060 16136 22324 16164
rect 22423 16136 22468 16164
rect 22060 16124 22066 16136
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16096 20315 16099
rect 20530 16096 20536 16108
rect 20303 16068 20536 16096
rect 20303 16065 20315 16068
rect 20257 16059 20315 16065
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 22186 16096 22192 16108
rect 21315 16068 22192 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 17954 16028 17960 16040
rect 16684 16000 16988 16028
rect 17915 16000 17960 16028
rect 16960 15960 16988 16000
rect 17954 15988 17960 16000
rect 18012 15988 18018 16040
rect 18782 16028 18788 16040
rect 18743 16000 18788 16028
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 19061 16031 19119 16037
rect 19061 15997 19073 16031
rect 19107 16028 19119 16031
rect 22296 16028 22324 16136
rect 22462 16124 22468 16136
rect 22520 16124 22526 16176
rect 22554 16124 22560 16176
rect 22612 16164 22618 16176
rect 22612 16136 22657 16164
rect 22612 16124 22618 16136
rect 19107 16000 19141 16028
rect 22296 16000 23244 16028
rect 19107 15997 19119 16000
rect 19061 15991 19119 15997
rect 19076 15960 19104 15991
rect 23106 15960 23112 15972
rect 8680 15932 15884 15960
rect 16040 15932 16896 15960
rect 16960 15932 23112 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 7006 15892 7012 15904
rect 5224 15864 7012 15892
rect 5224 15852 5230 15864
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 12860 15864 13553 15892
rect 12860 15852 12866 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 16040 15892 16068 15932
rect 16868 15904 16896 15932
rect 23106 15920 23112 15932
rect 23164 15920 23170 15972
rect 13688 15864 16068 15892
rect 16209 15895 16267 15901
rect 13688 15852 13694 15864
rect 16209 15861 16221 15895
rect 16255 15892 16267 15895
rect 16758 15892 16764 15904
rect 16255 15864 16764 15892
rect 16255 15861 16267 15864
rect 16209 15855 16267 15861
rect 16758 15852 16764 15864
rect 16816 15852 16822 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 19610 15892 19616 15904
rect 16908 15864 19616 15892
rect 16908 15852 16914 15864
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 20312 15864 20361 15892
rect 20312 15852 20318 15864
rect 20349 15861 20361 15864
rect 20395 15861 20407 15895
rect 20349 15855 20407 15861
rect 21361 15895 21419 15901
rect 21361 15861 21373 15895
rect 21407 15892 21419 15895
rect 21818 15892 21824 15904
rect 21407 15864 21824 15892
rect 21407 15861 21419 15864
rect 21361 15855 21419 15861
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 23216 15892 23244 16000
rect 23400 15960 23428 16204
rect 24118 16192 24124 16204
rect 24176 16192 24182 16244
rect 27706 16232 27712 16244
rect 25976 16204 27712 16232
rect 23474 16124 23480 16176
rect 23532 16164 23538 16176
rect 24765 16167 24823 16173
rect 24765 16164 24777 16167
rect 23532 16136 24777 16164
rect 23532 16124 23538 16136
rect 24765 16133 24777 16136
rect 24811 16133 24823 16167
rect 24765 16127 24823 16133
rect 24026 16096 24032 16108
rect 23987 16068 24032 16096
rect 24026 16056 24032 16068
rect 24084 16056 24090 16108
rect 24670 16096 24676 16108
rect 24631 16068 24676 16096
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 24946 16056 24952 16108
rect 25004 16096 25010 16108
rect 25976 16105 26004 16204
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 28092 16204 29960 16232
rect 27341 16167 27399 16173
rect 27341 16133 27353 16167
rect 27387 16164 27399 16167
rect 27890 16164 27896 16176
rect 27387 16136 27896 16164
rect 27387 16133 27399 16136
rect 27341 16127 27399 16133
rect 27890 16124 27896 16136
rect 27948 16124 27954 16176
rect 25317 16099 25375 16105
rect 25317 16096 25329 16099
rect 25004 16068 25329 16096
rect 25004 16056 25010 16068
rect 25317 16065 25329 16068
rect 25363 16065 25375 16099
rect 25317 16059 25375 16065
rect 25961 16099 26019 16105
rect 25961 16065 25973 16099
rect 26007 16065 26019 16099
rect 25961 16059 26019 16065
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 23532 16000 23577 16028
rect 23532 15988 23538 16000
rect 26142 15988 26148 16040
rect 26200 16028 26206 16040
rect 26237 16031 26295 16037
rect 26237 16028 26249 16031
rect 26200 16000 26249 16028
rect 26200 15988 26206 16000
rect 26237 15997 26249 16000
rect 26283 15997 26295 16031
rect 27246 16028 27252 16040
rect 27159 16000 27252 16028
rect 26237 15991 26295 15997
rect 27246 15988 27252 16000
rect 27304 15988 27310 16040
rect 28092 16028 28120 16204
rect 29546 16124 29552 16176
rect 29604 16164 29610 16176
rect 29932 16164 29960 16204
rect 30098 16192 30104 16244
rect 30156 16232 30162 16244
rect 31021 16235 31079 16241
rect 31021 16232 31033 16235
rect 30156 16204 31033 16232
rect 30156 16192 30162 16204
rect 31021 16201 31033 16204
rect 31067 16201 31079 16235
rect 31021 16195 31079 16201
rect 31294 16192 31300 16244
rect 31352 16232 31358 16244
rect 31665 16235 31723 16241
rect 31665 16232 31677 16235
rect 31352 16204 31677 16232
rect 31352 16192 31358 16204
rect 31665 16201 31677 16204
rect 31711 16201 31723 16235
rect 31665 16195 31723 16201
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 34054 16232 34060 16244
rect 31812 16204 34060 16232
rect 31812 16192 31818 16204
rect 34054 16192 34060 16204
rect 34112 16192 34118 16244
rect 30834 16164 30840 16176
rect 29604 16136 29776 16164
rect 29932 16136 30840 16164
rect 29604 16124 29610 16136
rect 28626 16056 28632 16108
rect 28684 16096 28690 16108
rect 28721 16099 28779 16105
rect 28721 16096 28733 16099
rect 28684 16068 28733 16096
rect 28684 16056 28690 16068
rect 28721 16065 28733 16068
rect 28767 16065 28779 16099
rect 29638 16096 29644 16108
rect 29599 16068 29644 16096
rect 28721 16059 28779 16065
rect 29638 16056 29644 16068
rect 29696 16056 29702 16108
rect 29748 16096 29776 16136
rect 30834 16124 30840 16136
rect 30892 16124 30898 16176
rect 32493 16167 32551 16173
rect 32493 16164 32505 16167
rect 31680 16136 32505 16164
rect 31680 16108 31708 16136
rect 32493 16133 32505 16136
rect 32539 16133 32551 16167
rect 32493 16127 32551 16133
rect 30285 16099 30343 16105
rect 30285 16096 30297 16099
rect 29748 16068 30297 16096
rect 30285 16065 30297 16068
rect 30331 16065 30343 16099
rect 30285 16059 30343 16065
rect 30558 16056 30564 16108
rect 30616 16096 30622 16108
rect 30929 16099 30987 16105
rect 30929 16096 30941 16099
rect 30616 16068 30941 16096
rect 30616 16056 30622 16068
rect 30929 16065 30941 16068
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 31110 16056 31116 16108
rect 31168 16096 31174 16108
rect 31573 16099 31631 16105
rect 31573 16096 31585 16099
rect 31168 16068 31585 16096
rect 31168 16056 31174 16068
rect 31573 16065 31585 16068
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 31662 16056 31668 16108
rect 31720 16056 31726 16108
rect 37182 16056 37188 16108
rect 37240 16096 37246 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 37240 16068 38025 16096
rect 37240 16056 37246 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 27356 16000 28120 16028
rect 28261 16031 28319 16037
rect 27264 15960 27292 15988
rect 23400 15932 27292 15960
rect 24854 15892 24860 15904
rect 23216 15864 24860 15892
rect 24854 15852 24860 15864
rect 24912 15852 24918 15904
rect 25222 15852 25228 15904
rect 25280 15892 25286 15904
rect 25409 15895 25467 15901
rect 25409 15892 25421 15895
rect 25280 15864 25421 15892
rect 25280 15852 25286 15864
rect 25409 15861 25421 15864
rect 25455 15861 25467 15895
rect 25409 15855 25467 15861
rect 25498 15852 25504 15904
rect 25556 15892 25562 15904
rect 27356 15892 27384 16000
rect 28261 15997 28273 16031
rect 28307 16028 28319 16031
rect 28350 16028 28356 16040
rect 28307 16000 28356 16028
rect 28307 15997 28319 16000
rect 28261 15991 28319 15997
rect 28350 15988 28356 16000
rect 28408 15988 28414 16040
rect 28997 16031 29055 16037
rect 28997 15997 29009 16031
rect 29043 16028 29055 16031
rect 29043 16000 30604 16028
rect 29043 15997 29055 16000
rect 28997 15991 29055 15997
rect 30576 15972 30604 16000
rect 31938 15988 31944 16040
rect 31996 16028 32002 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 31996 16000 32413 16028
rect 31996 15988 32002 16000
rect 32401 15997 32413 16000
rect 32447 15997 32459 16031
rect 32401 15991 32459 15997
rect 33413 16031 33471 16037
rect 33413 15997 33425 16031
rect 33459 16028 33471 16031
rect 33502 16028 33508 16040
rect 33459 16000 33508 16028
rect 33459 15997 33471 16000
rect 33413 15991 33471 15997
rect 33502 15988 33508 16000
rect 33560 16028 33566 16040
rect 34514 16028 34520 16040
rect 33560 16000 34520 16028
rect 33560 15988 33566 16000
rect 34514 15988 34520 16000
rect 34572 15988 34578 16040
rect 27890 15920 27896 15972
rect 27948 15960 27954 15972
rect 30377 15963 30435 15969
rect 30377 15960 30389 15963
rect 27948 15932 30389 15960
rect 27948 15920 27954 15932
rect 30377 15929 30389 15932
rect 30423 15929 30435 15963
rect 30377 15923 30435 15929
rect 30558 15920 30564 15972
rect 30616 15920 30622 15972
rect 31386 15920 31392 15972
rect 31444 15960 31450 15972
rect 33134 15960 33140 15972
rect 31444 15932 33140 15960
rect 31444 15920 31450 15932
rect 33134 15920 33140 15932
rect 33192 15920 33198 15972
rect 25556 15864 27384 15892
rect 25556 15852 25562 15864
rect 27982 15852 27988 15904
rect 28040 15892 28046 15904
rect 29733 15895 29791 15901
rect 29733 15892 29745 15895
rect 28040 15864 29745 15892
rect 28040 15852 28046 15864
rect 29733 15861 29745 15864
rect 29779 15861 29791 15895
rect 29733 15855 29791 15861
rect 30650 15852 30656 15904
rect 30708 15892 30714 15904
rect 31754 15892 31760 15904
rect 30708 15864 31760 15892
rect 30708 15852 30714 15864
rect 31754 15852 31760 15864
rect 31812 15852 31818 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 9030 15688 9036 15700
rect 8352 15660 9036 15688
rect 8352 15648 8358 15660
rect 9030 15648 9036 15660
rect 9088 15688 9094 15700
rect 14550 15688 14556 15700
rect 9088 15660 14556 15688
rect 9088 15648 9094 15660
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 14918 15648 14924 15700
rect 14976 15688 14982 15700
rect 17678 15688 17684 15700
rect 14976 15660 17684 15688
rect 14976 15648 14982 15660
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 20070 15688 20076 15700
rect 17828 15660 20076 15688
rect 17828 15648 17834 15660
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 23106 15688 23112 15700
rect 21100 15660 23112 15688
rect 7006 15580 7012 15632
rect 7064 15620 7070 15632
rect 17954 15620 17960 15632
rect 7064 15592 17960 15620
rect 7064 15580 7070 15592
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 20714 15620 20720 15632
rect 18064 15592 20720 15620
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 7285 15555 7343 15561
rect 7285 15552 7297 15555
rect 6788 15524 7297 15552
rect 6788 15512 6794 15524
rect 7285 15521 7297 15524
rect 7331 15521 7343 15555
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 7285 15515 7343 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 9214 15512 9220 15564
rect 9272 15552 9278 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9272 15524 9689 15552
rect 9272 15512 9278 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9950 15552 9956 15564
rect 9911 15524 9956 15552
rect 9677 15515 9735 15521
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12989 15555 13047 15561
rect 12216 15524 12940 15552
rect 12216 15512 12222 15524
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 5040 15456 5181 15484
rect 5040 15444 5046 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 12250 15484 12256 15496
rect 11655 15456 12256 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 12250 15444 12256 15456
rect 12308 15484 12314 15496
rect 12434 15484 12440 15496
rect 12308 15456 12440 15484
rect 12308 15444 12314 15456
rect 12434 15444 12440 15456
rect 12492 15444 12498 15496
rect 12912 15493 12940 15524
rect 12989 15521 13001 15555
rect 13035 15552 13047 15555
rect 14274 15552 14280 15564
rect 13035 15524 14280 15552
rect 13035 15521 13047 15524
rect 12989 15515 13047 15521
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 15194 15552 15200 15564
rect 14844 15524 15200 15552
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 1670 15416 1676 15428
rect 1631 15388 1676 15416
rect 1670 15376 1676 15388
rect 1728 15376 1734 15428
rect 1854 15416 1860 15428
rect 1815 15388 1860 15416
rect 1854 15376 1860 15388
rect 1912 15376 1918 15428
rect 5261 15419 5319 15425
rect 5261 15385 5273 15419
rect 5307 15416 5319 15419
rect 5902 15416 5908 15428
rect 5307 15388 5908 15416
rect 5307 15385 5319 15388
rect 5261 15379 5319 15385
rect 5902 15376 5908 15388
rect 5960 15376 5966 15428
rect 5997 15419 6055 15425
rect 5997 15385 6009 15419
rect 6043 15385 6055 15419
rect 5997 15379 6055 15385
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 7006 15416 7012 15428
rect 6595 15388 7012 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 6012 15348 6040 15379
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 7432 15388 7477 15416
rect 7432 15376 7438 15388
rect 9766 15376 9772 15428
rect 9824 15416 9830 15428
rect 12912 15416 12940 15447
rect 13446 15444 13452 15496
rect 13504 15484 13510 15496
rect 14844 15493 14872 15524
rect 15194 15512 15200 15524
rect 15252 15552 15258 15564
rect 17770 15552 17776 15564
rect 15252 15524 17776 15552
rect 15252 15512 15258 15524
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 18064 15552 18092 15592
rect 17972 15524 18092 15552
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13504 15456 13553 15484
rect 13504 15444 13510 15456
rect 13541 15453 13553 15456
rect 13587 15484 13599 15487
rect 14829 15487 14887 15493
rect 13587 15456 14780 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14366 15416 14372 15428
rect 9824 15388 9869 15416
rect 12912 15388 14372 15416
rect 9824 15376 9830 15388
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 14752 15416 14780 15456
rect 14829 15453 14841 15487
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15484 15531 15487
rect 15838 15484 15844 15496
rect 15519 15456 15844 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15484 16175 15487
rect 16390 15484 16396 15496
rect 16163 15456 16396 15484
rect 16163 15453 16175 15456
rect 16117 15447 16175 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 16850 15484 16856 15496
rect 16807 15456 16856 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 17972 15484 18000 15524
rect 17451 15456 18000 15484
rect 18049 15487 18107 15493
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 18414 15484 18420 15496
rect 18095 15456 18420 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 15378 15416 15384 15428
rect 14752 15388 15384 15416
rect 15378 15376 15384 15388
rect 15436 15416 15442 15428
rect 17420 15416 17448 15447
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18524 15486 18552 15592
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 18966 15552 18972 15564
rect 18831 15524 18972 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 21100 15561 21128 15660
rect 23106 15648 23112 15660
rect 23164 15688 23170 15700
rect 25130 15688 25136 15700
rect 23164 15660 25136 15688
rect 23164 15648 23170 15660
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 25314 15648 25320 15700
rect 25372 15688 25378 15700
rect 26326 15688 26332 15700
rect 25372 15660 26332 15688
rect 25372 15648 25378 15660
rect 26326 15648 26332 15660
rect 26384 15648 26390 15700
rect 26881 15691 26939 15697
rect 26881 15657 26893 15691
rect 26927 15688 26939 15691
rect 27430 15688 27436 15700
rect 26927 15660 27436 15688
rect 26927 15657 26939 15660
rect 26881 15651 26939 15657
rect 27430 15648 27436 15660
rect 27488 15648 27494 15700
rect 28074 15648 28080 15700
rect 28132 15688 28138 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 28132 15660 29837 15688
rect 28132 15648 28138 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 30466 15688 30472 15700
rect 30427 15660 30472 15688
rect 29825 15651 29883 15657
rect 30466 15648 30472 15660
rect 30524 15648 30530 15700
rect 31757 15691 31815 15697
rect 31757 15657 31769 15691
rect 31803 15688 31815 15691
rect 32582 15688 32588 15700
rect 31803 15660 32588 15688
rect 31803 15657 31815 15660
rect 31757 15651 31815 15657
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 22554 15580 22560 15632
rect 22612 15620 22618 15632
rect 23014 15620 23020 15632
rect 22612 15592 23020 15620
rect 22612 15580 22618 15592
rect 23014 15580 23020 15592
rect 23072 15620 23078 15632
rect 25406 15620 25412 15632
rect 23072 15592 25412 15620
rect 23072 15580 23078 15592
rect 25406 15580 25412 15592
rect 25464 15580 25470 15632
rect 26142 15580 26148 15632
rect 26200 15620 26206 15632
rect 32766 15620 32772 15632
rect 26200 15592 32772 15620
rect 26200 15580 26206 15592
rect 32766 15580 32772 15592
rect 32824 15580 32830 15632
rect 21085 15555 21143 15561
rect 21085 15552 21097 15555
rect 19306 15524 21097 15552
rect 18685 15487 18743 15493
rect 18524 15484 18644 15486
rect 18685 15484 18697 15487
rect 18524 15458 18697 15484
rect 18616 15456 18697 15458
rect 18685 15453 18697 15456
rect 18731 15453 18743 15487
rect 18685 15447 18743 15453
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19306 15484 19334 15524
rect 21085 15521 21097 15524
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 22278 15512 22284 15564
rect 22336 15552 22342 15564
rect 22925 15555 22983 15561
rect 22925 15552 22937 15555
rect 22336 15524 22937 15552
rect 22336 15512 22342 15524
rect 22925 15521 22937 15524
rect 22971 15521 22983 15555
rect 23290 15552 23296 15564
rect 22925 15515 22983 15521
rect 23032 15524 23296 15552
rect 19610 15484 19616 15496
rect 18932 15456 19334 15484
rect 19523 15456 19616 15484
rect 18932 15444 18938 15456
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 20070 15444 20076 15496
rect 20128 15484 20134 15496
rect 20257 15487 20315 15493
rect 20257 15484 20269 15487
rect 20128 15456 20269 15484
rect 20128 15444 20134 15456
rect 20257 15453 20269 15456
rect 20303 15484 20315 15487
rect 20303 15456 20668 15484
rect 20303 15453 20315 15456
rect 20257 15447 20315 15453
rect 15436 15388 17448 15416
rect 17497 15419 17555 15425
rect 15436 15376 15442 15388
rect 17497 15385 17509 15419
rect 17543 15416 17555 15419
rect 19334 15416 19340 15428
rect 17543 15388 18644 15416
rect 17543 15385 17555 15388
rect 17497 15379 17555 15385
rect 5500 15320 6040 15348
rect 11701 15351 11759 15357
rect 5500 15308 5506 15320
rect 11701 15317 11713 15351
rect 11747 15348 11759 15351
rect 12066 15348 12072 15360
rect 11747 15320 12072 15348
rect 11747 15317 11759 15320
rect 11701 15311 11759 15317
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 12250 15308 12256 15360
rect 12308 15348 12314 15360
rect 12345 15351 12403 15357
rect 12345 15348 12357 15351
rect 12308 15320 12357 15348
rect 12308 15308 12314 15320
rect 12345 15317 12357 15320
rect 12391 15317 12403 15351
rect 12345 15311 12403 15317
rect 13633 15351 13691 15357
rect 13633 15317 13645 15351
rect 13679 15348 13691 15351
rect 13814 15348 13820 15360
rect 13679 15320 13820 15348
rect 13679 15317 13691 15320
rect 13633 15311 13691 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14921 15351 14979 15357
rect 14921 15317 14933 15351
rect 14967 15348 14979 15351
rect 15010 15348 15016 15360
rect 14967 15320 15016 15348
rect 14967 15317 14979 15320
rect 14921 15311 14979 15317
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15562 15348 15568 15360
rect 15523 15320 15568 15348
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 16206 15348 16212 15360
rect 16167 15320 16212 15348
rect 16206 15308 16212 15320
rect 16264 15308 16270 15360
rect 16853 15351 16911 15357
rect 16853 15317 16865 15351
rect 16899 15348 16911 15351
rect 17310 15348 17316 15360
rect 16899 15320 17316 15348
rect 16899 15317 16911 15320
rect 16853 15311 16911 15317
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 18138 15348 18144 15360
rect 18099 15320 18144 15348
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 18616 15348 18644 15388
rect 18800 15388 19340 15416
rect 18800 15348 18828 15388
rect 19334 15376 19340 15388
rect 19392 15376 19398 15428
rect 19628 15416 19656 15444
rect 20162 15416 20168 15428
rect 19628 15388 20168 15416
rect 20162 15376 20168 15388
rect 20220 15376 20226 15428
rect 18616 15320 18828 15348
rect 19705 15351 19763 15357
rect 19705 15317 19717 15351
rect 19751 15348 19763 15351
rect 20070 15348 20076 15360
rect 19751 15320 20076 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 20346 15348 20352 15360
rect 20307 15320 20352 15348
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 20640 15348 20668 15456
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 20864 15456 20913 15484
rect 20864 15444 20870 15456
rect 20901 15453 20913 15456
rect 20947 15484 20959 15487
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 20947 15456 21833 15484
rect 20947 15453 20959 15456
rect 20901 15447 20959 15453
rect 21821 15453 21833 15456
rect 21867 15453 21879 15487
rect 22097 15487 22155 15493
rect 22097 15484 22109 15487
rect 21821 15447 21879 15453
rect 22020 15456 22109 15484
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 22020 15416 22048 15456
rect 22097 15453 22109 15456
rect 22143 15453 22155 15487
rect 22097 15447 22155 15453
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15484 22799 15487
rect 23032 15484 23060 15524
rect 23290 15512 23296 15524
rect 23348 15552 23354 15564
rect 24854 15552 24860 15564
rect 23348 15524 24624 15552
rect 24815 15524 24860 15552
rect 23348 15512 23354 15524
rect 23658 15484 23664 15496
rect 22787 15456 23060 15484
rect 23619 15456 23664 15484
rect 22787 15453 22799 15456
rect 22741 15447 22799 15453
rect 20772 15388 22048 15416
rect 22112 15416 22140 15447
rect 23658 15444 23664 15456
rect 23716 15484 23722 15496
rect 24394 15484 24400 15496
rect 23716 15456 24400 15484
rect 23716 15444 23722 15456
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 24596 15493 24624 15524
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 25056 15524 27476 15552
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 25056 15484 25084 15524
rect 27448 15496 27476 15524
rect 27614 15512 27620 15564
rect 27672 15552 27678 15564
rect 27672 15524 30420 15552
rect 27672 15512 27678 15524
rect 24627 15456 25084 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 25130 15444 25136 15496
rect 25188 15484 25194 15496
rect 25501 15487 25559 15493
rect 25501 15484 25513 15487
rect 25188 15456 25513 15484
rect 25188 15444 25194 15456
rect 25501 15453 25513 15456
rect 25547 15484 25559 15487
rect 26145 15487 26203 15493
rect 26145 15484 26157 15487
rect 25547 15456 26157 15484
rect 25547 15453 25559 15456
rect 25501 15447 25559 15453
rect 26145 15453 26157 15456
rect 26191 15484 26203 15487
rect 26510 15484 26516 15496
rect 26191 15456 26516 15484
rect 26191 15453 26203 15456
rect 26145 15447 26203 15453
rect 26510 15444 26516 15456
rect 26568 15444 26574 15496
rect 26602 15444 26608 15496
rect 26660 15484 26666 15496
rect 26789 15487 26847 15493
rect 26789 15484 26801 15487
rect 26660 15456 26801 15484
rect 26660 15444 26666 15456
rect 26789 15453 26801 15456
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 27430 15444 27436 15496
rect 27488 15484 27494 15496
rect 27525 15487 27583 15493
rect 27525 15484 27537 15487
rect 27488 15456 27537 15484
rect 27488 15444 27494 15456
rect 27525 15453 27537 15456
rect 27571 15453 27583 15487
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 27525 15447 27583 15453
rect 27632 15456 28641 15484
rect 24486 15416 24492 15428
rect 22112 15388 24492 15416
rect 20772 15376 20778 15388
rect 24486 15376 24492 15388
rect 24544 15416 24550 15428
rect 27632 15416 27660 15456
rect 28629 15453 28641 15456
rect 28675 15484 28687 15487
rect 28994 15484 29000 15496
rect 28675 15456 29000 15484
rect 28675 15453 28687 15456
rect 28629 15447 28687 15453
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 29730 15484 29736 15496
rect 29691 15456 29736 15484
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 30392 15493 30420 15524
rect 33134 15512 33140 15564
rect 33192 15552 33198 15564
rect 33321 15555 33379 15561
rect 33321 15552 33333 15555
rect 33192 15524 33333 15552
rect 33192 15512 33198 15524
rect 33321 15521 33333 15524
rect 33367 15521 33379 15555
rect 33321 15515 33379 15521
rect 30377 15487 30435 15493
rect 30377 15453 30389 15487
rect 30423 15453 30435 15487
rect 31018 15484 31024 15496
rect 30979 15456 31024 15484
rect 30377 15447 30435 15453
rect 31018 15444 31024 15456
rect 31076 15444 31082 15496
rect 31570 15444 31576 15496
rect 31628 15484 31634 15496
rect 31665 15487 31723 15493
rect 31665 15484 31677 15487
rect 31628 15456 31677 15484
rect 31628 15444 31634 15456
rect 31665 15453 31677 15456
rect 31711 15453 31723 15487
rect 38010 15484 38016 15496
rect 37971 15456 38016 15484
rect 31665 15447 31723 15453
rect 38010 15444 38016 15456
rect 38068 15444 38074 15496
rect 28074 15416 28080 15428
rect 24544 15388 27660 15416
rect 28035 15388 28080 15416
rect 24544 15376 24550 15388
rect 28074 15376 28080 15388
rect 28132 15376 28138 15428
rect 28258 15376 28264 15428
rect 28316 15416 28322 15428
rect 32306 15416 32312 15428
rect 28316 15388 28856 15416
rect 28316 15376 28322 15388
rect 23474 15348 23480 15360
rect 20640 15320 23480 15348
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 23753 15351 23811 15357
rect 23753 15348 23765 15351
rect 23716 15320 23765 15348
rect 23716 15308 23722 15320
rect 23753 15317 23765 15320
rect 23799 15317 23811 15351
rect 23753 15311 23811 15317
rect 24026 15308 24032 15360
rect 24084 15348 24090 15360
rect 25593 15351 25651 15357
rect 25593 15348 25605 15351
rect 24084 15320 25605 15348
rect 24084 15308 24090 15320
rect 25593 15317 25605 15320
rect 25639 15317 25651 15351
rect 25593 15311 25651 15317
rect 25774 15308 25780 15360
rect 25832 15348 25838 15360
rect 26237 15351 26295 15357
rect 26237 15348 26249 15351
rect 25832 15320 26249 15348
rect 25832 15308 25838 15320
rect 26237 15317 26249 15320
rect 26283 15317 26295 15351
rect 26237 15311 26295 15317
rect 26326 15308 26332 15360
rect 26384 15348 26390 15360
rect 28721 15351 28779 15357
rect 28721 15348 28733 15351
rect 26384 15320 28733 15348
rect 26384 15308 26390 15320
rect 28721 15317 28733 15320
rect 28767 15317 28779 15351
rect 28828 15348 28856 15388
rect 28966 15388 32312 15416
rect 28966 15348 28994 15388
rect 32306 15376 32312 15388
rect 32364 15376 32370 15428
rect 33413 15419 33471 15425
rect 33413 15385 33425 15419
rect 33459 15385 33471 15419
rect 33413 15379 33471 15385
rect 34333 15419 34391 15425
rect 34333 15385 34345 15419
rect 34379 15416 34391 15419
rect 34514 15416 34520 15428
rect 34379 15388 34520 15416
rect 34379 15385 34391 15388
rect 34333 15379 34391 15385
rect 28828 15320 28994 15348
rect 28721 15311 28779 15317
rect 30650 15308 30656 15360
rect 30708 15348 30714 15360
rect 31113 15351 31171 15357
rect 31113 15348 31125 15351
rect 30708 15320 31125 15348
rect 30708 15308 30714 15320
rect 31113 15317 31125 15320
rect 31159 15317 31171 15351
rect 31113 15311 31171 15317
rect 32582 15308 32588 15360
rect 32640 15348 32646 15360
rect 33428 15348 33456 15379
rect 34514 15376 34520 15388
rect 34572 15416 34578 15428
rect 35710 15416 35716 15428
rect 34572 15388 35716 15416
rect 34572 15376 34578 15388
rect 35710 15376 35716 15388
rect 35768 15376 35774 15428
rect 38194 15348 38200 15360
rect 32640 15320 33456 15348
rect 38155 15320 38200 15348
rect 32640 15308 32646 15320
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 8478 15104 8484 15156
rect 8536 15144 8542 15156
rect 8536 15116 15608 15144
rect 8536 15104 8542 15116
rect 6914 15076 6920 15088
rect 6875 15048 6920 15076
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 8294 15076 8300 15088
rect 8255 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 10134 15076 10140 15088
rect 10095 15048 10140 15076
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 15378 15076 15384 15088
rect 13754 15048 15384 15076
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 5994 15008 6000 15020
rect 5955 14980 6000 15008
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 14458 14968 14464 15020
rect 14516 15008 14522 15020
rect 14829 15011 14887 15017
rect 14829 15008 14841 15011
rect 14516 14980 14841 15008
rect 14516 14968 14522 14980
rect 14829 14977 14841 14980
rect 14875 15008 14887 15011
rect 15470 15008 15476 15020
rect 14875 14980 15240 15008
rect 15431 14980 15476 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6748 14912 6837 14940
rect 6748 14884 6776 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7064 14912 7481 14940
rect 7064 14900 7070 14912
rect 7469 14909 7481 14912
rect 7515 14940 7527 14943
rect 7834 14940 7840 14952
rect 7515 14912 7840 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 8202 14940 8208 14952
rect 8163 14912 8208 14940
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 6730 14832 6736 14884
rect 6788 14832 6794 14884
rect 1118 14764 1124 14816
rect 1176 14804 1182 14816
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 1176 14776 5825 14804
rect 1176 14764 1182 14776
rect 5813 14773 5825 14776
rect 5859 14773 5871 14807
rect 5813 14767 5871 14773
rect 6086 14764 6092 14816
rect 6144 14804 6150 14816
rect 7650 14804 7656 14816
rect 6144 14776 7656 14804
rect 6144 14764 6150 14776
rect 7650 14764 7656 14776
rect 7708 14804 7714 14816
rect 8496 14804 8524 14903
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 9824 14912 10057 14940
rect 9824 14900 9830 14912
rect 10045 14909 10057 14912
rect 10091 14909 10103 14943
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10045 14903 10103 14909
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 13078 14940 13084 14952
rect 12299 14912 13084 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 14056 14912 14289 14940
rect 14056 14900 14062 14912
rect 14277 14909 14289 14912
rect 14323 14940 14335 14943
rect 15102 14940 15108 14952
rect 14323 14912 15108 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 7708 14776 8524 14804
rect 12516 14807 12574 14813
rect 7708 14764 7714 14776
rect 12516 14773 12528 14807
rect 12562 14804 12574 14807
rect 12894 14804 12900 14816
rect 12562 14776 12900 14804
rect 12562 14773 12574 14776
rect 12516 14767 12574 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 14918 14804 14924 14816
rect 14879 14776 14924 14804
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15212 14804 15240 14980
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 15580 14940 15608 15116
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 16482 15144 16488 15156
rect 15896 15116 16488 15144
rect 15896 15104 15902 15116
rect 16132 15017 16160 15116
rect 16482 15104 16488 15116
rect 16540 15144 16546 15156
rect 16540 15116 20392 15144
rect 16540 15104 16546 15116
rect 16209 15079 16267 15085
rect 16209 15045 16221 15079
rect 16255 15076 16267 15079
rect 18322 15076 18328 15088
rect 16255 15048 18328 15076
rect 16255 15045 16267 15048
rect 16209 15039 16267 15045
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 18690 15076 18696 15088
rect 18651 15048 18696 15076
rect 18690 15036 18696 15048
rect 18748 15036 18754 15088
rect 20364 15076 20392 15116
rect 24394 15104 24400 15156
rect 24452 15144 24458 15156
rect 27338 15144 27344 15156
rect 24452 15116 27344 15144
rect 24452 15104 24458 15116
rect 27338 15104 27344 15116
rect 27396 15104 27402 15156
rect 28166 15104 28172 15156
rect 28224 15144 28230 15156
rect 30098 15144 30104 15156
rect 28224 15116 30104 15144
rect 28224 15104 28230 15116
rect 30098 15104 30104 15116
rect 30156 15104 30162 15156
rect 32401 15147 32459 15153
rect 32401 15113 32413 15147
rect 32447 15144 32459 15147
rect 33410 15144 33416 15156
rect 32447 15116 33416 15144
rect 32447 15113 32459 15116
rect 32401 15107 32459 15113
rect 33410 15104 33416 15116
rect 33468 15104 33474 15156
rect 26142 15076 26148 15088
rect 20364 15048 26148 15076
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17770 15008 17776 15020
rect 17267 14980 17776 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17770 14968 17776 14980
rect 17828 15008 17834 15020
rect 20364 15017 20392 15048
rect 26142 15036 26148 15048
rect 26200 15036 26206 15088
rect 27246 15036 27252 15088
rect 27304 15076 27310 15088
rect 27890 15076 27896 15088
rect 27304 15048 27896 15076
rect 27304 15036 27310 15048
rect 27890 15036 27896 15048
rect 27948 15036 27954 15088
rect 28074 15036 28080 15088
rect 28132 15076 28138 15088
rect 29825 15079 29883 15085
rect 29825 15076 29837 15079
rect 28132 15048 29837 15076
rect 28132 15036 28138 15048
rect 29825 15045 29837 15048
rect 29871 15045 29883 15079
rect 30650 15076 30656 15088
rect 30611 15048 30656 15076
rect 29825 15039 29883 15045
rect 30650 15036 30656 15048
rect 30708 15036 30714 15088
rect 31205 15079 31263 15085
rect 31205 15045 31217 15079
rect 31251 15076 31263 15079
rect 32214 15076 32220 15088
rect 31251 15048 32220 15076
rect 31251 15045 31263 15048
rect 31205 15039 31263 15045
rect 32214 15036 32220 15048
rect 32272 15036 32278 15088
rect 17865 15011 17923 15017
rect 17865 15008 17877 15011
rect 17828 14980 17877 15008
rect 17828 14968 17834 14980
rect 17865 14977 17877 14980
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20806 14968 20812 15020
rect 20864 15008 20870 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 20864 14980 21005 15008
rect 20864 14968 20870 14980
rect 20993 14977 21005 14980
rect 21039 15008 21051 15011
rect 21726 15008 21732 15020
rect 21039 14980 21732 15008
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 21726 14968 21732 14980
rect 21784 15008 21790 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 21784 14980 22293 15008
rect 21784 14968 21790 14980
rect 22281 14977 22293 14980
rect 22327 15008 22339 15011
rect 23661 15011 23719 15017
rect 23661 15008 23673 15011
rect 22327 14980 23673 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 23661 14977 23673 14980
rect 23707 14977 23719 15011
rect 23661 14971 23719 14977
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 24581 15011 24639 15017
rect 24581 15008 24593 15011
rect 23808 14980 24593 15008
rect 23808 14968 23814 14980
rect 24581 14977 24593 14980
rect 24627 14977 24639 15011
rect 24581 14971 24639 14977
rect 25130 14968 25136 15020
rect 25188 15008 25194 15020
rect 25225 15011 25283 15017
rect 25225 15008 25237 15011
rect 25188 14980 25237 15008
rect 25188 14968 25194 14980
rect 25225 14977 25237 14980
rect 25271 14977 25283 15011
rect 25225 14971 25283 14977
rect 25869 15011 25927 15017
rect 25869 14977 25881 15011
rect 25915 14977 25927 15011
rect 25869 14971 25927 14977
rect 18601 14943 18659 14949
rect 18601 14940 18613 14943
rect 15580 14912 18613 14940
rect 18601 14909 18613 14912
rect 18647 14909 18659 14943
rect 18874 14940 18880 14952
rect 18835 14912 18880 14940
rect 18601 14903 18659 14909
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 18966 14900 18972 14952
rect 19024 14940 19030 14952
rect 20441 14943 20499 14949
rect 20441 14940 20453 14943
rect 19024 14912 20453 14940
rect 19024 14900 19030 14912
rect 20441 14909 20453 14912
rect 20487 14909 20499 14943
rect 20441 14903 20499 14909
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14940 21327 14943
rect 21450 14940 21456 14952
rect 21315 14912 21456 14940
rect 21315 14909 21327 14912
rect 21269 14903 21327 14909
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 22922 14900 22928 14952
rect 22980 14940 22986 14952
rect 23017 14943 23075 14949
rect 23017 14940 23029 14943
rect 22980 14912 23029 14940
rect 22980 14900 22986 14912
rect 23017 14909 23029 14912
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 23474 14900 23480 14952
rect 23532 14940 23538 14952
rect 23845 14943 23903 14949
rect 23845 14940 23857 14943
rect 23532 14912 23857 14940
rect 23532 14900 23538 14912
rect 23845 14909 23857 14912
rect 23891 14940 23903 14943
rect 24946 14940 24952 14952
rect 23891 14912 24952 14940
rect 23891 14909 23903 14912
rect 23845 14903 23903 14909
rect 24946 14900 24952 14912
rect 25004 14940 25010 14952
rect 25884 14940 25912 14971
rect 26510 14968 26516 15020
rect 26568 15008 26574 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26568 14980 27169 15008
rect 26568 14968 26574 14980
rect 27157 14977 27169 14980
rect 27203 15008 27215 15011
rect 27522 15008 27528 15020
rect 27203 14980 27528 15008
rect 27203 14977 27215 14980
rect 27157 14971 27215 14977
rect 27522 14968 27528 14980
rect 27580 15008 27586 15020
rect 27801 15011 27859 15017
rect 27801 15008 27813 15011
rect 27580 14980 27813 15008
rect 27580 14968 27586 14980
rect 27801 14977 27813 14980
rect 27847 15008 27859 15011
rect 28445 15011 28503 15017
rect 28445 15008 28457 15011
rect 27847 14980 28457 15008
rect 27847 14977 27859 14980
rect 27801 14971 27859 14977
rect 28445 14977 28457 14980
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 25004 14912 25912 14940
rect 25961 14943 26019 14949
rect 25004 14900 25010 14912
rect 25961 14909 25973 14943
rect 26007 14940 26019 14943
rect 26142 14940 26148 14952
rect 26007 14912 26148 14940
rect 26007 14909 26019 14912
rect 25961 14903 26019 14909
rect 26142 14900 26148 14912
rect 26200 14900 26206 14952
rect 28350 14940 28356 14952
rect 27356 14912 28356 14940
rect 15565 14875 15623 14881
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 17218 14872 17224 14884
rect 15611 14844 17224 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 18892 14872 18920 14900
rect 22554 14872 22560 14884
rect 18892 14844 22560 14872
rect 22554 14832 22560 14844
rect 22612 14832 22618 14884
rect 24302 14832 24308 14884
rect 24360 14872 24366 14884
rect 27356 14872 27384 14912
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 28460 14940 28488 14971
rect 28994 14968 29000 15020
rect 29052 15008 29058 15020
rect 29089 15011 29147 15017
rect 29089 15008 29101 15011
rect 29052 14980 29101 15008
rect 29052 14968 29058 14980
rect 29089 14977 29101 14980
rect 29135 14977 29147 15011
rect 29730 15008 29736 15020
rect 29691 14980 29736 15008
rect 29089 14971 29147 14977
rect 29730 14968 29736 14980
rect 29788 14968 29794 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 31726 14980 32321 15008
rect 29638 14940 29644 14952
rect 28460 14912 29644 14940
rect 29638 14900 29644 14912
rect 29696 14900 29702 14952
rect 29822 14900 29828 14952
rect 29880 14940 29886 14952
rect 30561 14943 30619 14949
rect 30561 14940 30573 14943
rect 29880 14912 30573 14940
rect 29880 14900 29886 14912
rect 30561 14909 30573 14912
rect 30607 14909 30619 14943
rect 30561 14903 30619 14909
rect 24360 14844 27384 14872
rect 24360 14832 24366 14844
rect 27430 14832 27436 14884
rect 27488 14872 27494 14884
rect 29181 14875 29239 14881
rect 29181 14872 29193 14875
rect 27488 14844 29193 14872
rect 27488 14832 27494 14844
rect 29181 14841 29193 14844
rect 29227 14841 29239 14875
rect 29181 14835 29239 14841
rect 29362 14832 29368 14884
rect 29420 14872 29426 14884
rect 29914 14872 29920 14884
rect 29420 14844 29920 14872
rect 29420 14832 29426 14844
rect 29914 14832 29920 14844
rect 29972 14832 29978 14884
rect 16390 14804 16396 14816
rect 15212 14776 16396 14804
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17313 14807 17371 14813
rect 17313 14804 17325 14807
rect 17000 14776 17325 14804
rect 17000 14764 17006 14776
rect 17313 14773 17325 14776
rect 17359 14773 17371 14807
rect 17313 14767 17371 14773
rect 17957 14807 18015 14813
rect 17957 14773 17969 14807
rect 18003 14804 18015 14807
rect 19058 14804 19064 14816
rect 18003 14776 19064 14804
rect 18003 14773 18015 14776
rect 17957 14767 18015 14773
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 20530 14804 20536 14816
rect 19392 14776 20536 14804
rect 19392 14764 19398 14776
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 24118 14764 24124 14816
rect 24176 14804 24182 14816
rect 24673 14807 24731 14813
rect 24673 14804 24685 14807
rect 24176 14776 24685 14804
rect 24176 14764 24182 14776
rect 24673 14773 24685 14776
rect 24719 14773 24731 14807
rect 24673 14767 24731 14773
rect 24946 14764 24952 14816
rect 25004 14804 25010 14816
rect 25317 14807 25375 14813
rect 25317 14804 25329 14807
rect 25004 14776 25329 14804
rect 25004 14764 25010 14776
rect 25317 14773 25329 14776
rect 25363 14773 25375 14807
rect 25317 14767 25375 14773
rect 26050 14764 26056 14816
rect 26108 14804 26114 14816
rect 27249 14807 27307 14813
rect 27249 14804 27261 14807
rect 26108 14776 27261 14804
rect 26108 14764 26114 14776
rect 27249 14773 27261 14776
rect 27295 14773 27307 14807
rect 27249 14767 27307 14773
rect 27706 14764 27712 14816
rect 27764 14804 27770 14816
rect 27893 14807 27951 14813
rect 27893 14804 27905 14807
rect 27764 14776 27905 14804
rect 27764 14764 27770 14776
rect 27893 14773 27905 14776
rect 27939 14773 27951 14807
rect 27893 14767 27951 14773
rect 28442 14764 28448 14816
rect 28500 14804 28506 14816
rect 28537 14807 28595 14813
rect 28537 14804 28549 14807
rect 28500 14776 28549 14804
rect 28500 14764 28506 14776
rect 28537 14773 28549 14776
rect 28583 14773 28595 14807
rect 28537 14767 28595 14773
rect 28994 14764 29000 14816
rect 29052 14804 29058 14816
rect 31726 14804 31754 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 38013 15011 38071 15017
rect 38013 14977 38025 15011
rect 38059 15008 38071 15011
rect 38102 15008 38108 15020
rect 38059 14980 38108 15008
rect 38059 14977 38071 14980
rect 38013 14971 38071 14977
rect 38102 14968 38108 14980
rect 38160 14968 38166 15020
rect 37826 14804 37832 14816
rect 29052 14776 31754 14804
rect 37787 14776 37832 14804
rect 29052 14764 29058 14776
rect 37826 14764 37832 14776
rect 37884 14764 37890 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 2225 14603 2283 14609
rect 2225 14569 2237 14603
rect 2271 14600 2283 14603
rect 2314 14600 2320 14612
rect 2271 14572 2320 14600
rect 2271 14569 2283 14572
rect 2225 14563 2283 14569
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 2240 14396 2268 14563
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 9030 14600 9036 14612
rect 6604 14572 9036 14600
rect 6604 14560 6610 14572
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 17221 14603 17279 14609
rect 10100 14572 16160 14600
rect 10100 14560 10106 14572
rect 8570 14532 8576 14544
rect 5552 14504 8576 14532
rect 5552 14473 5580 14504
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 11974 14492 11980 14544
rect 12032 14532 12038 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 12032 14504 13645 14532
rect 12032 14492 12038 14504
rect 13633 14501 13645 14504
rect 13679 14501 13691 14535
rect 13633 14495 13691 14501
rect 14016 14504 16068 14532
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14433 5595 14467
rect 5537 14427 5595 14433
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 5960 14436 7573 14464
rect 5960 14424 5966 14436
rect 7561 14433 7573 14436
rect 7607 14464 7619 14467
rect 8202 14464 8208 14476
rect 7607 14436 8208 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8478 14464 8484 14476
rect 8439 14436 8484 14464
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 11057 14467 11115 14473
rect 9732 14436 9777 14464
rect 9732 14424 9738 14436
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 13906 14464 13912 14476
rect 11103 14436 13912 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 1627 14368 2268 14396
rect 10965 14399 11023 14405
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11011 14368 11621 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11609 14365 11621 14368
rect 11655 14396 11667 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 11655 14368 12265 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 5629 14331 5687 14337
rect 5629 14297 5641 14331
rect 5675 14328 5687 14331
rect 5902 14328 5908 14340
rect 5675 14300 5908 14328
rect 5675 14297 5687 14300
rect 5629 14291 5687 14297
rect 5902 14288 5908 14300
rect 5960 14288 5966 14340
rect 6546 14328 6552 14340
rect 6507 14300 6552 14328
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 7558 14288 7564 14340
rect 7616 14328 7622 14340
rect 7653 14331 7711 14337
rect 7653 14328 7665 14331
rect 7616 14300 7665 14328
rect 7616 14288 7622 14300
rect 7653 14297 7665 14300
rect 7699 14297 7711 14331
rect 9306 14328 9312 14340
rect 9267 14300 9312 14328
rect 7653 14291 7711 14297
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 9416 14260 9444 14291
rect 7524 14232 9444 14260
rect 11701 14263 11759 14269
rect 7524 14220 7530 14232
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12158 14260 12164 14272
rect 11747 14232 12164 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 12268 14260 12296 14359
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12894 14396 12900 14408
rect 12492 14368 12900 14396
rect 12492 14356 12498 14368
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 13262 14396 13268 14408
rect 13035 14368 13268 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 14016 14396 14044 14504
rect 15930 14464 15936 14476
rect 14568 14436 15936 14464
rect 14568 14405 14596 14436
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 13587 14368 14044 14396
rect 14108 14368 14565 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 12345 14331 12403 14337
rect 12345 14297 12357 14331
rect 12391 14328 12403 14331
rect 13998 14328 14004 14340
rect 12391 14300 14004 14328
rect 12391 14297 12403 14300
rect 12345 14291 12403 14297
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 14108 14260 14136 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 15194 14396 15200 14408
rect 15155 14368 15200 14396
rect 14553 14359 14611 14365
rect 15194 14356 15200 14368
rect 15252 14396 15258 14408
rect 15470 14396 15476 14408
rect 15252 14368 15476 14396
rect 15252 14356 15258 14368
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16040 14396 16068 14504
rect 15887 14368 16068 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 16040 14272 16068 14368
rect 16132 14328 16160 14572
rect 17221 14569 17233 14603
rect 17267 14600 17279 14603
rect 18690 14600 18696 14612
rect 17267 14572 18696 14600
rect 17267 14569 17279 14572
rect 17221 14563 17279 14569
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 19334 14600 19340 14612
rect 18800 14572 19340 14600
rect 18800 14532 18828 14572
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 20162 14560 20168 14612
rect 20220 14600 20226 14612
rect 21266 14600 21272 14612
rect 20220 14572 21272 14600
rect 20220 14560 20226 14572
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 23845 14603 23903 14609
rect 23845 14600 23857 14603
rect 22612 14572 23857 14600
rect 22612 14560 22618 14572
rect 23845 14569 23857 14572
rect 23891 14569 23903 14603
rect 23845 14563 23903 14569
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 26786 14600 26792 14612
rect 25188 14572 26792 14600
rect 25188 14560 25194 14572
rect 26786 14560 26792 14572
rect 26844 14560 26850 14612
rect 28902 14600 28908 14612
rect 28863 14572 28908 14600
rect 28902 14560 28908 14572
rect 28960 14560 28966 14612
rect 37369 14603 37427 14609
rect 37369 14569 37381 14603
rect 37415 14600 37427 14603
rect 38010 14600 38016 14612
rect 37415 14572 38016 14600
rect 37415 14569 37427 14572
rect 37369 14563 37427 14569
rect 38010 14560 38016 14572
rect 38068 14560 38074 14612
rect 16500 14504 18828 14532
rect 16500 14408 16528 14504
rect 22370 14492 22376 14544
rect 22428 14532 22434 14544
rect 23750 14532 23756 14544
rect 22428 14504 23756 14532
rect 22428 14492 22434 14504
rect 23750 14492 23756 14504
rect 23808 14492 23814 14544
rect 27338 14492 27344 14544
rect 27396 14532 27402 14544
rect 29730 14532 29736 14544
rect 27396 14504 29736 14532
rect 27396 14492 27402 14504
rect 29730 14492 29736 14504
rect 29788 14532 29794 14544
rect 29788 14504 31248 14532
rect 29788 14492 29794 14504
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 16908 14436 19461 14464
rect 16908 14424 16914 14436
rect 16482 14396 16488 14408
rect 16395 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 17126 14396 17132 14408
rect 16632 14368 16677 14396
rect 17087 14368 17132 14396
rect 16632 14356 16638 14368
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 19334 14396 19340 14408
rect 18708 14368 19340 14396
rect 17865 14331 17923 14337
rect 17865 14328 17877 14331
rect 16132 14300 17877 14328
rect 17865 14297 17877 14300
rect 17911 14297 17923 14331
rect 17865 14291 17923 14297
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 18708 14328 18736 14368
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19433 14405 19461 14436
rect 22186 14424 22192 14476
rect 22244 14464 22250 14476
rect 23014 14464 23020 14476
rect 22244 14436 23020 14464
rect 22244 14424 22250 14436
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25501 14467 25559 14473
rect 25501 14464 25513 14467
rect 24912 14436 25513 14464
rect 24912 14424 24918 14436
rect 25501 14433 25513 14436
rect 25547 14464 25559 14467
rect 26234 14464 26240 14476
rect 25547 14436 26240 14464
rect 25547 14433 25559 14436
rect 25501 14427 25559 14433
rect 26234 14424 26240 14436
rect 26292 14424 26298 14476
rect 27246 14424 27252 14476
rect 27304 14464 27310 14476
rect 27304 14436 28856 14464
rect 27304 14424 27310 14436
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 21726 14396 21732 14408
rect 21687 14368 21732 14396
rect 19429 14359 19487 14365
rect 21726 14356 21732 14368
rect 21784 14396 21790 14408
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 21784 14368 22845 14396
rect 21784 14356 21790 14368
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 23750 14396 23756 14408
rect 23711 14368 23756 14396
rect 22833 14359 22891 14365
rect 23750 14356 23756 14368
rect 23808 14356 23814 14408
rect 24486 14356 24492 14408
rect 24544 14396 24550 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24544 14368 24593 14396
rect 24544 14356 24550 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 27154 14396 27160 14408
rect 26910 14368 27160 14396
rect 24581 14359 24639 14365
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 27525 14399 27583 14405
rect 27525 14396 27537 14399
rect 27448 14368 27537 14396
rect 18874 14328 18880 14340
rect 18012 14300 18057 14328
rect 18156 14300 18736 14328
rect 18835 14300 18880 14328
rect 18012 14288 18018 14300
rect 14642 14260 14648 14272
rect 12268 14232 14136 14260
rect 14603 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 15286 14260 15292 14272
rect 15247 14232 15292 14260
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15896 14232 15945 14260
rect 15896 14220 15902 14232
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 15933 14223 15991 14229
rect 16022 14220 16028 14272
rect 16080 14260 16086 14272
rect 16298 14260 16304 14272
rect 16080 14232 16304 14260
rect 16080 14220 16086 14232
rect 16298 14220 16304 14232
rect 16356 14260 16362 14272
rect 18156 14260 18184 14300
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 19242 14288 19248 14340
rect 19300 14328 19306 14340
rect 19705 14331 19763 14337
rect 19705 14328 19717 14331
rect 19300 14300 19717 14328
rect 19300 14288 19306 14300
rect 19705 14297 19717 14300
rect 19751 14297 19763 14331
rect 22281 14331 22339 14337
rect 19705 14291 19763 14297
rect 19812 14300 20194 14328
rect 16356 14232 18184 14260
rect 16356 14220 16362 14232
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 19260 14260 19288 14288
rect 18748 14232 19288 14260
rect 18748 14220 18754 14232
rect 19518 14220 19524 14272
rect 19576 14260 19582 14272
rect 19812 14260 19840 14300
rect 22281 14297 22293 14331
rect 22327 14328 22339 14331
rect 22462 14328 22468 14340
rect 22327 14300 22468 14328
rect 22327 14297 22339 14300
rect 22281 14291 22339 14297
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 24673 14331 24731 14337
rect 24673 14328 24685 14331
rect 23400 14300 24685 14328
rect 19576 14232 19840 14260
rect 19576 14220 19582 14232
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 21177 14263 21235 14269
rect 21177 14260 21189 14263
rect 20036 14232 21189 14260
rect 20036 14220 20042 14232
rect 21177 14229 21189 14232
rect 21223 14229 21235 14263
rect 21177 14223 21235 14229
rect 21726 14220 21732 14272
rect 21784 14260 21790 14272
rect 23400 14260 23428 14300
rect 24673 14297 24685 14300
rect 24719 14297 24731 14331
rect 24673 14291 24731 14297
rect 25777 14331 25835 14337
rect 25777 14297 25789 14331
rect 25823 14297 25835 14331
rect 25777 14291 25835 14297
rect 21784 14232 23428 14260
rect 25792 14260 25820 14291
rect 27338 14288 27344 14340
rect 27396 14328 27402 14340
rect 27448 14328 27476 14368
rect 27525 14365 27537 14368
rect 27571 14365 27583 14399
rect 27525 14359 27583 14365
rect 27614 14356 27620 14408
rect 27672 14396 27678 14408
rect 28828 14405 28856 14436
rect 31220 14405 31248 14504
rect 27985 14399 28043 14405
rect 27985 14396 27997 14399
rect 27672 14368 27997 14396
rect 27672 14356 27678 14368
rect 27985 14365 27997 14368
rect 28031 14365 28043 14399
rect 27985 14359 28043 14365
rect 28813 14399 28871 14405
rect 28813 14365 28825 14399
rect 28859 14365 28871 14399
rect 28813 14359 28871 14365
rect 31205 14399 31263 14405
rect 31205 14365 31217 14399
rect 31251 14396 31263 14399
rect 33042 14396 33048 14408
rect 31251 14368 33048 14396
rect 31251 14365 31263 14368
rect 31205 14359 31263 14365
rect 33042 14356 33048 14368
rect 33100 14356 33106 14408
rect 37550 14396 37556 14408
rect 37511 14368 37556 14396
rect 37550 14356 37556 14368
rect 37608 14356 37614 14408
rect 37918 14356 37924 14408
rect 37976 14396 37982 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 37976 14368 38025 14396
rect 37976 14356 37982 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 29362 14328 29368 14340
rect 27396 14300 27476 14328
rect 27540 14300 29368 14328
rect 27396 14288 27402 14300
rect 27540 14260 27568 14300
rect 29362 14288 29368 14300
rect 29420 14288 29426 14340
rect 29822 14288 29828 14340
rect 29880 14328 29886 14340
rect 30101 14331 30159 14337
rect 30101 14328 30113 14331
rect 29880 14300 30113 14328
rect 29880 14288 29886 14300
rect 30101 14297 30113 14300
rect 30147 14297 30159 14331
rect 30101 14291 30159 14297
rect 30190 14288 30196 14340
rect 30248 14328 30254 14340
rect 30745 14331 30803 14337
rect 30248 14300 30293 14328
rect 30248 14288 30254 14300
rect 30745 14297 30757 14331
rect 30791 14328 30803 14331
rect 31478 14328 31484 14340
rect 30791 14300 31484 14328
rect 30791 14297 30803 14300
rect 30745 14291 30803 14297
rect 31478 14288 31484 14300
rect 31536 14288 31542 14340
rect 25792 14232 27568 14260
rect 21784 14220 21790 14232
rect 27614 14220 27620 14272
rect 27672 14260 27678 14272
rect 28077 14263 28135 14269
rect 28077 14260 28089 14263
rect 27672 14232 28089 14260
rect 27672 14220 27678 14232
rect 28077 14229 28089 14232
rect 28123 14229 28135 14263
rect 28077 14223 28135 14229
rect 30650 14220 30656 14272
rect 30708 14260 30714 14272
rect 31297 14263 31355 14269
rect 31297 14260 31309 14263
rect 30708 14232 31309 14260
rect 30708 14220 30714 14232
rect 31297 14229 31309 14232
rect 31343 14229 31355 14263
rect 31297 14223 31355 14229
rect 37458 14220 37464 14272
rect 37516 14260 37522 14272
rect 37918 14260 37924 14272
rect 37516 14232 37924 14260
rect 37516 14220 37522 14232
rect 37918 14220 37924 14232
rect 37976 14220 37982 14272
rect 38194 14260 38200 14272
rect 38155 14232 38200 14260
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 5902 14056 5908 14068
rect 5863 14028 5908 14056
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 7432 14028 7481 14056
rect 7432 14016 7438 14028
rect 7469 14025 7481 14028
rect 7515 14025 7527 14059
rect 7469 14019 7527 14025
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8294 14056 8300 14068
rect 8159 14028 8300 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8444 14028 8769 14056
rect 8444 14016 8450 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 10042 14056 10048 14068
rect 8757 14019 8815 14025
rect 9232 14028 10048 14056
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5500 13892 5825 13920
rect 5500 13880 5506 13892
rect 5813 13889 5825 13892
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7006 13920 7012 13932
rect 6779 13892 7012 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 8018 13920 8024 13932
rect 7979 13892 8024 13920
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 9232 13920 9260 14028
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 11882 14056 11888 14068
rect 11103 14028 11888 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 15286 14056 15292 14068
rect 11992 14028 15292 14056
rect 9490 13988 9496 14000
rect 9451 13960 9496 13988
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 10410 13948 10416 14000
rect 10468 13988 10474 14000
rect 11992 13988 12020 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18690 14056 18696 14068
rect 18647 14028 18696 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 18874 14016 18880 14068
rect 18932 14056 18938 14068
rect 19150 14056 19156 14068
rect 18932 14028 19156 14056
rect 18932 14016 18938 14028
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21416 14028 21465 14056
rect 21416 14016 21422 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 21542 14016 21548 14068
rect 21600 14056 21606 14068
rect 22278 14056 22284 14068
rect 21600 14028 22284 14056
rect 21600 14016 21606 14028
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 23750 14016 23756 14068
rect 23808 14056 23814 14068
rect 23845 14059 23903 14065
rect 23845 14056 23857 14059
rect 23808 14028 23857 14056
rect 23808 14016 23814 14028
rect 23845 14025 23857 14028
rect 23891 14056 23903 14059
rect 23934 14056 23940 14068
rect 23891 14028 23940 14056
rect 23891 14025 23903 14028
rect 23845 14019 23903 14025
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 27706 14056 27712 14068
rect 25516 14028 27712 14056
rect 13354 13988 13360 14000
rect 10468 13960 12020 13988
rect 13315 13960 13360 13988
rect 10468 13948 10474 13960
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 13814 13948 13820 14000
rect 13872 13948 13878 14000
rect 15102 13948 15108 14000
rect 15160 13988 15166 14000
rect 17129 13991 17187 13997
rect 15160 13960 15240 13988
rect 15160 13948 15166 13960
rect 8711 13892 9260 13920
rect 10965 13923 11023 13929
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 10965 13889 10977 13923
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12986 13920 12992 13932
rect 12299 13892 12992 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 8680 13824 9168 13852
rect 8680 13796 8708 13824
rect 8662 13744 8668 13796
rect 8720 13744 8726 13796
rect 9140 13784 9168 13824
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9401 13855 9459 13861
rect 9401 13852 9413 13855
rect 9272 13824 9413 13852
rect 9272 13812 9278 13824
rect 9401 13821 9413 13824
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9640 13824 9689 13852
rect 9640 13812 9646 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 10980 13852 11008 13883
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 12342 13852 12348 13864
rect 9677 13815 9735 13821
rect 9784 13824 11008 13852
rect 12303 13824 12348 13852
rect 9784 13784 9812 13824
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 13078 13852 13084 13864
rect 13039 13824 13084 13852
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13188 13824 14412 13852
rect 9140 13756 9812 13784
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 13188 13784 13216 13824
rect 12584 13756 13216 13784
rect 14384 13784 14412 13824
rect 14826 13812 14832 13864
rect 14884 13852 14890 13864
rect 15105 13855 15163 13861
rect 15105 13852 15117 13855
rect 14884 13824 15117 13852
rect 14884 13812 14890 13824
rect 15105 13821 15117 13824
rect 15151 13821 15163 13855
rect 15212 13852 15240 13960
rect 17129 13957 17141 13991
rect 17175 13988 17187 13991
rect 17402 13988 17408 14000
rect 17175 13960 17408 13988
rect 17175 13957 17187 13960
rect 17129 13951 17187 13957
rect 17402 13948 17408 13960
rect 17460 13948 17466 14000
rect 17678 13948 17684 14000
rect 17736 13948 17742 14000
rect 18782 13948 18788 14000
rect 18840 13988 18846 14000
rect 19334 13988 19340 14000
rect 18840 13960 19340 13988
rect 18840 13948 18846 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 20714 13948 20720 14000
rect 20772 13948 20778 14000
rect 25516 13988 25544 14028
rect 27706 14016 27712 14028
rect 27764 14016 27770 14068
rect 28442 14056 28448 14068
rect 27816 14028 28448 14056
rect 27816 13988 27844 14028
rect 28442 14016 28448 14028
rect 28500 14016 28506 14068
rect 30009 14059 30067 14065
rect 30009 14025 30021 14059
rect 30055 14056 30067 14059
rect 30190 14056 30196 14068
rect 30055 14028 30196 14056
rect 30055 14025 30067 14028
rect 30009 14019 30067 14025
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 23598 13960 25544 13988
rect 26358 13960 27844 13988
rect 27982 13948 27988 14000
rect 28040 13948 28046 14000
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16482 13920 16488 13932
rect 16163 13892 16488 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16850 13920 16856 13932
rect 16811 13892 16856 13920
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13920 19119 13923
rect 19610 13920 19616 13932
rect 19107 13892 19616 13920
rect 19107 13889 19119 13892
rect 19061 13883 19119 13889
rect 19610 13880 19616 13892
rect 19668 13880 19674 13932
rect 24854 13920 24860 13932
rect 24815 13892 24860 13920
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 29086 13880 29092 13932
rect 29144 13920 29150 13932
rect 29917 13923 29975 13929
rect 29917 13920 29929 13923
rect 29144 13892 29929 13920
rect 29144 13880 29150 13892
rect 29917 13889 29929 13892
rect 29963 13889 29975 13923
rect 30558 13920 30564 13932
rect 30519 13892 30564 13920
rect 29917 13883 29975 13889
rect 30558 13880 30564 13892
rect 30616 13920 30622 13932
rect 30926 13920 30932 13932
rect 30616 13892 30932 13920
rect 30616 13880 30622 13892
rect 30926 13880 30932 13892
rect 30984 13880 30990 13932
rect 18414 13852 18420 13864
rect 15212 13824 18420 13852
rect 15105 13815 15163 13821
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 19153 13855 19211 13861
rect 19153 13821 19165 13855
rect 19199 13852 19211 13855
rect 19334 13852 19340 13864
rect 19199 13824 19340 13852
rect 19199 13821 19211 13824
rect 19153 13815 19211 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19484 13824 19717 13852
rect 19484 13812 19490 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19978 13852 19984 13864
rect 19939 13824 19984 13852
rect 19705 13815 19763 13821
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 22152 13824 22197 13852
rect 24964 13824 26617 13852
rect 22152 13812 22158 13824
rect 14384 13756 16344 13784
rect 12584 13744 12590 13756
rect 7282 13676 7288 13728
rect 7340 13716 7346 13728
rect 11606 13716 11612 13728
rect 7340 13688 11612 13716
rect 7340 13676 7346 13688
rect 11606 13676 11612 13688
rect 11664 13716 11670 13728
rect 14458 13716 14464 13728
rect 11664 13688 14464 13716
rect 11664 13676 11670 13688
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15930 13716 15936 13728
rect 15252 13688 15936 13716
rect 15252 13676 15258 13688
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16206 13716 16212 13728
rect 16167 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 16316 13716 16344 13756
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 18690 13784 18696 13796
rect 18288 13756 18696 13784
rect 18288 13744 18294 13756
rect 18690 13744 18696 13756
rect 18748 13744 18754 13796
rect 21174 13744 21180 13796
rect 21232 13784 21238 13796
rect 22002 13784 22008 13796
rect 21232 13756 22008 13784
rect 21232 13744 21238 13756
rect 22002 13744 22008 13756
rect 22060 13744 22066 13796
rect 24964 13784 24992 13824
rect 26605 13821 26617 13824
rect 26651 13852 26663 13855
rect 26694 13852 26700 13864
rect 26651 13824 26700 13852
rect 26651 13821 26663 13824
rect 26605 13815 26663 13821
rect 26694 13812 26700 13824
rect 26752 13812 26758 13864
rect 27154 13852 27160 13864
rect 26804 13824 27160 13852
rect 24412 13756 24992 13784
rect 21192 13716 21220 13744
rect 16316 13688 21220 13716
rect 22360 13719 22418 13725
rect 22360 13685 22372 13719
rect 22406 13716 22418 13719
rect 24412 13716 24440 13756
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 26804 13784 26832 13824
rect 27154 13812 27160 13824
rect 27212 13812 27218 13864
rect 27433 13855 27491 13861
rect 27433 13852 27445 13855
rect 27264 13824 27445 13852
rect 26292 13756 26832 13784
rect 26292 13744 26298 13756
rect 26970 13744 26976 13796
rect 27028 13784 27034 13796
rect 27264 13784 27292 13824
rect 27433 13821 27445 13824
rect 27479 13852 27491 13855
rect 27522 13852 27528 13864
rect 27479 13824 27528 13852
rect 27479 13821 27491 13824
rect 27433 13815 27491 13821
rect 27522 13812 27528 13824
rect 27580 13812 27586 13864
rect 28442 13812 28448 13864
rect 28500 13852 28506 13864
rect 29181 13855 29239 13861
rect 29181 13852 29193 13855
rect 28500 13824 29193 13852
rect 28500 13812 28506 13824
rect 29181 13821 29193 13824
rect 29227 13821 29239 13855
rect 30653 13855 30711 13861
rect 30653 13852 30665 13855
rect 29181 13815 29239 13821
rect 29288 13824 30665 13852
rect 27028 13756 27292 13784
rect 27028 13744 27034 13756
rect 28902 13744 28908 13796
rect 28960 13784 28966 13796
rect 29086 13784 29092 13796
rect 28960 13756 29092 13784
rect 28960 13744 28966 13756
rect 29086 13744 29092 13756
rect 29144 13744 29150 13796
rect 25130 13725 25136 13728
rect 22406 13688 24440 13716
rect 25120 13719 25136 13725
rect 22406 13685 22418 13688
rect 22360 13679 22418 13685
rect 25120 13685 25132 13719
rect 25120 13679 25136 13685
rect 25130 13676 25136 13679
rect 25188 13676 25194 13728
rect 25498 13676 25504 13728
rect 25556 13716 25562 13728
rect 29288 13716 29316 13824
rect 30653 13821 30665 13824
rect 30699 13821 30711 13855
rect 30653 13815 30711 13821
rect 30558 13744 30564 13796
rect 30616 13784 30622 13796
rect 30834 13784 30840 13796
rect 30616 13756 30840 13784
rect 30616 13744 30622 13756
rect 30834 13744 30840 13756
rect 30892 13744 30898 13796
rect 25556 13688 29316 13716
rect 25556 13676 25562 13688
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 9217 13515 9275 13521
rect 9217 13481 9229 13515
rect 9263 13512 9275 13515
rect 9306 13512 9312 13524
rect 9263 13484 9312 13512
rect 9263 13481 9275 13484
rect 9217 13475 9275 13481
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13444 1823 13447
rect 2038 13444 2044 13456
rect 1811 13416 2044 13444
rect 1811 13413 1823 13416
rect 1765 13407 1823 13413
rect 2038 13404 2044 13416
rect 2096 13444 2102 13456
rect 5534 13444 5540 13456
rect 2096 13416 5540 13444
rect 2096 13404 2102 13416
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 8386 13376 8392 13388
rect 7607 13348 8392 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 8386 13336 8392 13348
rect 8444 13376 8450 13388
rect 9232 13376 9260 13475
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9490 13472 9496 13524
rect 9548 13512 9554 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 9548 13484 10057 13512
rect 9548 13472 9554 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10192 13484 10701 13512
rect 10192 13472 10198 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 11964 13515 12022 13521
rect 11964 13481 11976 13515
rect 12010 13512 12022 13515
rect 12526 13512 12532 13524
rect 12010 13484 12532 13512
rect 12010 13481 12022 13484
rect 11964 13475 12022 13481
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 15933 13515 15991 13521
rect 15933 13512 15945 13515
rect 15436 13484 15945 13512
rect 15436 13472 15442 13484
rect 15933 13481 15945 13484
rect 15979 13481 15991 13515
rect 15933 13475 15991 13481
rect 16592 13484 18000 13512
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 16592 13444 16620 13484
rect 13412 13416 16620 13444
rect 13412 13404 13418 13416
rect 8444 13348 9260 13376
rect 11701 13379 11759 13385
rect 8444 13336 8450 13348
rect 11701 13345 11713 13379
rect 11747 13376 11759 13379
rect 12986 13376 12992 13388
rect 11747 13348 12992 13376
rect 11747 13345 11759 13348
rect 11701 13339 11759 13345
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 16206 13376 16212 13388
rect 13096 13348 16212 13376
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13308 4399 13311
rect 5166 13308 5172 13320
rect 4387 13280 5172 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 7190 13308 7196 13320
rect 6871 13280 7196 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13308 10011 13311
rect 10042 13308 10048 13320
rect 9999 13280 10048 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10870 13308 10876 13320
rect 10643 13280 10876 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 13096 13294 13124 13348
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 16850 13376 16856 13388
rect 16531 13348 16856 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 16850 13336 16856 13348
rect 16908 13376 16914 13388
rect 17770 13376 17776 13388
rect 16908 13348 17776 13376
rect 16908 13336 16914 13348
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 17972 13376 18000 13484
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18506 13512 18512 13524
rect 18104 13484 18512 13512
rect 18104 13472 18110 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 20714 13512 20720 13524
rect 20180 13484 20720 13512
rect 20180 13444 20208 13484
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 21266 13512 21272 13524
rect 20824 13484 21272 13512
rect 18524 13416 20208 13444
rect 18524 13385 18552 13416
rect 18509 13379 18567 13385
rect 18509 13376 18521 13379
rect 17972 13348 18521 13376
rect 18509 13345 18521 13348
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13688 13280 13737 13308
rect 13688 13268 13694 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 15194 13308 15200 13320
rect 15155 13280 15200 13308
rect 13725 13271 13783 13277
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15344 13280 15389 13308
rect 15344 13268 15350 13280
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 15528 13280 15853 13308
rect 15528 13268 15534 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19610 13308 19616 13320
rect 19475 13280 19616 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19610 13268 19616 13280
rect 19668 13268 19674 13320
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20254 13308 20260 13320
rect 20119 13280 20260 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 20254 13268 20260 13280
rect 20312 13308 20318 13320
rect 20530 13308 20536 13320
rect 20312 13280 20536 13308
rect 20312 13268 20318 13280
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 20824 13308 20852 13484
rect 21266 13472 21272 13484
rect 21324 13512 21330 13524
rect 22370 13512 22376 13524
rect 21324 13484 22376 13512
rect 21324 13472 21330 13484
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 23198 13472 23204 13524
rect 23256 13512 23262 13524
rect 23256 13484 24900 13512
rect 23256 13472 23262 13484
rect 22922 13404 22928 13456
rect 22980 13444 22986 13456
rect 24486 13444 24492 13456
rect 22980 13416 24492 13444
rect 22980 13404 22986 13416
rect 24486 13404 24492 13416
rect 24544 13404 24550 13456
rect 20898 13336 20904 13388
rect 20956 13336 20962 13388
rect 22186 13376 22192 13388
rect 21376 13348 22192 13376
rect 20763 13280 20852 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 7653 13243 7711 13249
rect 7653 13209 7665 13243
rect 7699 13209 7711 13243
rect 8570 13240 8576 13252
rect 8531 13212 8576 13240
rect 7653 13203 7711 13209
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4028 13144 4353 13172
rect 4028 13132 4034 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7668 13172 7696 13203
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 14332 13212 14964 13240
rect 14332 13200 14338 13212
rect 6963 13144 7696 13172
rect 14936 13172 14964 13212
rect 16482 13200 16488 13252
rect 16540 13240 16546 13252
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 16540 13212 16773 13240
rect 16540 13200 16546 13212
rect 16761 13209 16773 13212
rect 16807 13209 16819 13243
rect 16761 13203 16819 13209
rect 17218 13200 17224 13252
rect 17276 13200 17282 13252
rect 20916 13240 20944 13336
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 21376 13317 21404 13348
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 23382 13376 23388 13388
rect 22704 13348 23388 13376
rect 22704 13336 22710 13348
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 24762 13376 24768 13388
rect 24723 13348 24768 13376
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 24872 13376 24900 13484
rect 37550 13472 37556 13524
rect 37608 13512 37614 13524
rect 38105 13515 38163 13521
rect 38105 13512 38117 13515
rect 37608 13484 38117 13512
rect 37608 13472 37614 13484
rect 38105 13481 38117 13484
rect 38151 13481 38163 13515
rect 38105 13475 38163 13481
rect 26326 13444 26332 13456
rect 26068 13416 26332 13444
rect 26068 13376 26096 13416
rect 26326 13404 26332 13416
rect 26384 13444 26390 13456
rect 26878 13444 26884 13456
rect 26384 13416 26884 13444
rect 26384 13404 26390 13416
rect 26878 13404 26884 13416
rect 26936 13404 26942 13456
rect 27706 13404 27712 13456
rect 27764 13444 27770 13456
rect 27890 13444 27896 13456
rect 27764 13416 27896 13444
rect 27764 13404 27770 13416
rect 27890 13404 27896 13416
rect 27948 13404 27954 13456
rect 24872 13348 26096 13376
rect 27154 13336 27160 13388
rect 27212 13376 27218 13388
rect 27985 13379 28043 13385
rect 27985 13376 27997 13379
rect 27212 13348 27997 13376
rect 27212 13336 27218 13348
rect 27985 13345 27997 13348
rect 28031 13345 28043 13379
rect 27985 13339 28043 13345
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 21232 13280 21373 13308
rect 21232 13268 21238 13280
rect 21361 13277 21373 13280
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23845 13311 23903 13317
rect 23845 13308 23857 13311
rect 23532 13280 23857 13308
rect 23532 13268 23538 13280
rect 23845 13277 23857 13280
rect 23891 13277 23903 13311
rect 28074 13308 28080 13320
rect 26174 13280 28080 13308
rect 23845 13271 23903 13277
rect 28074 13268 28080 13280
rect 28132 13268 28138 13320
rect 33321 13311 33379 13317
rect 33321 13277 33333 13311
rect 33367 13308 33379 13311
rect 33870 13308 33876 13320
rect 33367 13280 33876 13308
rect 33367 13277 33379 13280
rect 33321 13271 33379 13277
rect 33870 13268 33876 13280
rect 33928 13268 33934 13320
rect 38286 13308 38292 13320
rect 38247 13280 38292 13308
rect 38286 13268 38292 13280
rect 38344 13268 38350 13320
rect 18064 13212 20944 13240
rect 21637 13243 21695 13249
rect 16206 13172 16212 13184
rect 14936 13144 16212 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 17770 13132 17776 13184
rect 17828 13172 17834 13184
rect 18064 13172 18092 13212
rect 21637 13209 21649 13243
rect 21683 13209 21695 13243
rect 24946 13240 24952 13252
rect 22862 13212 24952 13240
rect 21637 13203 21695 13209
rect 17828 13144 18092 13172
rect 19521 13175 19579 13181
rect 17828 13132 17834 13144
rect 19521 13141 19533 13175
rect 19567 13172 19579 13175
rect 19978 13172 19984 13184
rect 19567 13144 19984 13172
rect 19567 13141 19579 13144
rect 19521 13135 19579 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20165 13175 20223 13181
rect 20165 13141 20177 13175
rect 20211 13172 20223 13175
rect 20530 13172 20536 13184
rect 20211 13144 20536 13172
rect 20211 13141 20223 13144
rect 20165 13135 20223 13141
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 20806 13172 20812 13184
rect 20767 13144 20812 13172
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 21652 13172 21680 13203
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 25096 13212 25141 13240
rect 25096 13200 25102 13212
rect 26510 13200 26516 13252
rect 26568 13240 26574 13252
rect 26789 13243 26847 13249
rect 26789 13240 26801 13243
rect 26568 13212 26801 13240
rect 26568 13200 26574 13212
rect 26789 13209 26801 13212
rect 26835 13240 26847 13243
rect 26970 13240 26976 13252
rect 26835 13212 26976 13240
rect 26835 13209 26847 13212
rect 26789 13203 26847 13209
rect 26970 13200 26976 13212
rect 27028 13200 27034 13252
rect 27249 13243 27307 13249
rect 27249 13209 27261 13243
rect 27295 13240 27307 13243
rect 27890 13240 27896 13252
rect 27295 13212 27896 13240
rect 27295 13209 27307 13212
rect 27249 13203 27307 13209
rect 27890 13200 27896 13212
rect 27948 13200 27954 13252
rect 28810 13200 28816 13252
rect 28868 13240 28874 13252
rect 30006 13240 30012 13252
rect 28868 13212 30012 13240
rect 28868 13200 28874 13212
rect 30006 13200 30012 13212
rect 30064 13200 30070 13252
rect 23198 13172 23204 13184
rect 21652 13144 23204 13172
rect 23198 13132 23204 13144
rect 23256 13132 23262 13184
rect 23934 13172 23940 13184
rect 23895 13144 23940 13172
rect 23934 13132 23940 13144
rect 23992 13132 23998 13184
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 29546 13172 29552 13184
rect 24544 13144 29552 13172
rect 24544 13132 24550 13144
rect 29546 13132 29552 13144
rect 29604 13172 29610 13184
rect 30282 13172 30288 13184
rect 29604 13144 30288 13172
rect 29604 13132 29610 13144
rect 30282 13132 30288 13144
rect 30340 13132 30346 13184
rect 33137 13175 33195 13181
rect 33137 13141 33149 13175
rect 33183 13172 33195 13175
rect 35986 13172 35992 13184
rect 33183 13144 35992 13172
rect 33183 13141 33195 13144
rect 33137 13135 33195 13141
rect 35986 13132 35992 13144
rect 36044 13132 36050 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 9272 12940 9505 12968
rect 9272 12928 9278 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 12526 12968 12532 12980
rect 9493 12931 9551 12937
rect 12360 12940 12532 12968
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12900 1915 12903
rect 1946 12900 1952 12912
rect 1903 12872 1952 12900
rect 1903 12869 1915 12872
rect 1857 12863 1915 12869
rect 1946 12860 1952 12872
rect 2004 12860 2010 12912
rect 7282 12860 7288 12912
rect 7340 12900 7346 12912
rect 7561 12903 7619 12909
rect 7561 12900 7573 12903
rect 7340 12872 7573 12900
rect 7340 12860 7346 12872
rect 7561 12869 7573 12872
rect 7607 12869 7619 12903
rect 7561 12863 7619 12869
rect 8481 12903 8539 12909
rect 8481 12869 8493 12903
rect 8527 12900 8539 12903
rect 8846 12900 8852 12912
rect 8527 12872 8852 12900
rect 8527 12869 8539 12872
rect 8481 12863 8539 12869
rect 8846 12860 8852 12872
rect 8904 12900 8910 12912
rect 9030 12900 9036 12912
rect 8904 12872 9036 12900
rect 8904 12860 8910 12872
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 10134 12860 10140 12912
rect 10192 12900 10198 12912
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 10192 12872 11805 12900
rect 10192 12860 10198 12872
rect 11793 12869 11805 12872
rect 11839 12869 11851 12903
rect 11793 12863 11851 12869
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 3970 12832 3976 12844
rect 3931 12804 3976 12832
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 5074 12832 5080 12844
rect 5035 12804 5080 12832
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 6779 12804 7328 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 5828 12764 5856 12795
rect 3936 12736 5856 12764
rect 3936 12724 3942 12736
rect 5905 12699 5963 12705
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 7098 12696 7104 12708
rect 5951 12668 7104 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7300 12696 7328 12804
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 9180 12804 9413 12832
rect 9180 12792 9186 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 10505 12795 10563 12801
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12764 7527 12767
rect 8386 12764 8392 12776
rect 7515 12736 8392 12764
rect 7515 12733 7527 12736
rect 7469 12727 7527 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 7374 12696 7380 12708
rect 7287 12668 7380 12696
rect 7374 12656 7380 12668
rect 7432 12696 7438 12708
rect 8018 12696 8024 12708
rect 7432 12668 8024 12696
rect 7432 12656 7438 12668
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 10520 12696 10548 12795
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12360 12832 12388 12940
rect 12526 12928 12532 12940
rect 12584 12968 12590 12980
rect 13078 12968 13084 12980
rect 12584 12940 13084 12968
rect 12584 12928 12590 12940
rect 13078 12928 13084 12940
rect 13136 12968 13142 12980
rect 13136 12940 15700 12968
rect 13136 12928 13142 12940
rect 13998 12900 14004 12912
rect 13938 12872 14004 12900
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 14458 12900 14464 12912
rect 14419 12872 14464 12900
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 15672 12909 15700 12940
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 15988 12940 19334 12968
rect 15988 12928 15994 12940
rect 15657 12903 15715 12909
rect 15657 12869 15669 12903
rect 15703 12869 15715 12903
rect 17770 12900 17776 12912
rect 17731 12872 17776 12900
rect 15657 12863 15715 12869
rect 17770 12860 17776 12872
rect 17828 12860 17834 12912
rect 18322 12860 18328 12912
rect 18380 12860 18386 12912
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 12360 12804 12449 12832
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 12437 12795 12495 12801
rect 14752 12804 14933 12832
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12764 12771 12767
rect 13078 12764 13084 12776
rect 12759 12736 13084 12764
rect 12759 12733 12771 12736
rect 12713 12727 12771 12733
rect 13078 12724 13084 12736
rect 13136 12764 13142 12776
rect 14458 12764 14464 12776
rect 13136 12736 14464 12764
rect 13136 12724 13142 12736
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 14752 12696 14780 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 16908 12804 17509 12832
rect 16908 12792 16914 12804
rect 17497 12801 17509 12804
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 19306 12764 19334 12940
rect 20254 12928 20260 12980
rect 20312 12968 20318 12980
rect 25225 12971 25283 12977
rect 20312 12940 25176 12968
rect 20312 12928 20318 12940
rect 21082 12900 21088 12912
rect 19433 12872 21088 12900
rect 19433 12764 19461 12872
rect 21082 12860 21088 12872
rect 21140 12860 21146 12912
rect 23934 12900 23940 12912
rect 23506 12872 23940 12900
rect 23934 12860 23940 12872
rect 23992 12860 23998 12912
rect 20530 12832 20536 12844
rect 20491 12804 20536 12832
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 24394 12792 24400 12844
rect 24452 12832 24458 12844
rect 25148 12841 25176 12940
rect 25225 12937 25237 12971
rect 25271 12968 25283 12971
rect 27982 12968 27988 12980
rect 25271 12940 27988 12968
rect 25271 12937 25283 12940
rect 25225 12931 25283 12937
rect 27982 12928 27988 12940
rect 28040 12928 28046 12980
rect 28258 12928 28264 12980
rect 28316 12968 28322 12980
rect 34514 12968 34520 12980
rect 28316 12940 34520 12968
rect 28316 12928 28322 12940
rect 34514 12928 34520 12940
rect 34572 12928 34578 12980
rect 24489 12835 24547 12841
rect 24489 12832 24501 12835
rect 24452 12804 24501 12832
rect 24452 12792 24458 12804
rect 24489 12801 24501 12804
rect 24535 12801 24547 12835
rect 24489 12795 24547 12801
rect 25133 12835 25191 12841
rect 25133 12801 25145 12835
rect 25179 12832 25191 12835
rect 28810 12832 28816 12844
rect 25179 12804 28816 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 28810 12792 28816 12804
rect 28868 12792 28874 12844
rect 30282 12792 30288 12844
rect 30340 12832 30346 12844
rect 30745 12835 30803 12841
rect 30745 12832 30757 12835
rect 30340 12804 30757 12832
rect 30340 12792 30346 12804
rect 30745 12801 30757 12804
rect 30791 12832 30803 12835
rect 33134 12832 33140 12844
rect 30791 12804 33140 12832
rect 30791 12801 30803 12804
rect 30745 12795 30803 12801
rect 33134 12792 33140 12804
rect 33192 12792 33198 12844
rect 34790 12792 34796 12844
rect 34848 12832 34854 12844
rect 34885 12835 34943 12841
rect 34885 12832 34897 12835
rect 34848 12804 34897 12832
rect 34848 12792 34854 12804
rect 34885 12801 34897 12804
rect 34931 12801 34943 12835
rect 38102 12832 38108 12844
rect 38063 12804 38108 12832
rect 34885 12795 34943 12801
rect 38102 12792 38108 12804
rect 38160 12792 38166 12844
rect 19306 12736 19461 12764
rect 19521 12767 19579 12773
rect 19521 12733 19533 12767
rect 19567 12764 19579 12767
rect 19702 12764 19708 12776
rect 19567 12736 19708 12764
rect 19567 12733 19579 12736
rect 19521 12727 19579 12733
rect 19702 12724 19708 12736
rect 19760 12724 19766 12776
rect 21174 12724 21180 12776
rect 21232 12764 21238 12776
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 21232 12736 21281 12764
rect 21232 12724 21238 12736
rect 21269 12733 21281 12736
rect 21315 12764 21327 12767
rect 22005 12767 22063 12773
rect 22005 12764 22017 12767
rect 21315 12736 22017 12764
rect 21315 12733 21327 12736
rect 21269 12727 21327 12733
rect 22005 12733 22017 12736
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 22281 12767 22339 12773
rect 22281 12733 22293 12767
rect 22327 12764 22339 12767
rect 22370 12764 22376 12776
rect 22327 12736 22376 12764
rect 22327 12733 22339 12736
rect 22281 12727 22339 12733
rect 22370 12724 22376 12736
rect 22428 12764 22434 12776
rect 24029 12767 24087 12773
rect 22428 12736 23980 12764
rect 22428 12724 22434 12736
rect 17402 12696 17408 12708
rect 10520 12668 12572 12696
rect 14752 12668 17408 12696
rect 3786 12628 3792 12640
rect 3747 12600 3792 12628
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6788 12600 6837 12628
rect 6788 12588 6794 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9582 12628 9588 12640
rect 9456 12600 9588 12628
rect 9456 12588 9462 12600
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10008 12600 10609 12628
rect 10008 12588 10014 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 12544 12628 12572 12668
rect 17402 12656 17408 12668
rect 17460 12656 17466 12708
rect 19150 12656 19156 12708
rect 19208 12696 19214 12708
rect 21542 12696 21548 12708
rect 19208 12668 21548 12696
rect 19208 12656 19214 12668
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 23952 12696 23980 12736
rect 24029 12733 24041 12767
rect 24075 12764 24087 12767
rect 24210 12764 24216 12776
rect 24075 12736 24216 12764
rect 24075 12733 24087 12736
rect 24029 12727 24087 12733
rect 24210 12724 24216 12736
rect 24268 12764 24274 12776
rect 34146 12764 34152 12776
rect 24268 12736 34152 12764
rect 24268 12724 24274 12736
rect 34146 12724 34152 12736
rect 34204 12724 34210 12776
rect 32398 12696 32404 12708
rect 23952 12668 32404 12696
rect 32398 12656 32404 12668
rect 32456 12656 32462 12708
rect 15930 12628 15936 12640
rect 12544 12600 15936 12628
rect 10597 12591 10655 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 17420 12628 17448 12656
rect 19334 12628 19340 12640
rect 17420 12600 19340 12628
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 19702 12588 19708 12640
rect 19760 12628 19766 12640
rect 21910 12628 21916 12640
rect 19760 12600 21916 12628
rect 19760 12588 19766 12600
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 24581 12631 24639 12637
rect 24581 12597 24593 12631
rect 24627 12628 24639 12631
rect 24946 12628 24952 12640
rect 24627 12600 24952 12628
rect 24627 12597 24639 12600
rect 24581 12591 24639 12597
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 25590 12588 25596 12640
rect 25648 12628 25654 12640
rect 27338 12628 27344 12640
rect 25648 12600 27344 12628
rect 25648 12588 25654 12600
rect 27338 12588 27344 12600
rect 27396 12588 27402 12640
rect 29086 12588 29092 12640
rect 29144 12628 29150 12640
rect 30837 12631 30895 12637
rect 30837 12628 30849 12631
rect 29144 12600 30849 12628
rect 29144 12588 29150 12600
rect 30837 12597 30849 12600
rect 30883 12597 30895 12631
rect 30837 12591 30895 12597
rect 34701 12631 34759 12637
rect 34701 12597 34713 12631
rect 34747 12628 34759 12631
rect 38010 12628 38016 12640
rect 34747 12600 38016 12628
rect 34747 12597 34759 12600
rect 34701 12591 34759 12597
rect 38010 12588 38016 12600
rect 38068 12588 38074 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5074 12424 5080 12436
rect 5035 12396 5080 12424
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 6052 12396 9904 12424
rect 6052 12384 6058 12396
rect 7024 12368 7052 12396
rect 7006 12316 7012 12368
rect 7064 12316 7070 12368
rect 9876 12356 9904 12396
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10284 12396 10701 12424
rect 10284 12384 10290 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11974 12424 11980 12436
rect 11388 12396 11980 12424
rect 11388 12384 11394 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 15736 12427 15794 12433
rect 15736 12393 15748 12427
rect 15782 12424 15794 12427
rect 17954 12424 17960 12436
rect 15782 12396 17960 12424
rect 15782 12393 15794 12396
rect 15736 12387 15794 12393
rect 17954 12384 17960 12396
rect 18012 12384 18018 12436
rect 19426 12384 19432 12436
rect 19484 12384 19490 12436
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 21174 12424 21180 12436
rect 19668 12396 21180 12424
rect 19668 12384 19674 12396
rect 19444 12356 19472 12384
rect 19978 12356 19984 12368
rect 7760 12328 9720 12356
rect 9876 12328 9989 12356
rect 19444 12328 19984 12356
rect 5994 12288 6000 12300
rect 5092 12260 6000 12288
rect 5092 12229 5120 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 5500 12192 6929 12220
rect 5500 12180 5506 12192
rect 6917 12189 6929 12192
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7760 12229 7788 12328
rect 9692 12300 9720 12328
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9582 12288 9588 12300
rect 9263 12260 9588 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12288 9919 12291
rect 9961 12288 9989 12328
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 9907 12260 9989 12288
rect 9907 12257 9919 12260
rect 9861 12251 9919 12257
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10502 12288 10508 12300
rect 10100 12260 10508 12288
rect 10100 12248 10106 12260
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12526 12288 12532 12300
rect 11747 12260 12532 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 12986 12288 12992 12300
rect 12768 12260 12992 12288
rect 12768 12248 12774 12260
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 13630 12248 13636 12300
rect 13688 12288 13694 12300
rect 13725 12291 13783 12297
rect 13725 12288 13737 12291
rect 13688 12260 13737 12288
rect 13688 12248 13694 12260
rect 13725 12257 13737 12260
rect 13771 12257 13783 12291
rect 13725 12251 13783 12257
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15252 12260 15485 12288
rect 15252 12248 15258 12260
rect 15473 12257 15485 12260
rect 15519 12288 15531 12291
rect 17862 12288 17868 12300
rect 15519 12260 17868 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 17862 12248 17868 12260
rect 17920 12288 17926 12300
rect 18693 12291 18751 12297
rect 18693 12288 18705 12291
rect 17920 12260 18705 12288
rect 17920 12248 17926 12260
rect 18693 12257 18705 12260
rect 18739 12257 18751 12291
rect 18693 12251 18751 12257
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 20180 12297 20208 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 22612 12396 25544 12424
rect 22612 12384 22618 12396
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 25516 12356 25544 12396
rect 26418 12384 26424 12436
rect 26476 12424 26482 12436
rect 26970 12424 26976 12436
rect 26476 12396 26976 12424
rect 26476 12384 26482 12396
rect 26970 12384 26976 12396
rect 27028 12384 27034 12436
rect 28626 12424 28632 12436
rect 28587 12396 28632 12424
rect 28626 12384 28632 12396
rect 28684 12384 28690 12436
rect 31018 12384 31024 12436
rect 31076 12424 31082 12436
rect 34149 12427 34207 12433
rect 34149 12424 34161 12427
rect 31076 12396 34161 12424
rect 31076 12384 31082 12396
rect 34149 12393 34161 12396
rect 34195 12393 34207 12427
rect 34149 12387 34207 12393
rect 34790 12384 34796 12436
rect 34848 12424 34854 12436
rect 34977 12427 35035 12433
rect 34977 12424 34989 12427
rect 34848 12396 34989 12424
rect 34848 12384 34854 12396
rect 34977 12393 34989 12396
rect 35023 12393 35035 12427
rect 34977 12387 35035 12393
rect 25590 12356 25596 12368
rect 23164 12328 23244 12356
rect 25516 12328 25596 12356
rect 23164 12316 23170 12328
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 19484 12260 20177 12288
rect 19484 12248 19490 12260
rect 20165 12257 20177 12260
rect 20211 12257 20223 12291
rect 20165 12251 20223 12257
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7248 12192 7757 12220
rect 7248 12180 7254 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8478 12220 8484 12232
rect 8435 12192 8484 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 11514 12220 11520 12232
rect 10643 12192 11520 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17460 12192 17969 12220
rect 17460 12180 17466 12192
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 22646 12220 22652 12232
rect 21574 12192 22652 12220
rect 17957 12183 18015 12189
rect 22646 12180 22652 12192
rect 22704 12180 22710 12232
rect 23216 12229 23244 12328
rect 25590 12316 25596 12328
rect 25648 12316 25654 12368
rect 30558 12316 30564 12368
rect 30616 12356 30622 12368
rect 31570 12356 31576 12368
rect 30616 12328 31576 12356
rect 30616 12316 30622 12328
rect 31570 12316 31576 12328
rect 31628 12356 31634 12368
rect 31628 12328 31892 12356
rect 31628 12316 31634 12328
rect 24486 12248 24492 12300
rect 24544 12288 24550 12300
rect 25498 12288 25504 12300
rect 24544 12260 25504 12288
rect 24544 12248 24550 12260
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 25685 12291 25743 12297
rect 25685 12257 25697 12291
rect 25731 12288 25743 12291
rect 27154 12288 27160 12300
rect 25731 12260 27160 12288
rect 25731 12257 25743 12260
rect 25685 12251 25743 12257
rect 27154 12248 27160 12260
rect 27212 12248 27218 12300
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 31864 12297 31892 12328
rect 31849 12291 31907 12297
rect 27396 12260 31754 12288
rect 27396 12248 27402 12260
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 28350 12180 28356 12232
rect 28408 12220 28414 12232
rect 28537 12223 28595 12229
rect 28537 12220 28549 12223
rect 28408 12192 28549 12220
rect 28408 12180 28414 12192
rect 28537 12189 28549 12192
rect 28583 12189 28595 12223
rect 31726 12220 31754 12260
rect 31849 12257 31861 12291
rect 31895 12288 31907 12291
rect 31895 12260 34928 12288
rect 31895 12257 31907 12260
rect 31849 12251 31907 12257
rect 34900 12229 34928 12260
rect 34057 12223 34115 12229
rect 31726 12192 33640 12220
rect 28537 12183 28595 12189
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 5776 12124 9321 12152
rect 5776 12112 5782 12124
rect 9309 12121 9321 12124
rect 9355 12121 9367 12155
rect 9309 12115 9367 12121
rect 11698 12112 11704 12164
rect 11756 12112 11762 12164
rect 11974 12152 11980 12164
rect 11935 12124 11980 12152
rect 11974 12112 11980 12124
rect 12032 12112 12038 12164
rect 12434 12112 12440 12164
rect 12492 12112 12498 12164
rect 15654 12152 15660 12164
rect 13372 12124 15660 12152
rect 7009 12087 7067 12093
rect 7009 12053 7021 12087
rect 7055 12084 7067 12087
rect 7558 12084 7564 12096
rect 7055 12056 7564 12084
rect 7055 12053 7067 12056
rect 7009 12047 7067 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 7837 12087 7895 12093
rect 7837 12053 7849 12087
rect 7883 12084 7895 12087
rect 8294 12084 8300 12096
rect 7883 12056 8300 12084
rect 7883 12053 7895 12056
rect 7837 12047 7895 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 8444 12056 8493 12084
rect 8444 12044 8450 12056
rect 8481 12053 8493 12056
rect 8527 12053 8539 12087
rect 8481 12047 8539 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 11716 12084 11744 12112
rect 9824 12056 11744 12084
rect 11992 12084 12020 12112
rect 13372 12084 13400 12124
rect 15654 12112 15660 12124
rect 15712 12112 15718 12164
rect 16206 12112 16212 12164
rect 16264 12112 16270 12164
rect 17126 12112 17132 12164
rect 17184 12152 17190 12164
rect 17497 12155 17555 12161
rect 17497 12152 17509 12155
rect 17184 12124 17509 12152
rect 17184 12112 17190 12124
rect 17497 12121 17509 12124
rect 17543 12121 17555 12155
rect 20438 12152 20444 12164
rect 20399 12124 20444 12152
rect 17497 12115 17555 12121
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 22189 12155 22247 12161
rect 22189 12152 22201 12155
rect 22066 12124 22201 12152
rect 11992 12056 13400 12084
rect 9824 12044 9830 12056
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 18874 12084 18880 12096
rect 18380 12056 18880 12084
rect 18380 12044 18386 12056
rect 18874 12044 18880 12056
rect 18932 12084 18938 12096
rect 22066 12084 22094 12124
rect 22189 12121 22201 12124
rect 22235 12121 22247 12155
rect 22189 12115 22247 12121
rect 22462 12112 22468 12164
rect 22520 12152 22526 12164
rect 23106 12152 23112 12164
rect 22520 12124 23112 12152
rect 22520 12112 22526 12124
rect 23106 12112 23112 12124
rect 23164 12152 23170 12164
rect 25498 12152 25504 12164
rect 23164 12124 25504 12152
rect 23164 12112 23170 12124
rect 25498 12112 25504 12124
rect 25556 12112 25562 12164
rect 25958 12152 25964 12164
rect 25919 12124 25964 12152
rect 25958 12112 25964 12124
rect 26016 12112 26022 12164
rect 27709 12155 27767 12161
rect 26068 12124 26450 12152
rect 18932 12056 22094 12084
rect 23293 12087 23351 12093
rect 18932 12044 18938 12056
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 26068 12084 26096 12124
rect 27709 12121 27721 12155
rect 27755 12152 27767 12155
rect 28902 12152 28908 12164
rect 27755 12124 28908 12152
rect 27755 12121 27767 12124
rect 27709 12115 27767 12121
rect 23339 12056 26096 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 26326 12044 26332 12096
rect 26384 12084 26390 12096
rect 27724 12084 27752 12115
rect 28902 12112 28908 12124
rect 28960 12112 28966 12164
rect 30837 12155 30895 12161
rect 30837 12121 30849 12155
rect 30883 12121 30895 12155
rect 30837 12115 30895 12121
rect 30929 12155 30987 12161
rect 30929 12121 30941 12155
rect 30975 12152 30987 12155
rect 33502 12152 33508 12164
rect 30975 12124 33508 12152
rect 30975 12121 30987 12124
rect 30929 12115 30987 12121
rect 26384 12056 27752 12084
rect 26384 12044 26390 12056
rect 29730 12044 29736 12096
rect 29788 12084 29794 12096
rect 30466 12084 30472 12096
rect 29788 12056 30472 12084
rect 29788 12044 29794 12056
rect 30466 12044 30472 12056
rect 30524 12044 30530 12096
rect 30852 12084 30880 12115
rect 33502 12112 33508 12124
rect 33560 12112 33566 12164
rect 31754 12084 31760 12096
rect 30852 12056 31760 12084
rect 31754 12044 31760 12056
rect 31812 12044 31818 12096
rect 32122 12044 32128 12096
rect 32180 12084 32186 12096
rect 32674 12084 32680 12096
rect 32180 12056 32680 12084
rect 32180 12044 32186 12056
rect 32674 12044 32680 12056
rect 32732 12044 32738 12096
rect 33612 12084 33640 12192
rect 34057 12189 34069 12223
rect 34103 12189 34115 12223
rect 34057 12183 34115 12189
rect 34885 12223 34943 12229
rect 34885 12189 34897 12223
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 34072 12152 34100 12183
rect 37366 12180 37372 12232
rect 37424 12220 37430 12232
rect 38105 12223 38163 12229
rect 38105 12220 38117 12223
rect 37424 12192 38117 12220
rect 37424 12180 37430 12192
rect 38105 12189 38117 12192
rect 38151 12189 38163 12223
rect 38105 12183 38163 12189
rect 36998 12152 37004 12164
rect 34072 12124 37004 12152
rect 36998 12112 37004 12124
rect 37056 12112 37062 12164
rect 36170 12084 36176 12096
rect 33612 12056 36176 12084
rect 36170 12044 36176 12056
rect 36228 12044 36234 12096
rect 38197 12087 38255 12093
rect 38197 12053 38209 12087
rect 38243 12084 38255 12087
rect 39022 12084 39028 12096
rect 38243 12056 39028 12084
rect 38243 12053 38255 12056
rect 38197 12047 38255 12053
rect 39022 12044 39028 12056
rect 39080 12044 39086 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 9766 11880 9772 11892
rect 4172 11852 9772 11880
rect 4172 11753 4200 11852
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10134 11880 10140 11892
rect 9961 11852 10140 11880
rect 5445 11815 5503 11821
rect 5445 11781 5457 11815
rect 5491 11812 5503 11815
rect 6270 11812 6276 11824
rect 5491 11784 6276 11812
rect 5491 11781 5503 11784
rect 5445 11775 5503 11781
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 7374 11772 7380 11824
rect 7432 11812 7438 11824
rect 8386 11812 8392 11824
rect 7432 11784 7512 11812
rect 8347 11784 8392 11812
rect 7432 11772 7438 11784
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 2516 11676 2544 11707
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6917 11747 6975 11753
rect 6052 11716 6097 11744
rect 6052 11704 6058 11716
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7190 11744 7196 11756
rect 6963 11716 7196 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 7484 11744 7512 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 9674 11812 9680 11824
rect 9140 11784 9680 11812
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7484 11716 7573 11744
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 7800 11716 7880 11744
rect 7800 11704 7806 11716
rect 4614 11676 4620 11688
rect 2516 11648 4620 11676
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 5810 11676 5816 11688
rect 5399 11648 5816 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 6604 11648 7788 11676
rect 6604 11636 6610 11648
rect 6822 11568 6828 11620
rect 6880 11608 6886 11620
rect 7653 11611 7711 11617
rect 7653 11608 7665 11611
rect 6880 11580 7665 11608
rect 6880 11568 6886 11580
rect 7653 11577 7665 11580
rect 7699 11577 7711 11611
rect 7653 11571 7711 11577
rect 2314 11540 2320 11552
rect 2275 11512 2320 11540
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 3973 11543 4031 11549
rect 3973 11540 3985 11543
rect 3292 11512 3985 11540
rect 3292 11500 3298 11512
rect 3973 11509 3985 11512
rect 4019 11509 4031 11543
rect 3973 11503 4031 11509
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7190 11540 7196 11552
rect 7055 11512 7196 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 7760 11540 7788 11648
rect 7852 11608 7880 11716
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8386 11676 8392 11688
rect 8343 11648 8392 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 8536 11648 8585 11676
rect 8536 11636 8542 11648
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 9140 11608 9168 11784
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 9961 11821 9989 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 10284 11852 14780 11880
rect 10284 11840 10290 11852
rect 14752 11824 14780 11852
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 18230 11880 18236 11892
rect 15712 11852 18236 11880
rect 15712 11840 15718 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 19426 11880 19432 11892
rect 18432 11852 19432 11880
rect 9946 11815 10004 11821
rect 9946 11781 9958 11815
rect 9992 11781 10004 11815
rect 9946 11775 10004 11781
rect 10778 11772 10784 11824
rect 10836 11812 10842 11824
rect 10873 11815 10931 11821
rect 10873 11812 10885 11815
rect 10836 11784 10885 11812
rect 10836 11772 10842 11784
rect 10873 11781 10885 11784
rect 10919 11781 10931 11815
rect 10873 11775 10931 11781
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 12124 11784 13110 11812
rect 12124 11772 12130 11784
rect 14734 11772 14740 11824
rect 14792 11772 14798 11824
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 18432 11812 18460 11852
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 26970 11880 26976 11892
rect 20496 11852 26976 11880
rect 20496 11840 20502 11852
rect 26970 11840 26976 11852
rect 27028 11840 27034 11892
rect 31202 11880 31208 11892
rect 27080 11852 31208 11880
rect 14884 11784 15318 11812
rect 18340 11784 18460 11812
rect 14884 11772 14890 11784
rect 18340 11753 18368 11784
rect 18506 11772 18512 11824
rect 18564 11812 18570 11824
rect 18601 11815 18659 11821
rect 18601 11812 18613 11815
rect 18564 11784 18613 11812
rect 18564 11772 18570 11784
rect 18601 11781 18613 11784
rect 18647 11781 18659 11815
rect 18601 11775 18659 11781
rect 19058 11772 19064 11824
rect 19116 11772 19122 11824
rect 20254 11772 20260 11824
rect 20312 11812 20318 11824
rect 20349 11815 20407 11821
rect 20349 11812 20361 11815
rect 20312 11784 20361 11812
rect 20312 11772 20318 11784
rect 20349 11781 20361 11784
rect 20395 11781 20407 11815
rect 23750 11812 23756 11824
rect 23711 11784 23756 11812
rect 20349 11775 20407 11781
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 26050 11812 26056 11824
rect 24978 11784 26056 11812
rect 26050 11772 26056 11784
rect 26108 11772 26114 11824
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 10704 11716 11713 11744
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 7852 11580 9168 11608
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 9674 11608 9680 11620
rect 9364 11580 9680 11608
rect 9364 11568 9370 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 9876 11608 9904 11639
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10704 11676 10732 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 18325 11747 18383 11753
rect 18325 11713 18337 11747
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 23477 11747 23535 11753
rect 23477 11744 23489 11747
rect 22152 11716 23489 11744
rect 22152 11704 22158 11716
rect 23477 11713 23489 11716
rect 23523 11713 23535 11747
rect 23477 11707 23535 11713
rect 25498 11704 25504 11756
rect 25556 11744 25562 11756
rect 27080 11744 27108 11852
rect 31202 11840 31208 11852
rect 31260 11840 31266 11892
rect 31573 11883 31631 11889
rect 31573 11849 31585 11883
rect 31619 11880 31631 11883
rect 31662 11880 31668 11892
rect 31619 11852 31668 11880
rect 31619 11849 31631 11852
rect 31573 11843 31631 11849
rect 31662 11840 31668 11852
rect 31720 11840 31726 11892
rect 32582 11880 32588 11892
rect 32543 11852 32588 11880
rect 32582 11840 32588 11852
rect 32640 11840 32646 11892
rect 33152 11852 38148 11880
rect 27338 11772 27344 11824
rect 27396 11812 27402 11824
rect 27706 11812 27712 11824
rect 27396 11784 27712 11812
rect 27396 11772 27402 11784
rect 27706 11772 27712 11784
rect 27764 11772 27770 11824
rect 30650 11812 30656 11824
rect 28658 11784 30656 11812
rect 30650 11772 30656 11784
rect 30708 11772 30714 11824
rect 32674 11812 32680 11824
rect 30852 11784 32680 11812
rect 25556 11716 27108 11744
rect 25556 11704 25562 11716
rect 30006 11704 30012 11756
rect 30064 11744 30070 11756
rect 30852 11753 30880 11784
rect 32674 11772 32680 11784
rect 32732 11772 32738 11824
rect 30193 11747 30251 11753
rect 30193 11744 30205 11747
rect 30064 11716 30205 11744
rect 30064 11704 30070 11716
rect 30193 11713 30205 11716
rect 30239 11744 30251 11747
rect 30837 11747 30895 11753
rect 30837 11744 30849 11747
rect 30239 11716 30849 11744
rect 30239 11713 30251 11716
rect 30193 11707 30251 11713
rect 30837 11713 30849 11716
rect 30883 11713 30895 11747
rect 30837 11707 30895 11713
rect 31386 11704 31392 11756
rect 31444 11744 31450 11756
rect 31481 11747 31539 11753
rect 31481 11744 31493 11747
rect 31444 11716 31493 11744
rect 31444 11704 31450 11716
rect 31481 11713 31493 11716
rect 31527 11713 31539 11747
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 31481 11707 31539 11713
rect 31726 11716 32505 11744
rect 12342 11676 12348 11688
rect 10100 11648 10732 11676
rect 12303 11648 12348 11676
rect 10100 11636 10106 11648
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 12618 11676 12624 11688
rect 12579 11648 12624 11676
rect 12618 11636 12624 11648
rect 12676 11676 12682 11688
rect 13262 11676 13268 11688
rect 12676 11648 13268 11676
rect 12676 11636 12682 11648
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 14829 11679 14887 11685
rect 14829 11645 14841 11679
rect 14875 11676 14887 11679
rect 14875 11648 15884 11676
rect 14875 11645 14887 11648
rect 14829 11639 14887 11645
rect 10134 11608 10140 11620
rect 9876 11580 10140 11608
rect 10134 11568 10140 11580
rect 10192 11568 10198 11620
rect 10686 11568 10692 11620
rect 10744 11608 10750 11620
rect 11054 11608 11060 11620
rect 10744 11580 11060 11608
rect 10744 11568 10750 11580
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 7760 11512 11805 11540
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 13906 11540 13912 11552
rect 12124 11512 13912 11540
rect 12124 11500 12130 11512
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 14056 11512 14105 11540
rect 14056 11500 14062 11512
rect 14093 11509 14105 11512
rect 14139 11540 14151 11543
rect 14274 11540 14280 11552
rect 14139 11512 14280 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14568 11540 14596 11639
rect 15856 11608 15884 11648
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 21266 11676 21272 11688
rect 18012 11648 21272 11676
rect 18012 11636 18018 11648
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 27154 11676 27160 11688
rect 21416 11648 25268 11676
rect 27115 11648 27160 11676
rect 21416 11636 21422 11648
rect 15856 11580 18460 11608
rect 15194 11540 15200 11552
rect 14568 11512 15200 11540
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 15896 11512 16313 11540
rect 15896 11500 15902 11512
rect 16301 11509 16313 11512
rect 16347 11540 16359 11543
rect 16666 11540 16672 11552
rect 16347 11512 16672 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 18432 11540 18460 11580
rect 18690 11540 18696 11552
rect 18432 11512 18696 11540
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 24302 11540 24308 11552
rect 19760 11512 24308 11540
rect 19760 11500 19766 11512
rect 24302 11500 24308 11512
rect 24360 11500 24366 11552
rect 25240 11549 25268 11648
rect 27154 11636 27160 11648
rect 27212 11636 27218 11688
rect 27433 11679 27491 11685
rect 27433 11676 27445 11679
rect 27264 11648 27445 11676
rect 26418 11568 26424 11620
rect 26476 11608 26482 11620
rect 27062 11608 27068 11620
rect 26476 11580 27068 11608
rect 26476 11568 26482 11580
rect 27062 11568 27068 11580
rect 27120 11608 27126 11620
rect 27264 11608 27292 11648
rect 27433 11645 27445 11648
rect 27479 11645 27491 11679
rect 29178 11676 29184 11688
rect 29139 11648 29184 11676
rect 27433 11639 27491 11645
rect 29178 11636 29184 11648
rect 29236 11636 29242 11688
rect 30650 11636 30656 11688
rect 30708 11676 30714 11688
rect 31726 11676 31754 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 30708 11648 31754 11676
rect 30708 11636 30714 11648
rect 32306 11636 32312 11688
rect 32364 11676 32370 11688
rect 33152 11676 33180 11852
rect 35342 11772 35348 11824
rect 35400 11812 35406 11824
rect 36817 11815 36875 11821
rect 36817 11812 36829 11815
rect 35400 11784 36829 11812
rect 35400 11772 35406 11784
rect 36817 11781 36829 11784
rect 36863 11781 36875 11815
rect 36817 11775 36875 11781
rect 36078 11744 36084 11756
rect 36039 11716 36084 11744
rect 36078 11704 36084 11716
rect 36136 11704 36142 11756
rect 36725 11747 36783 11753
rect 36725 11713 36737 11747
rect 36771 11713 36783 11747
rect 36725 11707 36783 11713
rect 32364 11648 33180 11676
rect 32364 11636 32370 11648
rect 29730 11608 29736 11620
rect 27120 11580 27292 11608
rect 28460 11580 29736 11608
rect 27120 11568 27126 11580
rect 25225 11543 25283 11549
rect 25225 11509 25237 11543
rect 25271 11540 25283 11543
rect 28460 11540 28488 11580
rect 29730 11568 29736 11580
rect 29788 11568 29794 11620
rect 30006 11568 30012 11620
rect 30064 11608 30070 11620
rect 36740 11608 36768 11707
rect 37274 11704 37280 11756
rect 37332 11744 37338 11756
rect 38120 11753 38148 11852
rect 37461 11747 37519 11753
rect 37461 11744 37473 11747
rect 37332 11716 37473 11744
rect 37332 11704 37338 11716
rect 37461 11713 37473 11716
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 38105 11747 38163 11753
rect 38105 11713 38117 11747
rect 38151 11713 38163 11747
rect 38105 11707 38163 11713
rect 30064 11580 36768 11608
rect 37553 11611 37611 11617
rect 30064 11568 30070 11580
rect 37553 11577 37565 11611
rect 37599 11608 37611 11611
rect 38930 11608 38936 11620
rect 37599 11580 38936 11608
rect 37599 11577 37611 11580
rect 37553 11571 37611 11577
rect 38930 11568 38936 11580
rect 38988 11568 38994 11620
rect 25271 11512 28488 11540
rect 25271 11509 25283 11512
rect 25225 11503 25283 11509
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 30285 11543 30343 11549
rect 30285 11540 30297 11543
rect 30156 11512 30297 11540
rect 30156 11500 30162 11512
rect 30285 11509 30297 11512
rect 30331 11509 30343 11543
rect 30285 11503 30343 11509
rect 30834 11500 30840 11552
rect 30892 11540 30898 11552
rect 30929 11543 30987 11549
rect 30929 11540 30941 11543
rect 30892 11512 30941 11540
rect 30892 11500 30898 11512
rect 30929 11509 30941 11512
rect 30975 11509 30987 11543
rect 30929 11503 30987 11509
rect 36173 11543 36231 11549
rect 36173 11509 36185 11543
rect 36219 11540 36231 11543
rect 38102 11540 38108 11552
rect 36219 11512 38108 11540
rect 36219 11509 36231 11512
rect 36173 11503 36231 11509
rect 38102 11500 38108 11512
rect 38160 11500 38166 11552
rect 38197 11543 38255 11549
rect 38197 11509 38209 11543
rect 38243 11540 38255 11543
rect 38286 11540 38292 11552
rect 38243 11512 38292 11540
rect 38243 11509 38255 11512
rect 38197 11503 38255 11509
rect 38286 11500 38292 11512
rect 38344 11500 38350 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 3200 11308 5181 11336
rect 3200 11296 3206 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 5169 11299 5227 11305
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 7282 11336 7288 11348
rect 6871 11308 7288 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 7708 11308 9229 11336
rect 7708 11296 7714 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 10042 11336 10048 11348
rect 9217 11299 9275 11305
rect 9324 11308 10048 11336
rect 1026 11228 1032 11280
rect 1084 11268 1090 11280
rect 2317 11271 2375 11277
rect 2317 11268 2329 11271
rect 1084 11240 2329 11268
rect 1084 11228 1090 11240
rect 2317 11237 2329 11240
rect 2363 11237 2375 11271
rect 2317 11231 2375 11237
rect 3329 11271 3387 11277
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 7374 11268 7380 11280
rect 3375 11240 5212 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 5184 11212 5212 11240
rect 6748 11240 7380 11268
rect 4982 11200 4988 11212
rect 2746 11172 4988 11200
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 2746 11132 2774 11172
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 5166 11160 5172 11212
rect 5224 11160 5230 11212
rect 5810 11200 5816 11212
rect 5771 11172 5816 11200
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 2547 11104 2774 11132
rect 3237 11135 3295 11141
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 4062 11132 4068 11144
rect 3283 11104 4068 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 1596 11064 1624 11095
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 5353 11135 5411 11141
rect 4203 11104 5304 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4890 11064 4896 11076
rect 1596 11036 4896 11064
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 5074 11064 5080 11076
rect 5000 11036 5080 11064
rect 1762 10996 1768 11008
rect 1723 10968 1768 10996
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 3973 10999 4031 11005
rect 3973 10965 3985 10999
rect 4019 10996 4031 10999
rect 4614 10996 4620 11008
rect 4019 10968 4620 10996
rect 4019 10965 4031 10968
rect 3973 10959 4031 10965
rect 4614 10956 4620 10968
rect 4672 10996 4678 11008
rect 5000 10996 5028 11036
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 5276 11064 5304 11104
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 6086 11132 6092 11144
rect 5399 11104 6092 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6748 11141 6776 11240
rect 7374 11228 7380 11240
rect 7432 11228 7438 11280
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 9324 11268 9352 11308
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 11238 11336 11244 11348
rect 10192 11308 11244 11336
rect 10192 11296 10198 11308
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 11698 11336 11704 11348
rect 11563 11308 11704 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12434 11336 12440 11348
rect 11992 11308 12440 11336
rect 7800 11240 9352 11268
rect 7800 11228 7806 11240
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11200 7527 11203
rect 7650 11200 7656 11212
rect 7515 11172 7656 11200
rect 7515 11169 7527 11172
rect 7469 11163 7527 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 7834 11200 7840 11212
rect 7795 11172 7840 11200
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 11992 11209 12020 11308
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 14090 11336 14096 11348
rect 13771 11308 14096 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 18138 11336 18144 11348
rect 15528 11308 18144 11336
rect 15528 11296 15534 11308
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 23106 11336 23112 11348
rect 19306 11308 23112 11336
rect 17126 11228 17132 11280
rect 17184 11268 17190 11280
rect 19306 11268 19334 11308
rect 23106 11296 23112 11308
rect 23164 11296 23170 11348
rect 24029 11339 24087 11345
rect 24029 11305 24041 11339
rect 24075 11336 24087 11339
rect 25130 11336 25136 11348
rect 24075 11308 25136 11336
rect 24075 11305 24087 11308
rect 24029 11299 24087 11305
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 25240 11308 28994 11336
rect 17184 11240 19334 11268
rect 17184 11228 17190 11240
rect 23750 11228 23756 11280
rect 23808 11268 23814 11280
rect 25240 11268 25268 11308
rect 23808 11240 25268 11268
rect 28966 11268 28994 11308
rect 30469 11271 30527 11277
rect 30469 11268 30481 11271
rect 28966 11240 30481 11268
rect 23808 11228 23814 11240
rect 30469 11237 30481 11240
rect 30515 11237 30527 11271
rect 37458 11268 37464 11280
rect 37419 11240 37464 11268
rect 30469 11231 30527 11237
rect 37458 11228 37464 11240
rect 37516 11228 37522 11280
rect 38289 11271 38347 11277
rect 38289 11237 38301 11271
rect 38335 11268 38347 11271
rect 38654 11268 38660 11280
rect 38335 11240 38660 11268
rect 38335 11237 38347 11240
rect 38289 11231 38347 11237
rect 38654 11228 38660 11240
rect 38712 11228 38718 11280
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 9815 11172 11989 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 11977 11163 12035 11169
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 13998 11200 14004 11212
rect 12299 11172 14004 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 15470 11200 15476 11212
rect 15252 11172 15297 11200
rect 15431 11172 15476 11200
rect 15252 11160 15258 11172
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16942 11200 16948 11212
rect 16903 11172 16948 11200
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19702 11200 19708 11212
rect 19663 11172 19708 11200
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 21453 11203 21511 11209
rect 20312 11172 21036 11200
rect 20312 11160 20318 11172
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6512 11104 6745 11132
rect 6512 11092 6518 11104
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 9122 11132 9128 11144
rect 9083 11104 9128 11132
rect 6733 11095 6791 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 14274 11141 14280 11144
rect 14269 11132 14280 11141
rect 14235 11104 14280 11132
rect 14269 11095 14280 11104
rect 14274 11092 14280 11095
rect 14332 11092 14338 11144
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 15102 11132 15108 11144
rect 14415 11104 15108 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 5902 11064 5908 11076
rect 5276 11036 5908 11064
rect 5902 11024 5908 11036
rect 5960 11024 5966 11076
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 10045 11067 10103 11073
rect 7616 11036 7661 11064
rect 7616 11024 7622 11036
rect 10045 11033 10057 11067
rect 10091 11064 10103 11067
rect 10134 11064 10140 11076
rect 10091 11036 10140 11064
rect 10091 11033 10103 11036
rect 10045 11027 10103 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 11330 11064 11336 11076
rect 11270 11036 11336 11064
rect 11330 11024 11336 11036
rect 11388 11024 11394 11076
rect 12250 11024 12256 11076
rect 12308 11064 12314 11076
rect 12308 11036 12742 11064
rect 12308 11024 12314 11036
rect 14918 11024 14924 11076
rect 14976 11064 14982 11076
rect 14976 11036 15424 11064
rect 14976 11024 14982 11036
rect 4672 10968 5028 10996
rect 4672 10956 4678 10968
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 8478 10996 8484 11008
rect 6052 10968 8484 10996
rect 6052 10956 6058 10968
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 13630 10996 13636 11008
rect 9916 10968 13636 10996
rect 9916 10956 9922 10968
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 15396 10996 15424 11036
rect 15580 11036 15962 11064
rect 15580 10996 15608 11036
rect 20714 11024 20720 11076
rect 20772 11024 20778 11076
rect 21008 11064 21036 11172
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 22002 11200 22008 11212
rect 21499 11172 22008 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 22002 11160 22008 11172
rect 22060 11160 22066 11212
rect 22094 11160 22100 11212
rect 22152 11200 22158 11212
rect 22281 11203 22339 11209
rect 22281 11200 22293 11203
rect 22152 11172 22293 11200
rect 22152 11160 22158 11172
rect 22281 11169 22293 11172
rect 22327 11169 22339 11203
rect 22281 11163 22339 11169
rect 22557 11203 22615 11209
rect 22557 11169 22569 11203
rect 22603 11200 22615 11203
rect 22646 11200 22652 11212
rect 22603 11172 22652 11200
rect 22603 11169 22615 11172
rect 22557 11163 22615 11169
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 26234 11200 26240 11212
rect 26195 11172 26240 11200
rect 26234 11160 26240 11172
rect 26292 11160 26298 11212
rect 28261 11203 28319 11209
rect 28261 11169 28273 11203
rect 28307 11200 28319 11203
rect 29362 11200 29368 11212
rect 28307 11172 29368 11200
rect 28307 11169 28319 11172
rect 28261 11163 28319 11169
rect 29362 11160 29368 11172
rect 29420 11160 29426 11212
rect 29546 11160 29552 11212
rect 29604 11200 29610 11212
rect 30282 11200 30288 11212
rect 29604 11172 30288 11200
rect 29604 11160 29610 11172
rect 30282 11160 30288 11172
rect 30340 11200 30346 11212
rect 30340 11172 30420 11200
rect 30340 11160 30346 11172
rect 24578 11132 24584 11144
rect 23690 11104 24584 11132
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 24670 11092 24676 11144
rect 24728 11132 24734 11144
rect 29086 11132 29092 11144
rect 24728 11104 24992 11132
rect 24728 11092 24734 11104
rect 24762 11064 24768 11076
rect 21008 11036 22968 11064
rect 15396 10968 15608 10996
rect 18690 10956 18696 11008
rect 18748 10996 18754 11008
rect 18874 10996 18880 11008
rect 18748 10968 18880 10996
rect 18748 10956 18754 10968
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 22940 10996 22968 11036
rect 23860 11036 24768 11064
rect 23860 10996 23888 11036
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 24964 11064 24992 11104
rect 28966 11104 29092 11132
rect 26513 11067 26571 11073
rect 26513 11064 26525 11067
rect 24964 11036 26525 11064
rect 26513 11033 26525 11036
rect 26559 11033 26571 11067
rect 28966 11064 28994 11104
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 29914 11132 29920 11144
rect 29875 11104 29920 11132
rect 29914 11092 29920 11104
rect 29972 11092 29978 11144
rect 30392 11141 30420 11172
rect 30558 11160 30564 11212
rect 30616 11200 30622 11212
rect 30926 11200 30932 11212
rect 30616 11172 30932 11200
rect 30616 11160 30622 11172
rect 30926 11160 30932 11172
rect 30984 11200 30990 11212
rect 30984 11172 31524 11200
rect 30984 11160 30990 11172
rect 30377 11135 30435 11141
rect 30377 11101 30389 11135
rect 30423 11101 30435 11135
rect 30377 11095 30435 11101
rect 30466 11092 30472 11144
rect 30524 11132 30530 11144
rect 31021 11135 31079 11141
rect 31021 11132 31033 11135
rect 30524 11104 31033 11132
rect 30524 11092 30530 11104
rect 31021 11101 31033 11104
rect 31067 11101 31079 11135
rect 31496 11132 31524 11172
rect 31570 11160 31576 11212
rect 31628 11200 31634 11212
rect 32861 11203 32919 11209
rect 32861 11200 32873 11203
rect 31628 11172 32873 11200
rect 31628 11160 31634 11172
rect 32861 11169 32873 11172
rect 32907 11169 32919 11203
rect 32861 11163 32919 11169
rect 36262 11160 36268 11212
rect 36320 11160 36326 11212
rect 38102 11160 38108 11212
rect 38160 11200 38166 11212
rect 38160 11172 38700 11200
rect 38160 11160 38166 11172
rect 31665 11135 31723 11141
rect 31665 11132 31677 11135
rect 31496 11104 31677 11132
rect 31021 11095 31079 11101
rect 31665 11101 31677 11104
rect 31711 11132 31723 11135
rect 31938 11132 31944 11144
rect 31711 11104 31944 11132
rect 31711 11101 31723 11104
rect 31665 11095 31723 11101
rect 31938 11092 31944 11104
rect 31996 11092 32002 11144
rect 35894 11092 35900 11144
rect 35952 11132 35958 11144
rect 36173 11135 36231 11141
rect 36173 11132 36185 11135
rect 35952 11104 36185 11132
rect 35952 11092 35958 11104
rect 36173 11101 36185 11104
rect 36219 11101 36231 11135
rect 36280 11132 36308 11160
rect 38672 11144 38700 11172
rect 37366 11132 37372 11144
rect 36280 11104 37372 11132
rect 36173 11095 36231 11101
rect 37366 11092 37372 11104
rect 37424 11092 37430 11144
rect 38654 11092 38660 11144
rect 38712 11092 38718 11144
rect 27738 11036 28994 11064
rect 26513 11027 26571 11033
rect 31754 11024 31760 11076
rect 31812 11064 31818 11076
rect 32582 11064 32588 11076
rect 31812 11036 31857 11064
rect 32543 11036 32588 11064
rect 31812 11024 31818 11036
rect 32582 11024 32588 11036
rect 32640 11024 32646 11076
rect 32677 11067 32735 11073
rect 32677 11033 32689 11067
rect 32723 11064 32735 11067
rect 34054 11064 34060 11076
rect 32723 11036 34060 11064
rect 32723 11033 32735 11036
rect 32677 11027 32735 11033
rect 34054 11024 34060 11036
rect 34112 11024 34118 11076
rect 36265 11067 36323 11073
rect 36265 11033 36277 11067
rect 36311 11064 36323 11067
rect 36538 11064 36544 11076
rect 36311 11036 36544 11064
rect 36311 11033 36323 11036
rect 36265 11027 36323 11033
rect 36538 11024 36544 11036
rect 36596 11024 36602 11076
rect 38102 11064 38108 11076
rect 38063 11036 38108 11064
rect 38102 11024 38108 11036
rect 38160 11024 38166 11076
rect 22940 10968 23888 10996
rect 24394 10956 24400 11008
rect 24452 10996 24458 11008
rect 26326 10996 26332 11008
rect 24452 10968 26332 10996
rect 24452 10956 24458 10968
rect 26326 10956 26332 10968
rect 26384 10956 26390 11008
rect 26786 10956 26792 11008
rect 26844 10996 26850 11008
rect 29086 10996 29092 11008
rect 26844 10968 29092 10996
rect 26844 10956 26850 10968
rect 29086 10956 29092 10968
rect 29144 10956 29150 11008
rect 29730 10996 29736 11008
rect 29691 10968 29736 10996
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 31110 10996 31116 11008
rect 31071 10968 31116 10996
rect 31110 10956 31116 10968
rect 31168 10956 31174 11008
rect 32766 10956 32772 11008
rect 32824 10996 32830 11008
rect 36078 10996 36084 11008
rect 32824 10968 36084 10996
rect 32824 10956 32830 10968
rect 36078 10956 36084 10968
rect 36136 10956 36142 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 4617 10795 4675 10801
rect 2271 10764 4568 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 3326 10724 3332 10736
rect 2884 10696 3332 10724
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10625 2467 10659
rect 2774 10656 2780 10668
rect 2409 10619 2467 10625
rect 2424 10588 2452 10619
rect 2746 10616 2780 10656
rect 2832 10616 2838 10668
rect 2884 10665 2912 10696
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 4540 10724 4568 10764
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 5810 10792 5816 10804
rect 4663 10764 5816 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 7650 10792 7656 10804
rect 5951 10764 7656 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 9398 10792 9404 10804
rect 9324 10764 9404 10792
rect 5626 10724 5632 10736
rect 4540 10696 5632 10724
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 7190 10724 7196 10736
rect 7151 10696 7196 10724
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 7340 10696 7757 10724
rect 7340 10684 7346 10696
rect 7745 10693 7757 10696
rect 7791 10693 7803 10727
rect 7745 10687 7803 10693
rect 8294 10684 8300 10736
rect 8352 10724 8358 10736
rect 9324 10733 9352 10764
rect 9398 10752 9404 10764
rect 9456 10792 9462 10804
rect 10778 10792 10784 10804
rect 9456 10764 10784 10792
rect 9456 10752 9462 10764
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 14274 10792 14280 10804
rect 12032 10764 14280 10792
rect 12032 10752 12038 10764
rect 14274 10752 14280 10764
rect 14332 10792 14338 10804
rect 17126 10792 17132 10804
rect 14332 10764 17132 10792
rect 14332 10752 14338 10764
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 17862 10752 17868 10804
rect 17920 10752 17926 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 24394 10792 24400 10804
rect 21140 10764 24400 10792
rect 21140 10752 21146 10764
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 29178 10792 29184 10804
rect 24504 10764 29184 10792
rect 8389 10727 8447 10733
rect 8389 10724 8401 10727
rect 8352 10696 8401 10724
rect 8352 10684 8358 10696
rect 8389 10693 8401 10696
rect 8435 10693 8447 10727
rect 8389 10687 8447 10693
rect 9309 10727 9367 10733
rect 9309 10693 9321 10727
rect 9355 10693 9367 10727
rect 9950 10724 9956 10736
rect 9911 10696 9956 10724
rect 9309 10687 9367 10693
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 12618 10724 12624 10736
rect 11716 10696 12624 10724
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 2958 10616 2964 10668
rect 3016 10656 3022 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3016 10628 3525 10656
rect 3016 10616 3022 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 2746 10588 2774 10616
rect 2424 10560 2774 10588
rect 4540 10588 4568 10619
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 5169 10659 5227 10665
rect 5169 10656 5181 10659
rect 4672 10628 5181 10656
rect 4672 10616 4678 10628
rect 5169 10625 5181 10628
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 11716 10665 11744 10696
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 14458 10724 14464 10736
rect 14419 10696 14464 10724
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 17880 10724 17908 10752
rect 20806 10724 20812 10736
rect 17420 10696 17908 10724
rect 18906 10696 20812 10724
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5592 10628 5825 10656
rect 5592 10616 5598 10628
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 12437 10659 12495 10665
rect 12437 10652 12449 10659
rect 12483 10652 12495 10659
rect 11701 10619 11759 10625
rect 12434 10600 12440 10652
rect 12492 10600 12498 10652
rect 13814 10616 13820 10668
rect 13872 10616 13878 10668
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14424 10628 15117 10656
rect 14424 10616 14430 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 16482 10656 16488 10668
rect 15611 10628 16488 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 17420 10665 17448 10696
rect 20806 10684 20812 10696
rect 20864 10684 20870 10736
rect 24504 10733 24532 10764
rect 29178 10752 29184 10764
rect 29236 10752 29242 10804
rect 32398 10792 32404 10804
rect 29564 10764 32404 10792
rect 24489 10727 24547 10733
rect 24489 10693 24501 10727
rect 24535 10693 24547 10727
rect 24489 10687 24547 10693
rect 24946 10684 24952 10736
rect 25004 10684 25010 10736
rect 25958 10684 25964 10736
rect 26016 10724 26022 10736
rect 26786 10724 26792 10736
rect 26016 10696 26792 10724
rect 26016 10684 26022 10696
rect 26786 10684 26792 10696
rect 26844 10684 26850 10736
rect 29454 10724 29460 10736
rect 29415 10696 29460 10724
rect 29454 10684 29460 10696
rect 29512 10684 29518 10736
rect 29564 10733 29592 10764
rect 32398 10752 32404 10764
rect 32456 10752 32462 10804
rect 32582 10792 32588 10804
rect 32543 10764 32588 10792
rect 32582 10752 32588 10764
rect 32640 10752 32646 10804
rect 29549 10727 29607 10733
rect 29549 10693 29561 10727
rect 29595 10693 29607 10727
rect 29549 10687 29607 10693
rect 29914 10684 29920 10736
rect 29972 10724 29978 10736
rect 30098 10724 30104 10736
rect 29972 10696 30104 10724
rect 29972 10684 29978 10696
rect 30098 10684 30104 10696
rect 30156 10684 30162 10736
rect 30282 10684 30288 10736
rect 30340 10724 30346 10736
rect 30469 10727 30527 10733
rect 30469 10724 30481 10727
rect 30340 10696 30481 10724
rect 30340 10684 30346 10696
rect 30469 10693 30481 10696
rect 30515 10693 30527 10727
rect 30469 10687 30527 10693
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 6914 10588 6920 10600
rect 4540 10560 6920 10588
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7098 10588 7104 10600
rect 7059 10560 7104 10588
rect 7098 10548 7104 10560
rect 7156 10588 7162 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 7156 10560 8309 10588
rect 7156 10548 7162 10560
rect 8297 10557 8309 10560
rect 8343 10588 8355 10591
rect 8386 10588 8392 10600
rect 8343 10560 8392 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9732 10560 9873 10588
rect 9732 10548 9738 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 10008 10560 10149 10588
rect 10008 10548 10014 10560
rect 10137 10557 10149 10560
rect 10183 10588 10195 10591
rect 10226 10588 10232 10600
rect 10183 10560 10232 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 13170 10588 13176 10600
rect 12759 10560 13176 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 17681 10591 17739 10597
rect 13504 10560 17540 10588
rect 13504 10548 13510 10560
rect 3326 10480 3332 10532
rect 3384 10520 3390 10532
rect 3384 10492 12434 10520
rect 3384 10480 3390 10492
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 2498 10452 2504 10464
rect 1627 10424 2504 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3418 10452 3424 10464
rect 3007 10424 3424 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3602 10452 3608 10464
rect 3563 10424 3608 10452
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 5258 10452 5264 10464
rect 5219 10424 5264 10452
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 7374 10452 7380 10464
rect 5868 10424 7380 10452
rect 5868 10412 5874 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 11793 10455 11851 10461
rect 11793 10452 11805 10455
rect 9640 10424 11805 10452
rect 9640 10412 9646 10424
rect 11793 10421 11805 10424
rect 11839 10421 11851 10455
rect 12406 10452 12434 10492
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 12406 10424 14933 10452
rect 11793 10415 11851 10421
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 15654 10452 15660 10464
rect 15615 10424 15660 10452
rect 14921 10415 14979 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 17512 10452 17540 10560
rect 17681 10557 17693 10591
rect 17727 10588 17739 10591
rect 18322 10588 18328 10600
rect 17727 10560 18328 10588
rect 17727 10557 17739 10560
rect 17681 10551 17739 10557
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 18472 10560 19441 10588
rect 18472 10548 18478 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 24213 10591 24271 10597
rect 24213 10557 24225 10591
rect 24259 10588 24271 10591
rect 24259 10560 24348 10588
rect 24259 10557 24271 10560
rect 24213 10551 24271 10557
rect 18782 10480 18788 10532
rect 18840 10520 18846 10532
rect 22554 10520 22560 10532
rect 18840 10492 22560 10520
rect 18840 10480 18846 10492
rect 22554 10480 22560 10492
rect 22612 10480 22618 10532
rect 17862 10452 17868 10464
rect 17512 10424 17868 10452
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18322 10452 18328 10464
rect 18104 10424 18328 10452
rect 18104 10412 18110 10424
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 19886 10412 19892 10464
rect 19944 10452 19950 10464
rect 21910 10452 21916 10464
rect 19944 10424 21916 10452
rect 19944 10412 19950 10424
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 24320 10452 24348 10560
rect 25038 10548 25044 10600
rect 25096 10588 25102 10600
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 25096 10560 26249 10588
rect 25096 10548 25102 10560
rect 26237 10557 26249 10560
rect 26283 10557 26295 10591
rect 27154 10588 27160 10600
rect 27115 10560 27160 10588
rect 26237 10551 26295 10557
rect 27154 10548 27160 10560
rect 27212 10548 27218 10600
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10588 27491 10591
rect 28074 10588 28080 10600
rect 27479 10560 28080 10588
rect 27479 10557 27491 10560
rect 27433 10551 27491 10557
rect 28074 10548 28080 10560
rect 28132 10548 28138 10600
rect 28552 10588 28580 10642
rect 30374 10588 30380 10600
rect 28552 10560 30380 10588
rect 30374 10548 30380 10560
rect 30432 10548 30438 10600
rect 30484 10588 30512 10687
rect 30742 10684 30748 10736
rect 30800 10684 30806 10736
rect 38289 10727 38347 10733
rect 31404 10696 35480 10724
rect 30760 10656 30788 10684
rect 30929 10659 30987 10665
rect 30929 10656 30941 10659
rect 30760 10628 30941 10656
rect 30929 10625 30941 10628
rect 30975 10625 30987 10659
rect 30929 10619 30987 10625
rect 30742 10588 30748 10600
rect 30484 10560 30748 10588
rect 30742 10548 30748 10560
rect 30800 10548 30806 10600
rect 26050 10480 26056 10532
rect 26108 10520 26114 10532
rect 26108 10492 26464 10520
rect 26108 10480 26114 10492
rect 26326 10452 26332 10464
rect 24320 10424 26332 10452
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 26436 10452 26464 10492
rect 28460 10492 30236 10520
rect 28460 10452 28488 10492
rect 26436 10424 28488 10452
rect 28905 10455 28963 10461
rect 28905 10421 28917 10455
rect 28951 10452 28963 10455
rect 28994 10452 29000 10464
rect 28951 10424 29000 10452
rect 28951 10421 28963 10424
rect 28905 10415 28963 10421
rect 28994 10412 29000 10424
rect 29052 10412 29058 10464
rect 30208 10452 30236 10492
rect 30282 10480 30288 10532
rect 30340 10520 30346 10532
rect 31021 10523 31079 10529
rect 31021 10520 31033 10523
rect 30340 10492 31033 10520
rect 30340 10480 30346 10492
rect 31021 10489 31033 10492
rect 31067 10489 31079 10523
rect 31404 10520 31432 10696
rect 31573 10659 31631 10665
rect 31573 10625 31585 10659
rect 31619 10656 31631 10659
rect 32030 10656 32036 10668
rect 31619 10628 32036 10656
rect 31619 10625 31631 10628
rect 31573 10619 31631 10625
rect 32030 10616 32036 10628
rect 32088 10616 32094 10668
rect 33134 10616 33140 10668
rect 33192 10656 33198 10668
rect 35452 10665 35480 10696
rect 38289 10693 38301 10727
rect 38335 10724 38347 10727
rect 38746 10724 38752 10736
rect 38335 10696 38752 10724
rect 38335 10693 38347 10696
rect 38289 10687 38347 10693
rect 38746 10684 38752 10696
rect 38804 10684 38810 10736
rect 33229 10659 33287 10665
rect 33229 10656 33241 10659
rect 33192 10628 33241 10656
rect 33192 10616 33198 10628
rect 33229 10625 33241 10628
rect 33275 10625 33287 10659
rect 33229 10619 33287 10625
rect 35437 10659 35495 10665
rect 35437 10625 35449 10659
rect 35483 10625 35495 10659
rect 35437 10619 35495 10625
rect 35618 10616 35624 10668
rect 35676 10656 35682 10668
rect 36081 10659 36139 10665
rect 36081 10656 36093 10659
rect 35676 10628 36093 10656
rect 35676 10616 35682 10628
rect 36081 10625 36093 10628
rect 36127 10625 36139 10659
rect 36722 10656 36728 10668
rect 36683 10628 36728 10656
rect 36081 10619 36139 10625
rect 36722 10616 36728 10628
rect 36780 10616 36786 10668
rect 38102 10656 38108 10668
rect 38063 10628 38108 10656
rect 38102 10616 38108 10628
rect 38160 10616 38166 10668
rect 31662 10548 31668 10600
rect 31720 10588 31726 10600
rect 35529 10591 35587 10597
rect 35529 10588 35541 10591
rect 31720 10560 35541 10588
rect 31720 10548 31726 10560
rect 35529 10557 35541 10560
rect 35575 10557 35587 10591
rect 35529 10551 35587 10557
rect 36817 10523 36875 10529
rect 36817 10520 36829 10523
rect 31021 10483 31079 10489
rect 31128 10492 31432 10520
rect 35544 10492 36829 10520
rect 31128 10452 31156 10492
rect 35544 10464 35572 10492
rect 36817 10489 36829 10492
rect 36863 10489 36875 10523
rect 36817 10483 36875 10489
rect 30208 10424 31156 10452
rect 31202 10412 31208 10464
rect 31260 10452 31266 10464
rect 31665 10455 31723 10461
rect 31665 10452 31677 10455
rect 31260 10424 31677 10452
rect 31260 10412 31266 10424
rect 31665 10421 31677 10424
rect 31711 10421 31723 10455
rect 31665 10415 31723 10421
rect 33321 10455 33379 10461
rect 33321 10421 33333 10455
rect 33367 10452 33379 10455
rect 33410 10452 33416 10464
rect 33367 10424 33416 10452
rect 33367 10421 33379 10424
rect 33321 10415 33379 10421
rect 33410 10412 33416 10424
rect 33468 10412 33474 10464
rect 35526 10412 35532 10464
rect 35584 10412 35590 10464
rect 35894 10412 35900 10464
rect 35952 10452 35958 10464
rect 36173 10455 36231 10461
rect 36173 10452 36185 10455
rect 35952 10424 36185 10452
rect 35952 10412 35958 10424
rect 36173 10421 36185 10424
rect 36219 10421 36231 10455
rect 36173 10415 36231 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2958 10248 2964 10260
rect 1627 10220 2964 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 6270 10248 6276 10260
rect 6231 10220 6276 10248
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7466 10248 7472 10260
rect 6963 10220 7472 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 11974 10248 11980 10260
rect 7576 10220 11980 10248
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 2225 10183 2283 10189
rect 2225 10180 2237 10183
rect 1544 10152 2237 10180
rect 1544 10140 1550 10152
rect 2225 10149 2237 10152
rect 2271 10149 2283 10183
rect 2225 10143 2283 10149
rect 4341 10183 4399 10189
rect 4341 10149 4353 10183
rect 4387 10180 4399 10183
rect 7098 10180 7104 10192
rect 4387 10152 7104 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7576 10180 7604 10220
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 15654 10248 15660 10260
rect 12400 10220 15660 10248
rect 12400 10208 12406 10220
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 24118 10248 24124 10260
rect 18524 10220 24124 10248
rect 7208 10152 7604 10180
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 7208 10112 7236 10152
rect 7558 10112 7564 10124
rect 2648 10084 7236 10112
rect 7519 10084 7564 10112
rect 2648 10072 2654 10084
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2409 10047 2467 10053
rect 2409 10044 2421 10047
rect 2188 10016 2421 10044
rect 2188 10004 2194 10016
rect 2409 10013 2421 10016
rect 2455 10013 2467 10047
rect 2409 10007 2467 10013
rect 2498 10004 2504 10056
rect 2556 10044 2562 10056
rect 2866 10044 2872 10056
rect 2556 10016 2872 10044
rect 2556 10004 2562 10016
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 4264 10053 4292 10084
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8478 10112 8484 10124
rect 8439 10084 8484 10112
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10112 9827 10115
rect 9858 10112 9864 10124
rect 9815 10084 9864 10112
rect 9815 10081 9827 10084
rect 9769 10075 9827 10081
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 14277 10115 14335 10121
rect 14277 10112 14289 10115
rect 11716 10084 14289 10112
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 4982 10044 4988 10056
rect 4939 10016 4988 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 3436 9976 3464 10007
rect 4982 10004 4988 10016
rect 5040 10044 5046 10056
rect 5350 10044 5356 10056
rect 5040 10016 5356 10044
rect 5040 10004 5046 10016
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5810 10044 5816 10056
rect 5767 10016 5816 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 6270 10044 6276 10056
rect 6227 10016 6276 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 7190 10044 7196 10056
rect 6871 10016 7196 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 9456 10016 9505 10044
rect 9456 10004 9462 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11716 10053 11744 10084
rect 14277 10081 14289 10084
rect 14323 10112 14335 10115
rect 14550 10112 14556 10124
rect 14323 10084 14556 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16390 10112 16396 10124
rect 16347 10084 16396 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10112 17463 10115
rect 18414 10112 18420 10124
rect 17451 10084 18420 10112
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11572 10016 11713 10044
rect 11572 10004 11578 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13320 10016 13737 10044
rect 13320 10004 13326 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16908 10016 17141 10044
rect 16908 10004 16914 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 18524 10030 18552 10220
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 25038 10208 25044 10260
rect 25096 10248 25102 10260
rect 31202 10248 31208 10260
rect 25096 10220 31208 10248
rect 25096 10208 25102 10220
rect 31202 10208 31208 10220
rect 31260 10208 31266 10260
rect 32214 10208 32220 10260
rect 32272 10248 32278 10260
rect 32309 10251 32367 10257
rect 32309 10248 32321 10251
rect 32272 10220 32321 10248
rect 32272 10208 32278 10220
rect 32309 10217 32321 10220
rect 32355 10217 32367 10251
rect 32309 10211 32367 10217
rect 32490 10208 32496 10260
rect 32548 10248 32554 10260
rect 32953 10251 33011 10257
rect 32953 10248 32965 10251
rect 32548 10220 32965 10248
rect 32548 10208 32554 10220
rect 32953 10217 32965 10220
rect 32999 10217 33011 10251
rect 32953 10211 33011 10217
rect 33594 10208 33600 10260
rect 33652 10248 33658 10260
rect 35621 10251 35679 10257
rect 35621 10248 35633 10251
rect 33652 10220 35633 10248
rect 33652 10208 33658 10220
rect 35621 10217 35633 10220
rect 35667 10217 35679 10251
rect 35621 10211 35679 10217
rect 37550 10208 37556 10260
rect 37608 10248 37614 10260
rect 37918 10248 37924 10260
rect 37608 10220 37924 10248
rect 37608 10208 37614 10220
rect 37918 10208 37924 10220
rect 37976 10208 37982 10260
rect 18874 10180 18880 10192
rect 18835 10152 18880 10180
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 26970 10140 26976 10192
rect 27028 10180 27034 10192
rect 27028 10152 27568 10180
rect 27028 10140 27034 10152
rect 21082 10112 21088 10124
rect 21043 10084 21088 10112
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 22738 10072 22744 10124
rect 22796 10112 22802 10124
rect 22833 10115 22891 10121
rect 22833 10112 22845 10115
rect 22796 10084 22845 10112
rect 22796 10072 22802 10084
rect 22833 10081 22845 10084
rect 22879 10081 22891 10115
rect 22833 10075 22891 10081
rect 25501 10115 25559 10121
rect 25501 10081 25513 10115
rect 25547 10112 25559 10115
rect 26326 10112 26332 10124
rect 25547 10084 26332 10112
rect 25547 10081 25559 10084
rect 25501 10075 25559 10081
rect 26326 10072 26332 10084
rect 26384 10112 26390 10124
rect 27540 10121 27568 10152
rect 27614 10140 27620 10192
rect 27672 10180 27678 10192
rect 31478 10180 31484 10192
rect 27672 10152 31484 10180
rect 27672 10140 27678 10152
rect 31478 10140 31484 10152
rect 31536 10140 31542 10192
rect 31938 10140 31944 10192
rect 31996 10180 32002 10192
rect 31996 10152 33732 10180
rect 31996 10140 32002 10152
rect 27525 10115 27583 10121
rect 26384 10084 27200 10112
rect 26384 10072 26390 10084
rect 27172 10056 27200 10084
rect 27525 10081 27537 10115
rect 27571 10081 27583 10115
rect 27525 10075 27583 10081
rect 29822 10072 29828 10124
rect 29880 10112 29886 10124
rect 29917 10115 29975 10121
rect 29917 10112 29929 10115
rect 29880 10084 29929 10112
rect 29880 10072 29886 10084
rect 29917 10081 29929 10084
rect 29963 10081 29975 10115
rect 29917 10075 29975 10081
rect 30101 10115 30159 10121
rect 30101 10081 30113 10115
rect 30147 10112 30159 10115
rect 31110 10112 31116 10124
rect 30147 10084 31116 10112
rect 30147 10081 30159 10084
rect 30101 10075 30159 10081
rect 31110 10072 31116 10084
rect 31168 10072 31174 10124
rect 33597 10115 33655 10121
rect 33597 10112 33609 10115
rect 31726 10084 33609 10112
rect 20349 10047 20407 10053
rect 17129 10007 17187 10013
rect 20349 10013 20361 10047
rect 20395 10044 20407 10047
rect 20438 10044 20444 10056
rect 20395 10016 20444 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 20806 10044 20812 10056
rect 20767 10016 20812 10044
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 27154 10004 27160 10056
rect 27212 10044 27218 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 27212 10016 28733 10044
rect 27212 10004 27218 10016
rect 28721 10013 28733 10016
rect 28767 10013 28779 10047
rect 31726 10044 31754 10084
rect 33597 10081 33609 10084
rect 33643 10081 33655 10115
rect 33597 10075 33655 10081
rect 33704 10112 33732 10152
rect 34514 10140 34520 10192
rect 34572 10180 34578 10192
rect 38105 10183 38163 10189
rect 38105 10180 38117 10183
rect 34572 10152 38117 10180
rect 34572 10140 34578 10152
rect 38105 10149 38117 10152
rect 38151 10149 38163 10183
rect 38105 10143 38163 10149
rect 36262 10112 36268 10124
rect 33704 10084 36268 10112
rect 33704 10056 33732 10084
rect 36262 10072 36268 10084
rect 36320 10072 36326 10124
rect 28721 10007 28779 10013
rect 31312 10016 31754 10044
rect 6638 9976 6644 9988
rect 3436 9948 6644 9976
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 7650 9936 7656 9988
rect 7708 9976 7714 9988
rect 11974 9976 11980 9988
rect 7708 9948 7753 9976
rect 10994 9948 11376 9976
rect 11935 9948 11980 9976
rect 7708 9936 7714 9948
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 2464 9880 3249 9908
rect 2464 9868 2470 9880
rect 3237 9877 3249 9880
rect 3283 9877 3295 9911
rect 3237 9871 3295 9877
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 4985 9911 5043 9917
rect 4985 9908 4997 9911
rect 4856 9880 4997 9908
rect 4856 9868 4862 9880
rect 4985 9877 4997 9880
rect 5031 9877 5043 9911
rect 5534 9908 5540 9920
rect 5495 9880 5540 9908
rect 4985 9871 5043 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 11238 9908 11244 9920
rect 11199 9880 11244 9908
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11348 9908 11376 9948
rect 11974 9936 11980 9948
rect 12032 9976 12038 9988
rect 12250 9976 12256 9988
rect 12032 9948 12256 9976
rect 12032 9936 12038 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 14553 9979 14611 9985
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 14599 9948 14964 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 14642 9908 14648 9920
rect 11348 9880 14648 9908
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 14936 9908 14964 9948
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 25682 9976 25688 9988
rect 22310 9948 25688 9976
rect 25682 9936 25688 9948
rect 25740 9936 25746 9988
rect 25777 9979 25835 9985
rect 25777 9945 25789 9979
rect 25823 9976 25835 9979
rect 26050 9976 26056 9988
rect 25823 9948 26056 9976
rect 25823 9945 25835 9948
rect 25777 9939 25835 9945
rect 26050 9936 26056 9948
rect 26108 9936 26114 9988
rect 27430 9976 27436 9988
rect 27002 9948 27436 9976
rect 27430 9936 27436 9948
rect 27488 9936 27494 9988
rect 27890 9936 27896 9988
rect 27948 9976 27954 9988
rect 27985 9979 28043 9985
rect 27985 9976 27997 9979
rect 27948 9948 27997 9976
rect 27948 9936 27954 9948
rect 27985 9945 27997 9948
rect 28031 9945 28043 9979
rect 31312 9976 31340 10016
rect 32030 10004 32036 10056
rect 32088 10044 32094 10056
rect 32217 10047 32275 10053
rect 32217 10044 32229 10047
rect 32088 10016 32229 10044
rect 32088 10004 32094 10016
rect 32217 10013 32229 10016
rect 32263 10044 32275 10047
rect 32861 10047 32919 10053
rect 32861 10044 32873 10047
rect 32263 10016 32873 10044
rect 32263 10013 32275 10016
rect 32217 10007 32275 10013
rect 32861 10013 32873 10016
rect 32907 10044 32919 10047
rect 33318 10044 33324 10056
rect 32907 10016 33324 10044
rect 32907 10013 32919 10016
rect 32861 10007 32919 10013
rect 33318 10004 33324 10016
rect 33376 10004 33382 10056
rect 33505 10047 33563 10053
rect 33505 10013 33517 10047
rect 33551 10044 33563 10047
rect 33686 10044 33692 10056
rect 33551 10016 33692 10044
rect 33551 10013 33563 10016
rect 33505 10007 33563 10013
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 34146 10044 34152 10056
rect 34107 10016 34152 10044
rect 34146 10004 34152 10016
rect 34204 10004 34210 10056
rect 34885 10047 34943 10053
rect 34885 10013 34897 10047
rect 34931 10044 34943 10047
rect 34931 10016 35296 10044
rect 34931 10013 34943 10016
rect 34885 10007 34943 10013
rect 27985 9939 28043 9945
rect 28092 9948 31340 9976
rect 19886 9908 19892 9920
rect 14936 9880 19892 9908
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20165 9911 20223 9917
rect 20165 9877 20177 9911
rect 20211 9908 20223 9911
rect 20254 9908 20260 9920
rect 20211 9880 20260 9908
rect 20211 9877 20223 9880
rect 20165 9871 20223 9877
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 26694 9868 26700 9920
rect 26752 9908 26758 9920
rect 28092 9908 28120 9948
rect 31570 9936 31576 9988
rect 31628 9976 31634 9988
rect 31757 9979 31815 9985
rect 31757 9976 31769 9979
rect 31628 9948 31769 9976
rect 31628 9936 31634 9948
rect 31757 9945 31769 9948
rect 31803 9945 31815 9979
rect 31757 9939 31815 9945
rect 32582 9936 32588 9988
rect 32640 9976 32646 9988
rect 34977 9979 35035 9985
rect 34977 9976 34989 9979
rect 32640 9948 34989 9976
rect 32640 9936 32646 9948
rect 34977 9945 34989 9948
rect 35023 9945 35035 9979
rect 34977 9939 35035 9945
rect 26752 9880 28120 9908
rect 26752 9868 26758 9880
rect 29822 9868 29828 9920
rect 29880 9908 29886 9920
rect 33778 9908 33784 9920
rect 29880 9880 33784 9908
rect 29880 9868 29886 9880
rect 33778 9868 33784 9880
rect 33836 9868 33842 9920
rect 34241 9911 34299 9917
rect 34241 9877 34253 9911
rect 34287 9908 34299 9911
rect 34606 9908 34612 9920
rect 34287 9880 34612 9908
rect 34287 9877 34299 9880
rect 34241 9871 34299 9877
rect 34606 9868 34612 9880
rect 34664 9868 34670 9920
rect 35268 9908 35296 10016
rect 35434 10004 35440 10056
rect 35492 10044 35498 10056
rect 35529 10047 35587 10053
rect 35529 10044 35541 10047
rect 35492 10016 35541 10044
rect 35492 10004 35498 10016
rect 35529 10013 35541 10016
rect 35575 10013 35587 10047
rect 36906 10044 36912 10056
rect 36867 10016 36912 10044
rect 35529 10007 35587 10013
rect 36906 10004 36912 10016
rect 36964 10004 36970 10056
rect 37366 10044 37372 10056
rect 37327 10016 37372 10044
rect 37366 10004 37372 10016
rect 37424 10004 37430 10056
rect 38289 10047 38347 10053
rect 38289 10013 38301 10047
rect 38335 10044 38347 10047
rect 38378 10044 38384 10056
rect 38335 10016 38384 10044
rect 38335 10013 38347 10016
rect 38289 10007 38347 10013
rect 38378 10004 38384 10016
rect 38436 10004 38442 10056
rect 35802 9936 35808 9988
rect 35860 9976 35866 9988
rect 37461 9979 37519 9985
rect 37461 9976 37473 9979
rect 35860 9948 37473 9976
rect 35860 9936 35866 9948
rect 37461 9945 37473 9948
rect 37507 9945 37519 9979
rect 37461 9939 37519 9945
rect 36630 9908 36636 9920
rect 35268 9880 36636 9908
rect 36630 9868 36636 9880
rect 36688 9868 36694 9920
rect 36725 9911 36783 9917
rect 36725 9877 36737 9911
rect 36771 9908 36783 9911
rect 38102 9908 38108 9920
rect 36771 9880 38108 9908
rect 36771 9877 36783 9880
rect 36725 9871 36783 9877
rect 38102 9868 38108 9880
rect 38160 9868 38166 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 5534 9704 5540 9716
rect 1360 9676 5540 9704
rect 1360 9664 1366 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 17497 9707 17555 9713
rect 17497 9704 17509 9707
rect 6972 9676 17509 9704
rect 6972 9664 6978 9676
rect 17497 9673 17509 9676
rect 17543 9673 17555 9707
rect 26605 9707 26663 9713
rect 17497 9667 17555 9673
rect 25516 9676 26464 9704
rect 2608 9608 5580 9636
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 2608 9577 2636 9608
rect 5552 9580 5580 9608
rect 5902 9596 5908 9648
rect 5960 9596 5966 9648
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 7377 9639 7435 9645
rect 7377 9605 7389 9639
rect 7423 9636 7435 9639
rect 7742 9636 7748 9648
rect 7423 9608 7748 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 8018 9636 8024 9648
rect 7979 9608 8024 9636
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 9122 9636 9128 9648
rect 8812 9608 9128 9636
rect 8812 9596 8818 9608
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 10962 9636 10968 9648
rect 10902 9608 10968 9636
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11664 9608 11989 9636
rect 11664 9596 11670 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 12526 9596 12532 9648
rect 12584 9596 12590 9648
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13725 9639 13783 9645
rect 13725 9636 13737 9639
rect 13688 9608 13737 9636
rect 13688 9596 13694 9608
rect 13725 9605 13737 9608
rect 13771 9605 13783 9639
rect 14826 9636 14832 9648
rect 14787 9608 14832 9636
rect 13725 9599 13783 9605
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 16114 9596 16120 9648
rect 16172 9636 16178 9648
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 16172 9608 19257 9636
rect 16172 9596 16178 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 20990 9636 20996 9648
rect 20951 9608 20996 9636
rect 19245 9599 19303 9605
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 22281 9639 22339 9645
rect 22281 9605 22293 9639
rect 22327 9636 22339 9639
rect 22370 9636 22376 9648
rect 22327 9608 22376 9636
rect 22327 9605 22339 9608
rect 22281 9599 22339 9605
rect 22370 9596 22376 9608
rect 22428 9596 22434 9648
rect 22830 9596 22836 9648
rect 22888 9596 22894 9648
rect 24762 9596 24768 9648
rect 24820 9636 24826 9648
rect 25516 9636 25544 9676
rect 24820 9608 25544 9636
rect 26436 9636 26464 9676
rect 26605 9673 26617 9707
rect 26651 9704 26663 9707
rect 28442 9704 28448 9716
rect 26651 9676 27568 9704
rect 26651 9673 26663 9676
rect 26605 9667 26663 9673
rect 27433 9639 27491 9645
rect 27433 9636 27445 9639
rect 26436 9608 27445 9636
rect 24820 9596 24826 9608
rect 27433 9605 27445 9608
rect 27479 9605 27491 9639
rect 27540 9636 27568 9676
rect 27816 9676 28448 9704
rect 27706 9636 27712 9648
rect 27540 9608 27712 9636
rect 27433 9599 27491 9605
rect 27706 9596 27712 9608
rect 27764 9636 27770 9648
rect 27816 9636 27844 9676
rect 28442 9664 28448 9676
rect 28500 9664 28506 9716
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 34146 9704 34152 9716
rect 29144 9676 34152 9704
rect 29144 9664 29150 9676
rect 34146 9664 34152 9676
rect 34204 9664 34210 9716
rect 36630 9664 36636 9716
rect 36688 9704 36694 9716
rect 37090 9704 37096 9716
rect 36688 9676 37096 9704
rect 36688 9664 36694 9676
rect 37090 9664 37096 9676
rect 37148 9664 37154 9716
rect 30282 9636 30288 9648
rect 27764 9608 27844 9636
rect 30243 9608 30288 9636
rect 27764 9596 27770 9608
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 34514 9636 34520 9648
rect 32324 9608 34520 9636
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1452 9540 1777 9568
rect 1452 9528 1458 9540
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 2593 9531 2651 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 3927 9540 4537 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4525 9537 4537 9540
rect 4571 9568 4583 9571
rect 4614 9568 4620 9580
rect 4571 9540 4620 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 3896 9500 3924 9531
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4764 9540 5181 9568
rect 4764 9528 4770 9540
rect 5169 9537 5181 9540
rect 5215 9568 5227 9571
rect 5442 9568 5448 9580
rect 5215 9540 5448 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 5920 9568 5948 9596
rect 14550 9568 14556 9580
rect 5859 9540 5948 9568
rect 14511 9540 14556 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 16574 9568 16580 9580
rect 15962 9540 16580 9568
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9568 16911 9571
rect 17126 9568 17132 9580
rect 16899 9540 17132 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 17681 9531 17739 9537
rect 17788 9540 18153 9568
rect 2280 9472 3924 9500
rect 3973 9503 4031 9509
rect 2280 9460 2286 9472
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4890 9500 4896 9512
rect 4019 9472 4896 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 6733 9503 6791 9509
rect 6733 9500 6745 9503
rect 5960 9472 6745 9500
rect 5960 9460 5966 9472
rect 6733 9469 6745 9472
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7926 9500 7932 9512
rect 6880 9472 7788 9500
rect 7887 9472 7932 9500
rect 6880 9460 6886 9472
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 3878 9432 3884 9444
rect 1627 9404 3884 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 3878 9392 3884 9404
rect 3936 9392 3942 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4120 9404 6868 9432
rect 4120 9392 4126 9404
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 4614 9364 4620 9376
rect 4575 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 5261 9367 5319 9373
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 5442 9364 5448 9376
rect 5307 9336 5448 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6730 9364 6736 9376
rect 5951 9336 6736 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 6840 9364 6868 9404
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7282 9432 7288 9444
rect 6972 9404 7288 9432
rect 6972 9392 6978 9404
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 7760 9432 7788 9472
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9398 9500 9404 9512
rect 9359 9472 9404 9500
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 11698 9500 11704 9512
rect 9723 9472 11100 9500
rect 11659 9472 11704 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 8754 9432 8760 9444
rect 7760 9404 8760 9432
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 11072 9432 11100 9472
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 12434 9500 12440 9512
rect 11808 9472 12440 9500
rect 11808 9432 11836 9472
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 15838 9500 15844 9512
rect 14332 9472 15844 9500
rect 14332 9460 14338 9472
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 16206 9460 16212 9512
rect 16264 9500 16270 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 16264 9472 16313 9500
rect 16264 9460 16270 9472
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 17586 9500 17592 9512
rect 16540 9472 17592 9500
rect 16540 9460 16546 9472
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 11072 9404 11836 9432
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 17696 9432 17724 9531
rect 16816 9404 17724 9432
rect 16816 9392 16822 9404
rect 10962 9364 10968 9376
rect 6840 9336 10968 9364
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 13170 9364 13176 9376
rect 11195 9336 13176 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 14976 9336 16957 9364
rect 14976 9324 14982 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17788 9364 17816 9540
rect 18141 9537 18153 9540
rect 18187 9568 18199 9571
rect 18414 9568 18420 9580
rect 18187 9540 18420 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 18874 9528 18880 9580
rect 18932 9568 18938 9580
rect 18969 9571 19027 9577
rect 18969 9568 18981 9571
rect 18932 9540 18981 9568
rect 18932 9528 18938 9540
rect 18969 9537 18981 9540
rect 19015 9537 19027 9571
rect 18969 9531 19027 9537
rect 20346 9528 20352 9580
rect 20404 9528 20410 9580
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 22002 9568 22008 9580
rect 20864 9540 22008 9568
rect 20864 9528 20870 9540
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 26970 9568 26976 9580
rect 26266 9540 26976 9568
rect 26970 9528 26976 9540
rect 27028 9528 27034 9580
rect 27154 9568 27160 9580
rect 27115 9540 27160 9568
rect 27154 9528 27160 9540
rect 27212 9528 27218 9580
rect 29365 9571 29423 9577
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18506 9500 18512 9512
rect 18288 9472 18512 9500
rect 18288 9460 18294 9472
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 21450 9500 21456 9512
rect 19300 9472 21456 9500
rect 19300 9460 19306 9472
rect 21450 9460 21456 9472
rect 21508 9460 21514 9512
rect 22646 9500 22652 9512
rect 22066 9472 22652 9500
rect 18230 9364 18236 9376
rect 17368 9336 17816 9364
rect 18191 9336 18236 9364
rect 17368 9324 17374 9336
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19334 9364 19340 9376
rect 18932 9336 19340 9364
rect 18932 9324 18938 9336
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19610 9324 19616 9376
rect 19668 9364 19674 9376
rect 22066 9364 22094 9472
rect 22646 9460 22652 9472
rect 22704 9460 22710 9512
rect 23753 9503 23811 9509
rect 23753 9469 23765 9503
rect 23799 9500 23811 9503
rect 24670 9500 24676 9512
rect 23799 9472 24676 9500
rect 23799 9469 23811 9472
rect 23753 9463 23811 9469
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9469 24915 9503
rect 25130 9500 25136 9512
rect 25091 9472 25136 9500
rect 24857 9463 24915 9469
rect 19668 9336 22094 9364
rect 19668 9324 19674 9336
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 24762 9364 24768 9376
rect 22336 9336 24768 9364
rect 22336 9324 22342 9336
rect 24762 9324 24768 9336
rect 24820 9324 24826 9376
rect 24872 9364 24900 9463
rect 25130 9460 25136 9472
rect 25188 9460 25194 9512
rect 26142 9460 26148 9512
rect 26200 9500 26206 9512
rect 28552 9500 28580 9554
rect 29365 9537 29377 9571
rect 29411 9568 29423 9571
rect 29546 9568 29552 9580
rect 29411 9540 29552 9568
rect 29411 9537 29423 9540
rect 29365 9531 29423 9537
rect 29546 9528 29552 9540
rect 29604 9528 29610 9580
rect 32324 9577 32352 9608
rect 34514 9596 34520 9608
rect 34572 9596 34578 9648
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 32953 9571 33011 9577
rect 32953 9537 32965 9571
rect 32999 9568 33011 9571
rect 33042 9568 33048 9580
rect 32999 9540 33048 9568
rect 32999 9537 33011 9540
rect 32953 9531 33011 9537
rect 33042 9528 33048 9540
rect 33100 9528 33106 9580
rect 33134 9528 33140 9580
rect 33192 9568 33198 9580
rect 33597 9571 33655 9577
rect 33597 9568 33609 9571
rect 33192 9540 33609 9568
rect 33192 9528 33198 9540
rect 33597 9537 33609 9540
rect 33643 9568 33655 9571
rect 34146 9568 34152 9580
rect 33643 9540 34152 9568
rect 33643 9537 33655 9540
rect 33597 9531 33655 9537
rect 34146 9528 34152 9540
rect 34204 9528 34210 9580
rect 34238 9528 34244 9580
rect 34296 9568 34302 9580
rect 34296 9540 34341 9568
rect 34296 9528 34302 9540
rect 34422 9528 34428 9580
rect 34480 9568 34486 9580
rect 34885 9571 34943 9577
rect 34885 9568 34897 9571
rect 34480 9540 34897 9568
rect 34480 9528 34486 9540
rect 34885 9537 34897 9540
rect 34931 9537 34943 9571
rect 35802 9568 35808 9580
rect 35763 9540 35808 9568
rect 34885 9531 34943 9537
rect 35802 9528 35808 9540
rect 35860 9528 35866 9580
rect 36446 9568 36452 9580
rect 36407 9540 36452 9568
rect 36446 9528 36452 9540
rect 36504 9528 36510 9580
rect 36814 9528 36820 9580
rect 36872 9568 36878 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 36872 9540 37473 9568
rect 36872 9528 36878 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 37553 9571 37611 9577
rect 37553 9537 37565 9571
rect 37599 9568 37611 9571
rect 38289 9571 38347 9577
rect 38289 9568 38301 9571
rect 37599 9540 38301 9568
rect 37599 9537 37611 9540
rect 37553 9531 37611 9537
rect 38289 9537 38301 9540
rect 38335 9537 38347 9571
rect 38289 9531 38347 9537
rect 26200 9472 28580 9500
rect 26200 9460 26206 9472
rect 28626 9460 28632 9512
rect 28684 9500 28690 9512
rect 30193 9503 30251 9509
rect 28684 9472 30144 9500
rect 28684 9460 28690 9472
rect 29914 9432 29920 9444
rect 28828 9404 29920 9432
rect 26326 9364 26332 9376
rect 24872 9336 26332 9364
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 26970 9324 26976 9376
rect 27028 9364 27034 9376
rect 28828 9364 28856 9404
rect 29914 9392 29920 9404
rect 29972 9392 29978 9444
rect 27028 9336 28856 9364
rect 27028 9324 27034 9336
rect 28902 9324 28908 9376
rect 28960 9364 28966 9376
rect 29454 9364 29460 9376
rect 28960 9336 29005 9364
rect 29415 9336 29460 9364
rect 28960 9324 28966 9336
rect 29454 9324 29460 9336
rect 29512 9324 29518 9376
rect 30116 9364 30144 9472
rect 30193 9469 30205 9503
rect 30239 9469 30251 9503
rect 30193 9463 30251 9469
rect 30208 9432 30236 9463
rect 30282 9460 30288 9512
rect 30340 9500 30346 9512
rect 30469 9503 30527 9509
rect 30469 9500 30481 9503
rect 30340 9472 30481 9500
rect 30340 9460 30346 9472
rect 30469 9469 30481 9472
rect 30515 9469 30527 9503
rect 30469 9463 30527 9469
rect 31846 9460 31852 9512
rect 31904 9500 31910 9512
rect 33318 9500 33324 9512
rect 31904 9472 33324 9500
rect 31904 9460 31910 9472
rect 33318 9460 33324 9472
rect 33376 9460 33382 9512
rect 30374 9432 30380 9444
rect 30208 9404 30380 9432
rect 30374 9392 30380 9404
rect 30432 9432 30438 9444
rect 32401 9435 32459 9441
rect 32401 9432 32413 9435
rect 30432 9404 32413 9432
rect 30432 9392 30438 9404
rect 32401 9401 32413 9404
rect 32447 9401 32459 9435
rect 33686 9432 33692 9444
rect 33647 9404 33692 9432
rect 32401 9395 32459 9401
rect 33686 9392 33692 9404
rect 33744 9392 33750 9444
rect 35621 9435 35679 9441
rect 35621 9401 35633 9435
rect 35667 9432 35679 9435
rect 37366 9432 37372 9444
rect 35667 9404 37372 9432
rect 35667 9401 35679 9404
rect 35621 9395 35679 9401
rect 37366 9392 37372 9404
rect 37424 9392 37430 9444
rect 31754 9364 31760 9376
rect 30116 9336 31760 9364
rect 31754 9324 31760 9336
rect 31812 9324 31818 9376
rect 32214 9324 32220 9376
rect 32272 9364 32278 9376
rect 33045 9367 33103 9373
rect 33045 9364 33057 9367
rect 32272 9336 33057 9364
rect 32272 9324 32278 9336
rect 33045 9333 33057 9336
rect 33091 9333 33103 9367
rect 33045 9327 33103 9333
rect 33134 9324 33140 9376
rect 33192 9364 33198 9376
rect 33870 9364 33876 9376
rect 33192 9336 33876 9364
rect 33192 9324 33198 9336
rect 33870 9324 33876 9336
rect 33928 9324 33934 9376
rect 34330 9364 34336 9376
rect 34291 9336 34336 9364
rect 34330 9324 34336 9336
rect 34388 9324 34394 9376
rect 34790 9324 34796 9376
rect 34848 9364 34854 9376
rect 34977 9367 35035 9373
rect 34977 9364 34989 9367
rect 34848 9336 34989 9364
rect 34848 9324 34854 9336
rect 34977 9333 34989 9336
rect 35023 9333 35035 9367
rect 34977 9327 35035 9333
rect 36265 9367 36323 9373
rect 36265 9333 36277 9367
rect 36311 9364 36323 9367
rect 37458 9364 37464 9376
rect 36311 9336 37464 9364
rect 36311 9333 36323 9336
rect 36265 9327 36323 9333
rect 37458 9324 37464 9336
rect 37516 9324 37522 9376
rect 38010 9324 38016 9376
rect 38068 9364 38074 9376
rect 38105 9367 38163 9373
rect 38105 9364 38117 9367
rect 38068 9336 38117 9364
rect 38068 9324 38074 9336
rect 38105 9333 38117 9336
rect 38151 9333 38163 9367
rect 38105 9327 38163 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 8202 9160 8208 9172
rect 3292 9132 8208 9160
rect 3292 9120 3298 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 9324 9132 13553 9160
rect 4062 9092 4068 9104
rect 1964 9064 4068 9092
rect 1964 8965 1992 9064
rect 4062 9052 4068 9064
rect 4120 9052 4126 9104
rect 7926 9092 7932 9104
rect 4356 9064 7932 9092
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 4356 9033 4384 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 4341 9027 4399 9033
rect 2280 8996 2774 9024
rect 2280 8984 2286 8996
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 1949 8919 2007 8925
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2746 8956 2774 8996
rect 4341 8993 4353 9027
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 6178 9024 6184 9036
rect 5123 8996 6184 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6362 9024 6368 9036
rect 6323 8996 6368 9024
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 6512 8996 7573 9024
rect 6512 8984 6518 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 8168 8996 8585 9024
rect 8168 8984 8174 8996
rect 8573 8993 8585 8996
rect 8619 9024 8631 9027
rect 8938 9024 8944 9036
rect 8619 8996 8944 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 2746 8928 3249 8956
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5534 8956 5540 8968
rect 5031 8928 5540 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8956 5687 8959
rect 5994 8956 6000 8968
rect 5675 8928 6000 8956
rect 5675 8925 5687 8928
rect 5629 8919 5687 8925
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 9324 8956 9352 9132
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 17310 9160 17316 9172
rect 13541 9123 13599 9129
rect 14384 9132 17316 9160
rect 9398 9052 9404 9104
rect 9456 9052 9462 9104
rect 12250 9052 12256 9104
rect 12308 9092 12314 9104
rect 14182 9092 14188 9104
rect 12308 9064 14188 9092
rect 12308 9052 12314 9064
rect 14182 9052 14188 9064
rect 14240 9052 14246 9104
rect 9416 9024 9444 9052
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 9416 8996 10977 9024
rect 10965 8993 10977 8996
rect 11011 9024 11023 9027
rect 11790 9024 11796 9036
rect 11011 8996 11796 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 14384 9024 14412 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 19610 9160 19616 9172
rect 18288 9132 19616 9160
rect 18288 9120 18294 9132
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 22094 9160 22100 9172
rect 19720 9132 22100 9160
rect 19720 9092 19748 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22186 9120 22192 9172
rect 22244 9160 22250 9172
rect 23382 9160 23388 9172
rect 22244 9132 23388 9160
rect 22244 9120 22250 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 26050 9120 26056 9172
rect 26108 9160 26114 9172
rect 26108 9132 27752 9160
rect 26108 9120 26114 9132
rect 24026 9092 24032 9104
rect 18156 9064 19748 9092
rect 22204 9064 24032 9092
rect 12912 8996 14412 9024
rect 7064 8928 7109 8956
rect 8680 8928 9352 8956
rect 7064 8916 7070 8928
rect 2685 8891 2743 8897
rect 2685 8857 2697 8891
rect 2731 8888 2743 8891
rect 3050 8888 3056 8900
rect 2731 8860 3056 8888
rect 2731 8857 2743 8860
rect 2685 8851 2743 8857
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3252 8860 3924 8888
rect 2041 8823 2099 8829
rect 2041 8789 2053 8823
rect 2087 8820 2099 8823
rect 3252 8820 3280 8860
rect 2087 8792 3280 8820
rect 3329 8823 3387 8829
rect 2087 8789 2099 8792
rect 2041 8783 2099 8789
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 3510 8820 3516 8832
rect 3375 8792 3516 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3896 8820 3924 8860
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 6362 8888 6368 8900
rect 4028 8860 6368 8888
rect 4028 8848 4034 8860
rect 6362 8848 6368 8860
rect 6420 8848 6426 8900
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 7653 8891 7711 8897
rect 7653 8857 7665 8891
rect 7699 8888 7711 8891
rect 7834 8888 7840 8900
rect 7699 8860 7840 8888
rect 7699 8857 7711 8860
rect 7653 8851 7711 8857
rect 5534 8820 5540 8832
rect 3896 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5718 8820 5724 8832
rect 5679 8792 5724 8820
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 6472 8820 6500 8851
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 8680 8820 8708 8928
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9493 8891 9551 8897
rect 9493 8888 9505 8891
rect 9088 8860 9505 8888
rect 9088 8848 9094 8860
rect 9493 8857 9505 8860
rect 9539 8857 9551 8891
rect 9493 8851 9551 8857
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 9640 8860 9685 8888
rect 9640 8848 9646 8860
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 9950 8888 9956 8900
rect 9824 8860 9956 8888
rect 9824 8848 9830 8860
rect 9950 8848 9956 8860
rect 10008 8888 10014 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 10008 8860 10517 8888
rect 10008 8848 10014 8860
rect 10505 8857 10517 8860
rect 10551 8857 10563 8891
rect 10505 8851 10563 8857
rect 10870 8848 10876 8900
rect 10928 8888 10934 8900
rect 11241 8891 11299 8897
rect 11241 8888 11253 8891
rect 10928 8860 11253 8888
rect 10928 8848 10934 8860
rect 11241 8857 11253 8860
rect 11287 8888 11299 8891
rect 11514 8888 11520 8900
rect 11287 8860 11520 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 12250 8848 12256 8900
rect 12308 8848 12314 8900
rect 6472 8792 8708 8820
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 12912 8820 12940 8996
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 14608 8996 14657 9024
rect 14608 8984 14614 8996
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 16574 9024 16580 9036
rect 16439 8996 16580 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 16574 8984 16580 8996
rect 16632 9024 16638 9036
rect 17494 9024 17500 9036
rect 16632 8996 17500 9024
rect 16632 8984 16638 8996
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 18156 9024 18184 9064
rect 19978 9024 19984 9036
rect 17644 8996 18184 9024
rect 18248 8996 19984 9024
rect 17644 8984 17650 8996
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13412 8928 13461 8956
rect 13412 8916 13418 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 16850 8956 16856 8968
rect 16811 8928 16856 8956
rect 13449 8919 13507 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 18248 8942 18276 8996
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 20806 9024 20812 9036
rect 20767 8996 20812 9024
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 21085 9027 21143 9033
rect 21085 8993 21097 9027
rect 21131 9024 21143 9027
rect 22094 9024 22100 9036
rect 21131 8996 22100 9024
rect 21131 8993 21143 8996
rect 21085 8987 21143 8993
rect 22094 8984 22100 8996
rect 22152 8984 22158 9036
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 18877 8959 18935 8965
rect 18877 8956 18889 8959
rect 18564 8928 18889 8956
rect 18564 8916 18570 8928
rect 18877 8925 18889 8928
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 19392 8928 20177 8956
rect 19392 8916 19398 8928
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 22204 8942 22232 9064
rect 24026 9052 24032 9064
rect 24084 9052 24090 9104
rect 27724 9092 27752 9132
rect 27798 9120 27804 9172
rect 27856 9160 27862 9172
rect 28537 9163 28595 9169
rect 28537 9160 28549 9163
rect 27856 9132 28549 9160
rect 27856 9120 27862 9132
rect 28537 9129 28549 9132
rect 28583 9129 28595 9163
rect 34330 9160 34336 9172
rect 28537 9123 28595 9129
rect 29564 9132 34336 9160
rect 29454 9092 29460 9104
rect 27724 9064 29460 9092
rect 29454 9052 29460 9064
rect 29512 9052 29518 9104
rect 22830 9024 22836 9036
rect 22791 8996 22836 9024
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 23290 8984 23296 9036
rect 23348 9024 23354 9036
rect 23937 9027 23995 9033
rect 23937 9024 23949 9027
rect 23348 8996 23949 9024
rect 23348 8984 23354 8996
rect 23937 8993 23949 8996
rect 23983 8993 23995 9027
rect 24394 9024 24400 9036
rect 23937 8987 23995 8993
rect 24136 8996 24400 9024
rect 20165 8919 20223 8925
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 23845 8959 23903 8965
rect 23845 8956 23857 8959
rect 23072 8928 23857 8956
rect 23072 8916 23078 8928
rect 23845 8925 23857 8928
rect 23891 8956 23903 8959
rect 24136 8956 24164 8996
rect 24394 8984 24400 8996
rect 24452 8984 24458 9036
rect 25961 9027 26019 9033
rect 25961 8993 25973 9027
rect 26007 9024 26019 9027
rect 26326 9024 26332 9036
rect 26007 8996 26332 9024
rect 26007 8993 26019 8996
rect 25961 8987 26019 8993
rect 26326 8984 26332 8996
rect 26384 8984 26390 9036
rect 26878 8984 26884 9036
rect 26936 9024 26942 9036
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 26936 8996 27997 9024
rect 26936 8984 26942 8996
rect 27985 8993 27997 8996
rect 28031 8993 28043 9027
rect 27985 8987 28043 8993
rect 28166 8984 28172 9036
rect 28224 9024 28230 9036
rect 29564 9024 29592 9132
rect 34330 9120 34336 9132
rect 34388 9120 34394 9172
rect 35805 9163 35863 9169
rect 35805 9129 35817 9163
rect 35851 9160 35863 9163
rect 36446 9160 36452 9172
rect 35851 9132 36452 9160
rect 35851 9129 35863 9132
rect 35805 9123 35863 9129
rect 36446 9120 36452 9132
rect 36504 9120 36510 9172
rect 36998 9160 37004 9172
rect 36959 9132 37004 9160
rect 36998 9120 37004 9132
rect 37056 9120 37062 9172
rect 31110 9052 31116 9104
rect 31168 9092 31174 9104
rect 34974 9092 34980 9104
rect 31168 9064 34980 9092
rect 31168 9052 31174 9064
rect 34974 9052 34980 9064
rect 35032 9052 35038 9104
rect 36357 9095 36415 9101
rect 36357 9061 36369 9095
rect 36403 9092 36415 9095
rect 37274 9092 37280 9104
rect 36403 9064 37280 9092
rect 36403 9061 36415 9064
rect 36357 9055 36415 9061
rect 37274 9052 37280 9064
rect 37332 9052 37338 9104
rect 28224 8996 29592 9024
rect 28224 8984 28230 8996
rect 29638 8984 29644 9036
rect 29696 9024 29702 9036
rect 29917 9027 29975 9033
rect 29917 9024 29929 9027
rect 29696 8996 29929 9024
rect 29696 8984 29702 8996
rect 29917 8993 29929 8996
rect 29963 9024 29975 9027
rect 30282 9024 30288 9036
rect 29963 8996 30288 9024
rect 29963 8993 29975 8996
rect 29917 8987 29975 8993
rect 30282 8984 30288 8996
rect 30340 8984 30346 9036
rect 30742 9024 30748 9036
rect 30703 8996 30748 9024
rect 30742 8984 30748 8996
rect 30800 8984 30806 9036
rect 31754 9024 31760 9036
rect 30852 8996 31760 9024
rect 25317 8959 25375 8965
rect 25317 8956 25329 8959
rect 23891 8928 24164 8956
rect 24228 8928 25329 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 12989 8891 13047 8897
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13078 8888 13084 8900
rect 13035 8860 13084 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13078 8848 13084 8860
rect 13136 8888 13142 8900
rect 13722 8888 13728 8900
rect 13136 8860 13728 8888
rect 13136 8848 13142 8860
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 14550 8848 14556 8900
rect 14608 8888 14614 8900
rect 14921 8891 14979 8897
rect 14921 8888 14933 8891
rect 14608 8860 14933 8888
rect 14608 8848 14614 8860
rect 14921 8857 14933 8860
rect 14967 8857 14979 8891
rect 14921 8851 14979 8857
rect 15010 8848 15016 8900
rect 15068 8888 15074 8900
rect 17126 8888 17132 8900
rect 15068 8860 15410 8888
rect 17087 8860 17132 8888
rect 15068 8848 15074 8860
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 19426 8888 19432 8900
rect 19387 8860 19432 8888
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 24228 8888 24256 8928
rect 25317 8925 25329 8928
rect 25363 8925 25375 8959
rect 25317 8919 25375 8925
rect 27338 8916 27344 8968
rect 27396 8916 27402 8968
rect 28442 8956 28448 8968
rect 28403 8928 28448 8956
rect 28442 8916 28448 8928
rect 28500 8916 28506 8968
rect 28994 8916 29000 8968
rect 29052 8916 29058 8968
rect 23860 8860 24256 8888
rect 24581 8891 24639 8897
rect 23860 8832 23888 8860
rect 24581 8857 24593 8891
rect 24627 8888 24639 8891
rect 24854 8888 24860 8900
rect 24627 8860 24860 8888
rect 24627 8857 24639 8860
rect 24581 8851 24639 8857
rect 24854 8848 24860 8860
rect 24912 8848 24918 8900
rect 26237 8891 26295 8897
rect 26237 8857 26249 8891
rect 26283 8857 26295 8891
rect 26237 8851 26295 8857
rect 8812 8792 12940 8820
rect 8812 8780 8818 8792
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 21174 8820 21180 8832
rect 13228 8792 21180 8820
rect 13228 8780 13234 8792
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 22002 8780 22008 8832
rect 22060 8820 22066 8832
rect 23842 8820 23848 8832
rect 22060 8792 23848 8820
rect 22060 8780 22066 8792
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 24946 8780 24952 8832
rect 25004 8820 25010 8832
rect 25590 8820 25596 8832
rect 25004 8792 25596 8820
rect 25004 8780 25010 8792
rect 25590 8780 25596 8792
rect 25648 8780 25654 8832
rect 26252 8820 26280 8851
rect 27706 8848 27712 8900
rect 27764 8888 27770 8900
rect 29012 8888 29040 8916
rect 27764 8860 29040 8888
rect 30009 8891 30067 8897
rect 27764 8848 27770 8860
rect 30009 8857 30021 8891
rect 30055 8888 30067 8891
rect 30852 8888 30880 8996
rect 31754 8984 31760 8996
rect 31812 8984 31818 9036
rect 31846 8984 31852 9036
rect 31904 9024 31910 9036
rect 31904 8996 31949 9024
rect 31904 8984 31910 8996
rect 34238 8984 34244 9036
rect 34296 9024 34302 9036
rect 34296 8996 34928 9024
rect 34296 8984 34302 8996
rect 32585 8959 32643 8965
rect 32585 8925 32597 8959
rect 32631 8952 32643 8959
rect 32766 8952 32772 8968
rect 32631 8925 32772 8952
rect 32585 8924 32772 8925
rect 32585 8919 32643 8924
rect 32766 8916 32772 8924
rect 32824 8916 32830 8968
rect 33226 8956 33232 8968
rect 33187 8928 33232 8956
rect 33226 8916 33232 8928
rect 33284 8916 33290 8968
rect 33321 8959 33379 8965
rect 33321 8925 33333 8959
rect 33367 8956 33379 8959
rect 33502 8956 33508 8968
rect 33367 8928 33508 8956
rect 33367 8925 33379 8928
rect 33321 8919 33379 8925
rect 33502 8916 33508 8928
rect 33560 8916 33566 8968
rect 33870 8956 33876 8968
rect 33831 8928 33876 8956
rect 33870 8916 33876 8928
rect 33928 8956 33934 8968
rect 34514 8956 34520 8968
rect 33928 8928 34520 8956
rect 33928 8916 33934 8928
rect 34514 8916 34520 8928
rect 34572 8916 34578 8968
rect 34900 8965 34928 8996
rect 34885 8959 34943 8965
rect 34885 8925 34897 8959
rect 34931 8956 34943 8959
rect 35710 8956 35716 8968
rect 34931 8928 35388 8956
rect 35671 8928 35716 8956
rect 34931 8925 34943 8928
rect 34885 8919 34943 8925
rect 30055 8860 30880 8888
rect 31481 8891 31539 8897
rect 30055 8857 30067 8860
rect 30009 8851 30067 8857
rect 31481 8857 31493 8891
rect 31527 8857 31539 8891
rect 31481 8851 31539 8857
rect 31573 8891 31631 8897
rect 31573 8857 31585 8891
rect 31619 8888 31631 8891
rect 31619 8860 32996 8888
rect 31619 8857 31631 8860
rect 31573 8851 31631 8857
rect 26878 8820 26884 8832
rect 26252 8792 26884 8820
rect 26878 8780 26884 8792
rect 26936 8780 26942 8832
rect 27062 8780 27068 8832
rect 27120 8820 27126 8832
rect 28994 8820 29000 8832
rect 27120 8792 29000 8820
rect 27120 8780 27126 8792
rect 28994 8780 29000 8792
rect 29052 8780 29058 8832
rect 30466 8780 30472 8832
rect 30524 8820 30530 8832
rect 31496 8820 31524 8851
rect 30524 8792 31524 8820
rect 30524 8780 30530 8792
rect 31662 8780 31668 8832
rect 31720 8820 31726 8832
rect 32677 8823 32735 8829
rect 32677 8820 32689 8823
rect 31720 8792 32689 8820
rect 31720 8780 31726 8792
rect 32677 8789 32689 8792
rect 32723 8789 32735 8823
rect 32968 8820 32996 8860
rect 33134 8848 33140 8900
rect 33192 8888 33198 8900
rect 33965 8891 34023 8897
rect 33965 8888 33977 8891
rect 33192 8860 33977 8888
rect 33192 8848 33198 8860
rect 33965 8857 33977 8860
rect 34011 8857 34023 8891
rect 35250 8888 35256 8900
rect 33965 8851 34023 8857
rect 34716 8860 35256 8888
rect 34716 8820 34744 8860
rect 35250 8848 35256 8860
rect 35308 8848 35314 8900
rect 32968 8792 34744 8820
rect 32677 8783 32735 8789
rect 34790 8780 34796 8832
rect 34848 8820 34854 8832
rect 34977 8823 35035 8829
rect 34977 8820 34989 8823
rect 34848 8792 34989 8820
rect 34848 8780 34854 8792
rect 34977 8789 34989 8792
rect 35023 8789 35035 8823
rect 35360 8820 35388 8928
rect 35710 8916 35716 8928
rect 35768 8916 35774 8968
rect 36538 8956 36544 8968
rect 36499 8928 36544 8956
rect 36538 8916 36544 8928
rect 36596 8916 36602 8968
rect 37185 8959 37243 8965
rect 37185 8925 37197 8959
rect 37231 8925 37243 8959
rect 37185 8919 37243 8925
rect 35802 8848 35808 8900
rect 35860 8888 35866 8900
rect 37200 8888 37228 8919
rect 37826 8916 37832 8968
rect 37884 8956 37890 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 37884 8928 38025 8956
rect 37884 8916 37890 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 35860 8860 37228 8888
rect 35860 8848 35866 8860
rect 37182 8820 37188 8832
rect 35360 8792 37188 8820
rect 34977 8783 35035 8789
rect 37182 8780 37188 8792
rect 37240 8820 37246 8832
rect 37826 8820 37832 8832
rect 37240 8792 37832 8820
rect 37240 8780 37246 8792
rect 37826 8780 37832 8792
rect 37884 8780 37890 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 4764 8588 8064 8616
rect 4764 8576 4770 8588
rect 5442 8557 5448 8560
rect 5438 8511 5448 8557
rect 5500 8548 5506 8560
rect 6822 8557 6828 8560
rect 5500 8520 5538 8548
rect 5442 8508 5448 8511
rect 5500 8508 5506 8520
rect 6818 8511 6828 8557
rect 6880 8548 6886 8560
rect 8036 8557 8064 8588
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 9766 8616 9772 8628
rect 8168 8588 9772 8616
rect 8168 8576 8174 8588
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 11238 8616 11244 8628
rect 9876 8588 11244 8616
rect 8021 8551 8079 8557
rect 6880 8520 6918 8548
rect 6822 8508 6828 8511
rect 6880 8508 6886 8520
rect 8021 8517 8033 8551
rect 8067 8517 8079 8551
rect 8021 8511 8079 8517
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 8628 8520 8953 8548
rect 8628 8508 8634 8520
rect 8941 8517 8953 8520
rect 8987 8517 8999 8551
rect 8941 8511 8999 8517
rect 9677 8551 9735 8557
rect 9677 8517 9689 8551
rect 9723 8548 9735 8551
rect 9876 8548 9904 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 12434 8616 12440 8628
rect 11624 8588 12440 8616
rect 11624 8548 11652 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14274 8616 14280 8628
rect 12636 8588 14280 8616
rect 9723 8520 9904 8548
rect 10902 8520 11652 8548
rect 9723 8517 9735 8520
rect 9677 8511 9735 8517
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 12526 8548 12532 8560
rect 11940 8520 12532 8548
rect 11940 8508 11946 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 12636 8557 12664 8588
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 16574 8616 16580 8628
rect 14844 8588 16580 8616
rect 12621 8551 12679 8557
rect 12621 8517 12633 8551
rect 12667 8517 12679 8551
rect 12621 8511 12679 8517
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 14844 8557 14872 8588
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 16908 8588 19104 8616
rect 16908 8576 16914 8588
rect 14829 8551 14887 8557
rect 12952 8520 13110 8548
rect 12952 8508 12958 8520
rect 14829 8517 14841 8551
rect 14875 8517 14887 8551
rect 16298 8548 16304 8560
rect 16054 8520 16304 8548
rect 14829 8511 14887 8517
rect 16298 8508 16304 8520
rect 16356 8508 16362 8560
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 16448 8520 17141 8548
rect 16448 8508 16454 8520
rect 17129 8517 17141 8520
rect 17175 8517 17187 8551
rect 18966 8548 18972 8560
rect 18354 8520 18972 8548
rect 17129 8511 17187 8517
rect 18966 8508 18972 8520
rect 19024 8508 19030 8560
rect 19076 8548 19104 8588
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 24762 8616 24768 8628
rect 19484 8588 24768 8616
rect 19484 8576 19490 8588
rect 19334 8548 19340 8560
rect 19076 8520 19340 8548
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 1811 8452 2421 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 2409 8449 2421 8452
rect 2455 8480 2467 8483
rect 2590 8480 2596 8492
rect 2455 8452 2596 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 3234 8480 3240 8492
rect 3195 8452 3240 8480
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4246 8480 4252 8492
rect 3743 8452 4252 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 4356 8412 4384 8443
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 9398 8480 9404 8492
rect 9359 8452 9404 8480
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11664 8452 11713 8480
rect 11664 8440 11670 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 19076 8489 19104 8520
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 21726 8548 21732 8560
rect 20562 8520 21732 8548
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 23768 8557 23796 8588
rect 24762 8576 24768 8588
rect 24820 8576 24826 8628
rect 32398 8616 32404 8628
rect 25976 8588 27614 8616
rect 23753 8551 23811 8557
rect 23753 8517 23765 8551
rect 23799 8517 23811 8551
rect 25976 8548 26004 8588
rect 27062 8548 27068 8560
rect 25714 8520 26004 8548
rect 26620 8520 27068 8548
rect 23753 8511 23811 8517
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 11848 8452 12357 8480
rect 11848 8440 11854 8452
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21968 8452 22017 8480
rect 21968 8440 21974 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 26620 8489 26648 8520
rect 27062 8508 27068 8520
rect 27120 8508 27126 8560
rect 27338 8508 27344 8560
rect 27396 8548 27402 8560
rect 27433 8551 27491 8557
rect 27433 8548 27445 8551
rect 27396 8520 27445 8548
rect 27396 8508 27402 8520
rect 27433 8517 27445 8520
rect 27479 8517 27491 8551
rect 27586 8548 27614 8588
rect 27816 8588 31248 8616
rect 32359 8588 32404 8616
rect 27816 8548 27844 8588
rect 27586 8520 27844 8548
rect 29549 8551 29607 8557
rect 27433 8511 27491 8517
rect 29549 8517 29561 8551
rect 29595 8548 29607 8551
rect 30469 8551 30527 8557
rect 30469 8548 30481 8551
rect 29595 8520 30481 8548
rect 29595 8517 29607 8520
rect 29549 8511 29607 8517
rect 30469 8517 30481 8520
rect 30515 8517 30527 8551
rect 30469 8511 30527 8517
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 23900 8452 24225 8480
rect 23900 8440 23906 8452
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 26605 8483 26663 8489
rect 26605 8449 26617 8483
rect 26651 8449 26663 8483
rect 28566 8452 29132 8480
rect 26605 8443 26663 8449
rect 2924 8384 4384 8412
rect 4433 8415 4491 8421
rect 2924 8372 2930 8384
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 5353 8415 5411 8421
rect 5353 8412 5365 8415
rect 4479 8384 5365 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 5353 8381 5365 8384
rect 5399 8381 5411 8415
rect 6380 8412 6408 8440
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 6380 8384 6745 8412
rect 5353 8375 5411 8381
rect 6733 8381 6745 8384
rect 6779 8412 6791 8415
rect 6822 8412 6828 8424
rect 6779 8384 6828 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7006 8412 7012 8424
rect 6967 8384 7012 8412
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 8846 8412 8852 8424
rect 7975 8384 8852 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9766 8412 9772 8424
rect 8956 8384 9772 8412
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 1946 8344 1952 8356
rect 1903 8316 1952 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3234 8344 3240 8356
rect 3099 8316 3240 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 6914 8344 6920 8356
rect 5951 8316 6920 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 7650 8344 7656 8356
rect 7432 8316 7656 8344
rect 7432 8304 7438 8316
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8956 8344 8984 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 10134 8372 10140 8424
rect 10192 8412 10198 8424
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 10192 8384 11161 8412
rect 10192 8372 10198 8384
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 16850 8412 16856 8424
rect 14599 8384 16856 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 18414 8412 18420 8424
rect 17184 8384 18420 8412
rect 17184 8372 17190 8384
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 18601 8415 18659 8421
rect 18601 8381 18613 8415
rect 18647 8412 18659 8415
rect 21082 8412 21088 8424
rect 18647 8384 20392 8412
rect 21043 8384 21088 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 14090 8344 14096 8356
rect 8260 8316 8984 8344
rect 14051 8316 14096 8344
rect 8260 8304 8266 8316
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 16172 8316 16313 8344
rect 16172 8304 16178 8316
rect 16301 8313 16313 8316
rect 16347 8313 16359 8347
rect 20364 8344 20392 8384
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 21174 8372 21180 8424
rect 21232 8412 21238 8424
rect 22830 8412 22836 8424
rect 21232 8384 22836 8412
rect 21232 8372 21238 8384
rect 22830 8372 22836 8384
rect 22888 8372 22894 8424
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 24044 8384 24501 8412
rect 24044 8344 24072 8384
rect 24489 8381 24501 8384
rect 24535 8412 24547 8415
rect 24946 8412 24952 8424
rect 24535 8384 24952 8412
rect 24535 8381 24547 8384
rect 24489 8375 24547 8381
rect 24946 8372 24952 8384
rect 25004 8372 25010 8424
rect 25130 8372 25136 8424
rect 25188 8412 25194 8424
rect 27154 8412 27160 8424
rect 25188 8384 26556 8412
rect 27115 8384 27160 8412
rect 25188 8372 25194 8384
rect 20364 8316 24072 8344
rect 16301 8307 16359 8313
rect 25498 8304 25504 8356
rect 25556 8344 25562 8356
rect 25774 8344 25780 8356
rect 25556 8316 25780 8344
rect 25556 8304 25562 8316
rect 25774 8304 25780 8316
rect 25832 8344 25838 8356
rect 25961 8347 26019 8353
rect 25961 8344 25973 8347
rect 25832 8316 25973 8344
rect 25832 8304 25838 8316
rect 25961 8313 25973 8316
rect 26007 8313 26019 8347
rect 25961 8307 26019 8313
rect 26326 8304 26332 8356
rect 26384 8344 26390 8356
rect 26421 8347 26479 8353
rect 26421 8344 26433 8347
rect 26384 8316 26433 8344
rect 26384 8304 26390 8316
rect 26421 8313 26433 8316
rect 26467 8313 26479 8347
rect 26528 8344 26556 8384
rect 27154 8372 27160 8384
rect 27212 8372 27218 8424
rect 27982 8412 27988 8424
rect 27264 8384 27988 8412
rect 27264 8344 27292 8384
rect 27982 8372 27988 8384
rect 28040 8412 28046 8424
rect 28905 8415 28963 8421
rect 28905 8412 28917 8415
rect 28040 8384 28917 8412
rect 28040 8372 28046 8384
rect 28905 8381 28917 8384
rect 28951 8381 28963 8415
rect 28905 8375 28963 8381
rect 26528 8316 27292 8344
rect 29104 8344 29132 8452
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 29362 8480 29368 8492
rect 29236 8452 29368 8480
rect 29236 8440 29242 8452
rect 29362 8440 29368 8452
rect 29420 8480 29426 8492
rect 29457 8483 29515 8489
rect 29457 8480 29469 8483
rect 29420 8452 29469 8480
rect 29420 8440 29426 8452
rect 29457 8449 29469 8452
rect 29503 8449 29515 8483
rect 31220 8480 31248 8588
rect 32398 8576 32404 8588
rect 32456 8576 32462 8628
rect 32950 8576 32956 8628
rect 33008 8616 33014 8628
rect 34974 8616 34980 8628
rect 33008 8588 33180 8616
rect 34935 8588 34980 8616
rect 33008 8576 33014 8588
rect 32030 8508 32036 8560
rect 32088 8548 32094 8560
rect 33045 8551 33103 8557
rect 33045 8548 33057 8551
rect 32088 8520 33057 8548
rect 32088 8508 32094 8520
rect 33045 8517 33057 8520
rect 33091 8517 33103 8551
rect 33152 8548 33180 8588
rect 34974 8576 34980 8588
rect 35032 8576 35038 8628
rect 35621 8551 35679 8557
rect 35621 8548 35633 8551
rect 33152 8520 35633 8548
rect 33045 8511 33103 8517
rect 35621 8517 35633 8520
rect 35667 8517 35679 8551
rect 36262 8548 36268 8560
rect 35621 8511 35679 8517
rect 35728 8520 36268 8548
rect 32309 8483 32367 8489
rect 31220 8452 32260 8480
rect 29457 8443 29515 8449
rect 30374 8412 30380 8424
rect 30335 8384 30380 8412
rect 30374 8372 30380 8384
rect 30432 8372 30438 8424
rect 30558 8372 30564 8424
rect 30616 8412 30622 8424
rect 30653 8415 30711 8421
rect 30653 8412 30665 8415
rect 30616 8384 30665 8412
rect 30616 8372 30622 8384
rect 30653 8381 30665 8384
rect 30699 8381 30711 8415
rect 30653 8375 30711 8381
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 31662 8412 31668 8424
rect 31076 8384 31668 8412
rect 31076 8372 31082 8384
rect 31662 8372 31668 8384
rect 31720 8372 31726 8424
rect 32232 8412 32260 8452
rect 32309 8449 32321 8483
rect 32355 8480 32367 8483
rect 32674 8480 32680 8492
rect 32355 8452 32680 8480
rect 32355 8449 32367 8452
rect 32309 8443 32367 8449
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8480 33011 8483
rect 33226 8480 33232 8492
rect 32999 8452 33232 8480
rect 32999 8449 33011 8452
rect 32953 8443 33011 8449
rect 33226 8440 33232 8452
rect 33284 8480 33290 8492
rect 33597 8483 33655 8489
rect 33597 8480 33609 8483
rect 33284 8452 33609 8480
rect 33284 8440 33290 8452
rect 33597 8449 33609 8452
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 34241 8483 34299 8489
rect 34241 8449 34253 8483
rect 34287 8480 34299 8483
rect 34514 8480 34520 8492
rect 34287 8452 34520 8480
rect 34287 8449 34299 8452
rect 34241 8443 34299 8449
rect 34514 8440 34520 8452
rect 34572 8480 34578 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34572 8452 34897 8480
rect 34572 8440 34578 8452
rect 34885 8449 34897 8452
rect 34931 8480 34943 8483
rect 35434 8480 35440 8492
rect 34931 8452 35440 8480
rect 34931 8449 34943 8452
rect 34885 8443 34943 8449
rect 35434 8440 35440 8452
rect 35492 8440 35498 8492
rect 35529 8483 35587 8489
rect 35529 8449 35541 8483
rect 35575 8480 35587 8483
rect 35728 8480 35756 8520
rect 36262 8508 36268 8520
rect 36320 8508 36326 8560
rect 36170 8480 36176 8492
rect 35575 8452 35756 8480
rect 36131 8452 36176 8480
rect 35575 8449 35587 8452
rect 35529 8443 35587 8449
rect 36170 8440 36176 8452
rect 36228 8440 36234 8492
rect 38010 8480 38016 8492
rect 37971 8452 38016 8480
rect 38010 8440 38016 8452
rect 38068 8440 38074 8492
rect 35618 8412 35624 8424
rect 32232 8384 35624 8412
rect 35618 8372 35624 8384
rect 35676 8372 35682 8424
rect 30926 8344 30932 8356
rect 29104 8316 30932 8344
rect 26421 8307 26479 8313
rect 30926 8304 30932 8316
rect 30984 8304 30990 8356
rect 33689 8347 33747 8353
rect 33689 8344 33701 8347
rect 31036 8316 33701 8344
rect 2501 8279 2559 8285
rect 2501 8245 2513 8279
rect 2547 8276 2559 8279
rect 3694 8276 3700 8288
rect 2547 8248 3700 8276
rect 2547 8245 2559 8248
rect 2501 8239 2559 8245
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 3789 8279 3847 8285
rect 3789 8245 3801 8279
rect 3835 8276 3847 8279
rect 4062 8276 4068 8288
rect 3835 8248 4068 8276
rect 3835 8245 3847 8248
rect 3789 8239 3847 8245
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 9674 8276 9680 8288
rect 6420 8248 9680 8276
rect 6420 8236 6426 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 11793 8279 11851 8285
rect 11793 8245 11805 8279
rect 11839 8276 11851 8279
rect 11882 8276 11888 8288
rect 11839 8248 11888 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 14550 8276 14556 8288
rect 12308 8248 14556 8276
rect 12308 8236 12314 8248
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 16758 8236 16764 8288
rect 16816 8276 16822 8288
rect 19058 8276 19064 8288
rect 16816 8248 19064 8276
rect 16816 8236 16822 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 19318 8279 19376 8285
rect 19318 8276 19330 8279
rect 19208 8248 19330 8276
rect 19208 8236 19214 8248
rect 19318 8245 19330 8248
rect 19364 8245 19376 8279
rect 19318 8239 19376 8245
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 21082 8276 21088 8288
rect 19484 8248 21088 8276
rect 19484 8236 19490 8248
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 24946 8236 24952 8288
rect 25004 8276 25010 8288
rect 25866 8276 25872 8288
rect 25004 8248 25872 8276
rect 25004 8236 25010 8248
rect 25866 8236 25872 8248
rect 25924 8236 25930 8288
rect 26142 8236 26148 8288
rect 26200 8276 26206 8288
rect 28718 8276 28724 8288
rect 26200 8248 28724 8276
rect 26200 8236 26206 8248
rect 28718 8236 28724 8248
rect 28776 8236 28782 8288
rect 30282 8236 30288 8288
rect 30340 8276 30346 8288
rect 31036 8276 31064 8316
rect 33689 8313 33701 8316
rect 33735 8313 33747 8347
rect 33689 8307 33747 8313
rect 33870 8304 33876 8356
rect 33928 8344 33934 8356
rect 34333 8347 34391 8353
rect 34333 8344 34345 8347
rect 33928 8316 34345 8344
rect 33928 8304 33934 8316
rect 34333 8313 34345 8316
rect 34379 8313 34391 8347
rect 34333 8307 34391 8313
rect 34514 8304 34520 8356
rect 34572 8344 34578 8356
rect 34882 8344 34888 8356
rect 34572 8316 34888 8344
rect 34572 8304 34578 8316
rect 34882 8304 34888 8316
rect 34940 8304 34946 8356
rect 35250 8304 35256 8356
rect 35308 8344 35314 8356
rect 35434 8344 35440 8356
rect 35308 8316 35440 8344
rect 35308 8304 35314 8316
rect 35434 8304 35440 8316
rect 35492 8304 35498 8356
rect 36262 8344 36268 8356
rect 36223 8316 36268 8344
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 38194 8344 38200 8356
rect 38155 8316 38200 8344
rect 38194 8304 38200 8316
rect 38252 8304 38258 8356
rect 30340 8248 31064 8276
rect 30340 8236 30346 8248
rect 31662 8236 31668 8288
rect 31720 8276 31726 8288
rect 34238 8276 34244 8288
rect 31720 8248 34244 8276
rect 31720 8236 31726 8248
rect 34238 8236 34244 8248
rect 34296 8236 34302 8288
rect 34422 8236 34428 8288
rect 34480 8276 34486 8288
rect 36998 8276 37004 8288
rect 34480 8248 37004 8276
rect 34480 8236 34486 8248
rect 36998 8236 37004 8248
rect 37056 8236 37062 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1578 8072 1584 8084
rect 1452 8044 1584 8072
rect 1452 8032 1458 8044
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 4706 8072 4712 8084
rect 4667 8044 4712 8072
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 5350 8072 5356 8084
rect 5311 8044 5356 8072
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 15746 8072 15752 8084
rect 6236 8044 15752 8072
rect 6236 8032 6242 8044
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 20806 8072 20812 8084
rect 17000 8044 20812 8072
rect 17000 8032 17006 8044
rect 20806 8032 20812 8044
rect 20864 8032 20870 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 24762 8072 24768 8084
rect 21048 8044 24768 8072
rect 21048 8032 21054 8044
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 27890 8072 27896 8084
rect 24912 8044 27896 8072
rect 24912 8032 24918 8044
rect 27890 8032 27896 8044
rect 27948 8032 27954 8084
rect 28721 8075 28779 8081
rect 28721 8041 28733 8075
rect 28767 8072 28779 8075
rect 31938 8072 31944 8084
rect 28767 8044 31944 8072
rect 28767 8041 28779 8044
rect 28721 8035 28779 8041
rect 31938 8032 31944 8044
rect 31996 8032 32002 8084
rect 32030 8032 32036 8084
rect 32088 8072 32094 8084
rect 33134 8072 33140 8084
rect 32088 8044 33140 8072
rect 32088 8032 32094 8044
rect 33134 8032 33140 8044
rect 33192 8032 33198 8084
rect 33962 8032 33968 8084
rect 34020 8072 34026 8084
rect 34422 8072 34428 8084
rect 34020 8044 34428 8072
rect 34020 8032 34026 8044
rect 34422 8032 34428 8044
rect 34480 8032 34486 8084
rect 34698 8032 34704 8084
rect 34756 8072 34762 8084
rect 34977 8075 35035 8081
rect 34977 8072 34989 8075
rect 34756 8044 34989 8072
rect 34756 8032 34762 8044
rect 34977 8041 34989 8044
rect 35023 8041 35035 8075
rect 35618 8072 35624 8084
rect 35579 8044 35624 8072
rect 34977 8035 35035 8041
rect 35618 8032 35624 8044
rect 35676 8032 35682 8084
rect 3786 8004 3792 8016
rect 1596 7976 3792 8004
rect 1596 7877 1624 7976
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 8018 8004 8024 8016
rect 4111 7976 8024 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11241 8007 11299 8013
rect 11241 8004 11253 8007
rect 11112 7976 11253 8004
rect 11112 7964 11118 7976
rect 11241 7973 11253 7976
rect 11287 7973 11299 8007
rect 11241 7967 11299 7973
rect 13078 7964 13084 8016
rect 13136 7964 13142 8016
rect 16206 7964 16212 8016
rect 16264 8004 16270 8016
rect 16264 7976 17264 8004
rect 16264 7964 16270 7976
rect 2608 7908 5304 7936
rect 2608 7877 2636 7908
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 3108 7840 3249 7868
rect 3108 7828 3114 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4890 7868 4896 7880
rect 4663 7840 4896 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 3988 7800 4016 7831
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5276 7877 5304 7908
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 7006 7936 7012 7948
rect 5500 7908 7012 7936
rect 5500 7896 5506 7908
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7432 7908 7573 7936
rect 7432 7896 7438 7908
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 9214 7936 9220 7948
rect 7892 7908 9220 7936
rect 7892 7896 7898 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 12342 7936 12348 7948
rect 9815 7908 12348 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 13096 7936 13124 7964
rect 12492 7908 13124 7936
rect 12492 7896 12498 7908
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13596 7908 13737 7936
rect 13596 7896 13602 7908
rect 13725 7905 13737 7908
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 15197 7939 15255 7945
rect 15197 7905 15209 7939
rect 15243 7936 15255 7939
rect 15286 7936 15292 7948
rect 15243 7908 15292 7936
rect 15243 7905 15255 7908
rect 15197 7899 15255 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 15620 7908 16804 7936
rect 15620 7896 15626 7908
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5350 7868 5356 7880
rect 5307 7840 5356 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9456 7840 9505 7868
rect 9456 7828 9462 7840
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11514 7868 11520 7880
rect 11388 7840 11520 7868
rect 11388 7828 11394 7840
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13964 7840 14289 7868
rect 13964 7828 13970 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14642 7828 14648 7880
rect 14700 7868 14706 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14700 7840 14933 7868
rect 14700 7828 14706 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 16298 7828 16304 7880
rect 16356 7828 16362 7880
rect 16776 7868 16804 7908
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16908 7908 17141 7936
rect 16908 7896 16914 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17236 7936 17264 7976
rect 18506 7964 18512 8016
rect 18564 8004 18570 8016
rect 24673 8007 24731 8013
rect 18564 7976 19564 8004
rect 18564 7964 18570 7976
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17236 7908 17417 7936
rect 17129 7899 17187 7905
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 19392 7908 19441 7936
rect 19392 7896 19398 7908
rect 19429 7905 19441 7908
rect 19475 7905 19487 7939
rect 19536 7936 19564 7976
rect 24673 7973 24685 8007
rect 24719 8004 24731 8007
rect 26142 8004 26148 8016
rect 24719 7976 26148 8004
rect 24719 7973 24731 7976
rect 24673 7967 24731 7973
rect 26142 7964 26148 7976
rect 26200 7964 26206 8016
rect 28074 7964 28080 8016
rect 28132 8004 28138 8016
rect 28902 8004 28908 8016
rect 28132 7976 28908 8004
rect 28132 7964 28138 7976
rect 28902 7964 28908 7976
rect 28960 7964 28966 8016
rect 30926 7964 30932 8016
rect 30984 8004 30990 8016
rect 32490 8004 32496 8016
rect 30984 7976 32496 8004
rect 30984 7964 30990 7976
rect 32490 7964 32496 7976
rect 32548 7964 32554 8016
rect 34238 7964 34244 8016
rect 34296 8004 34302 8016
rect 36909 8007 36967 8013
rect 36909 8004 36921 8007
rect 34296 7976 36921 8004
rect 34296 7964 34302 7976
rect 36909 7973 36921 7976
rect 36955 7973 36967 8007
rect 36909 7967 36967 7973
rect 20162 7936 20168 7948
rect 19536 7908 20168 7936
rect 19429 7899 19487 7905
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 21453 7939 21511 7945
rect 21453 7936 21465 7939
rect 21232 7908 21465 7936
rect 21232 7896 21238 7908
rect 21453 7905 21465 7908
rect 21499 7905 21511 7939
rect 22002 7936 22008 7948
rect 21963 7908 22008 7936
rect 21453 7899 21511 7905
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 22281 7939 22339 7945
rect 22281 7905 22293 7939
rect 22327 7936 22339 7939
rect 23014 7936 23020 7948
rect 22327 7908 23020 7936
rect 22327 7905 22339 7908
rect 22281 7899 22339 7905
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 23753 7939 23811 7945
rect 23753 7905 23765 7939
rect 23799 7936 23811 7939
rect 26237 7939 26295 7945
rect 23799 7908 26188 7936
rect 23799 7905 23811 7908
rect 23753 7899 23811 7905
rect 17034 7868 17040 7880
rect 16776 7840 17040 7868
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 24394 7828 24400 7880
rect 24452 7868 24458 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24452 7840 24593 7868
rect 24452 7828 24458 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 25958 7868 25964 7880
rect 25639 7840 25964 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 25958 7828 25964 7840
rect 26016 7828 26022 7880
rect 26160 7868 26188 7908
rect 26237 7905 26249 7939
rect 26283 7936 26295 7939
rect 26970 7936 26976 7948
rect 26283 7908 26976 7936
rect 26283 7905 26295 7908
rect 26237 7899 26295 7905
rect 26970 7896 26976 7908
rect 27028 7936 27034 7948
rect 27154 7936 27160 7948
rect 27028 7908 27160 7936
rect 27028 7896 27034 7908
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 31662 7936 31668 7948
rect 27816 7908 31668 7936
rect 26160 7840 26280 7868
rect 26252 7812 26280 7840
rect 27614 7828 27620 7880
rect 27672 7828 27678 7880
rect 5718 7800 5724 7812
rect 3988 7772 5724 7800
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 5810 7760 5816 7812
rect 5868 7800 5874 7812
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 5868 7772 6009 7800
rect 5868 7760 5874 7772
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 5997 7763 6055 7769
rect 6086 7760 6092 7812
rect 6144 7800 6150 7812
rect 6144 7772 6189 7800
rect 6144 7760 6150 7772
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6880 7772 7021 7800
rect 6880 7760 6886 7772
rect 7009 7769 7021 7772
rect 7055 7800 7067 7803
rect 7374 7800 7380 7812
rect 7055 7772 7380 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 7653 7803 7711 7809
rect 7653 7769 7665 7803
rect 7699 7800 7711 7803
rect 8570 7800 8576 7812
rect 7699 7772 7785 7800
rect 8531 7772 8576 7800
rect 7699 7769 7711 7772
rect 7653 7763 7711 7769
rect 1762 7732 1768 7744
rect 1723 7704 1768 7732
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2556 7704 2697 7732
rect 2556 7692 2562 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 3326 7732 3332 7744
rect 3287 7704 3332 7732
rect 2685 7695 2743 7701
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 7190 7732 7196 7744
rect 4120 7704 7196 7732
rect 4120 7692 4126 7704
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7757 7732 7785 7772
rect 8570 7760 8576 7772
rect 8628 7760 8634 7812
rect 10502 7760 10508 7812
rect 10560 7760 10566 7812
rect 11977 7803 12035 7809
rect 11977 7769 11989 7803
rect 12023 7800 12035 7803
rect 12066 7800 12072 7812
rect 12023 7772 12072 7800
rect 12023 7769 12035 7772
rect 11977 7763 12035 7769
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 12986 7760 12992 7812
rect 13044 7760 13050 7812
rect 15470 7800 15476 7812
rect 14292 7772 15476 7800
rect 7834 7732 7840 7744
rect 7757 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 11238 7732 11244 7744
rect 9180 7704 11244 7732
rect 9180 7692 9186 7704
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 14292 7732 14320 7772
rect 15470 7760 15476 7772
rect 15528 7760 15534 7812
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 16540 7772 17356 7800
rect 16540 7760 16546 7772
rect 11388 7704 14320 7732
rect 14369 7735 14427 7741
rect 11388 7692 11394 7704
rect 14369 7701 14381 7735
rect 14415 7732 14427 7735
rect 16574 7732 16580 7744
rect 14415 7704 16580 7732
rect 14415 7701 14427 7704
rect 14369 7695 14427 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 17126 7732 17132 7744
rect 16715 7704 17132 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17328 7732 17356 7772
rect 18966 7760 18972 7812
rect 19024 7800 19030 7812
rect 19426 7800 19432 7812
rect 19024 7772 19432 7800
rect 19024 7760 19030 7772
rect 19426 7760 19432 7772
rect 19484 7760 19490 7812
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7769 19763 7803
rect 22186 7800 22192 7812
rect 20930 7772 22192 7800
rect 19705 7763 19763 7769
rect 18322 7732 18328 7744
rect 17328 7704 18328 7732
rect 18322 7692 18328 7704
rect 18380 7732 18386 7744
rect 18877 7735 18935 7741
rect 18877 7732 18889 7735
rect 18380 7704 18889 7732
rect 18380 7692 18386 7704
rect 18877 7701 18889 7704
rect 18923 7701 18935 7735
rect 19720 7732 19748 7763
rect 22186 7760 22192 7772
rect 22244 7760 22250 7812
rect 26142 7800 26148 7812
rect 23506 7772 26148 7800
rect 26142 7760 26148 7772
rect 26200 7760 26206 7812
rect 26234 7760 26240 7812
rect 26292 7760 26298 7812
rect 26510 7800 26516 7812
rect 26471 7772 26516 7800
rect 26510 7760 26516 7772
rect 26568 7760 26574 7812
rect 21266 7732 21272 7744
rect 19720 7704 21272 7732
rect 18877 7695 18935 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 21818 7692 21824 7744
rect 21876 7732 21882 7744
rect 22554 7732 22560 7744
rect 21876 7704 22560 7732
rect 21876 7692 21882 7704
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 25685 7735 25743 7741
rect 25685 7701 25697 7735
rect 25731 7732 25743 7735
rect 27816 7732 27844 7908
rect 31662 7896 31668 7908
rect 31720 7896 31726 7948
rect 32401 7939 32459 7945
rect 32401 7905 32413 7939
rect 32447 7936 32459 7939
rect 35710 7936 35716 7948
rect 32447 7908 35716 7936
rect 32447 7905 32459 7908
rect 32401 7899 32459 7905
rect 35710 7896 35716 7908
rect 35768 7896 35774 7948
rect 36078 7896 36084 7948
rect 36136 7896 36142 7948
rect 27890 7828 27896 7880
rect 27948 7868 27954 7880
rect 27948 7840 28396 7868
rect 27948 7828 27954 7840
rect 28258 7800 28264 7812
rect 28219 7772 28264 7800
rect 28258 7760 28264 7772
rect 28316 7760 28322 7812
rect 28368 7800 28396 7840
rect 28534 7828 28540 7880
rect 28592 7868 28598 7880
rect 28905 7871 28963 7877
rect 28905 7868 28917 7871
rect 28592 7840 28917 7868
rect 28592 7828 28598 7840
rect 28905 7837 28917 7840
rect 28951 7837 28963 7871
rect 28905 7831 28963 7837
rect 29362 7828 29368 7880
rect 29420 7868 29426 7880
rect 30469 7871 30527 7877
rect 30469 7868 30481 7871
rect 29420 7840 30481 7868
rect 29420 7828 29426 7840
rect 30469 7837 30481 7840
rect 30515 7837 30527 7871
rect 30469 7831 30527 7837
rect 32861 7871 32919 7877
rect 32861 7837 32873 7871
rect 32907 7868 32919 7871
rect 33226 7868 33232 7880
rect 32907 7840 33232 7868
rect 32907 7837 32919 7840
rect 32861 7831 32919 7837
rect 33226 7828 33232 7840
rect 33284 7828 33290 7880
rect 33502 7868 33508 7880
rect 33463 7840 33508 7868
rect 33502 7828 33508 7840
rect 33560 7828 33566 7880
rect 34149 7871 34207 7877
rect 34149 7837 34161 7871
rect 34195 7868 34207 7871
rect 34238 7868 34244 7880
rect 34195 7840 34244 7868
rect 34195 7837 34207 7840
rect 34149 7831 34207 7837
rect 34238 7828 34244 7840
rect 34296 7828 34302 7880
rect 34885 7871 34943 7877
rect 34885 7837 34897 7871
rect 34931 7837 34943 7871
rect 34885 7831 34943 7837
rect 35529 7871 35587 7877
rect 35529 7837 35541 7871
rect 35575 7868 35587 7871
rect 36096 7868 36124 7896
rect 36173 7871 36231 7877
rect 36173 7868 36185 7871
rect 35575 7840 36185 7868
rect 35575 7837 35587 7840
rect 35529 7831 35587 7837
rect 36173 7837 36185 7840
rect 36219 7837 36231 7871
rect 36814 7868 36820 7880
rect 36775 7840 36820 7868
rect 36173 7831 36231 7837
rect 29733 7803 29791 7809
rect 29733 7800 29745 7803
rect 28368 7772 29745 7800
rect 29733 7769 29745 7772
rect 29779 7769 29791 7803
rect 31389 7803 31447 7809
rect 31389 7800 31401 7803
rect 29733 7763 29791 7769
rect 31312 7772 31401 7800
rect 25731 7704 27844 7732
rect 25731 7701 25743 7704
rect 25685 7695 25743 7701
rect 27890 7692 27896 7744
rect 27948 7732 27954 7744
rect 30006 7732 30012 7744
rect 27948 7704 30012 7732
rect 27948 7692 27954 7704
rect 30006 7692 30012 7704
rect 30064 7692 30070 7744
rect 31312 7732 31340 7772
rect 31389 7769 31401 7772
rect 31435 7769 31447 7803
rect 31389 7763 31447 7769
rect 31481 7803 31539 7809
rect 31481 7769 31493 7803
rect 31527 7800 31539 7803
rect 33594 7800 33600 7812
rect 31527 7772 33456 7800
rect 33555 7772 33600 7800
rect 31527 7769 31539 7772
rect 31481 7763 31539 7769
rect 31570 7732 31576 7744
rect 31312 7704 31576 7732
rect 31570 7692 31576 7704
rect 31628 7692 31634 7744
rect 31662 7692 31668 7744
rect 31720 7732 31726 7744
rect 32953 7735 33011 7741
rect 32953 7732 32965 7735
rect 31720 7704 32965 7732
rect 31720 7692 31726 7704
rect 32953 7701 32965 7704
rect 32999 7701 33011 7735
rect 33428 7732 33456 7772
rect 33594 7760 33600 7772
rect 33652 7760 33658 7812
rect 34900 7800 34928 7831
rect 36814 7828 36820 7840
rect 36872 7828 36878 7880
rect 37918 7828 37924 7880
rect 37976 7868 37982 7880
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 37976 7840 38025 7868
rect 37976 7828 37982 7840
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 38102 7800 38108 7812
rect 33980 7772 34836 7800
rect 34900 7772 38108 7800
rect 33980 7732 34008 7772
rect 33428 7704 34008 7732
rect 32953 7695 33011 7701
rect 34054 7692 34060 7744
rect 34112 7732 34118 7744
rect 34241 7735 34299 7741
rect 34241 7732 34253 7735
rect 34112 7704 34253 7732
rect 34112 7692 34118 7704
rect 34241 7701 34253 7704
rect 34287 7701 34299 7735
rect 34808 7732 34836 7772
rect 38102 7760 38108 7772
rect 38160 7760 38166 7812
rect 35250 7732 35256 7744
rect 34808 7704 35256 7732
rect 34241 7695 34299 7701
rect 35250 7692 35256 7704
rect 35308 7692 35314 7744
rect 35710 7692 35716 7744
rect 35768 7732 35774 7744
rect 36265 7735 36323 7741
rect 36265 7732 36277 7735
rect 35768 7704 36277 7732
rect 35768 7692 35774 7704
rect 36265 7701 36277 7704
rect 36311 7701 36323 7735
rect 38194 7732 38200 7744
rect 38155 7704 38200 7732
rect 36265 7695 36323 7701
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 3970 7528 3976 7540
rect 3931 7500 3976 7528
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 6086 7528 6092 7540
rect 4663 7500 6092 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 11330 7528 11336 7540
rect 8956 7500 11336 7528
rect 2130 7460 2136 7472
rect 2091 7432 2136 7460
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 4856 7432 6837 7460
rect 4856 7420 4862 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 7558 7420 7564 7472
rect 7616 7460 7622 7472
rect 7929 7463 7987 7469
rect 7929 7460 7941 7463
rect 7616 7432 7941 7460
rect 7616 7420 7622 7432
rect 7929 7429 7941 7432
rect 7975 7429 7987 7463
rect 7929 7423 7987 7429
rect 8021 7463 8079 7469
rect 8021 7429 8033 7463
rect 8067 7460 8079 7463
rect 8386 7460 8392 7472
rect 8067 7432 8392 7460
rect 8067 7429 8079 7432
rect 8021 7423 8079 7429
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 8956 7469 8984 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 11839 7500 15700 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 8941 7463 8999 7469
rect 8941 7429 8953 7463
rect 8987 7429 8999 7463
rect 9950 7460 9956 7472
rect 8941 7423 8999 7429
rect 9048 7432 9956 7460
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2958 7392 2964 7404
rect 2823 7364 2964 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2056 7324 2084 7355
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3786 7392 3792 7404
rect 3283 7364 3792 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 3936 7364 3981 7392
rect 3936 7352 3942 7364
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4522 7392 4528 7404
rect 4212 7364 4528 7392
rect 4212 7352 4218 7364
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 5132 7364 5181 7392
rect 5132 7352 5138 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5684 7364 5825 7392
rect 5684 7352 5690 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 4614 7324 4620 7336
rect 2056 7296 4620 7324
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 6362 7324 6368 7336
rect 5307 7296 6368 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6730 7324 6736 7336
rect 6691 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7064 7296 7109 7324
rect 7064 7284 7070 7296
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 9048 7324 9076 7432
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 10410 7420 10416 7472
rect 10468 7420 10474 7472
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 11296 7432 12633 7460
rect 11296 7420 11302 7432
rect 12621 7429 12633 7432
rect 12667 7429 12679 7463
rect 12621 7423 12679 7429
rect 14369 7463 14427 7469
rect 14369 7429 14381 7463
rect 14415 7460 14427 7463
rect 14458 7460 14464 7472
rect 14415 7432 14464 7460
rect 14415 7429 14427 7432
rect 14369 7423 14427 7429
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 14642 7420 14648 7472
rect 14700 7460 14706 7472
rect 15565 7463 15623 7469
rect 15565 7460 15577 7463
rect 14700 7432 15577 7460
rect 14700 7420 14706 7432
rect 15565 7429 15577 7432
rect 15611 7429 15623 7463
rect 15672 7460 15700 7500
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 16942 7528 16948 7540
rect 15804 7500 16948 7528
rect 15804 7488 15810 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 17828 7500 19840 7528
rect 17828 7488 17834 7500
rect 18322 7460 18328 7472
rect 15672 7432 18328 7460
rect 15565 7423 15623 7429
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 18690 7420 18696 7472
rect 18748 7420 18754 7472
rect 19812 7469 19840 7500
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20864 7500 20913 7528
rect 20864 7488 20870 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 20901 7491 20959 7497
rect 23566 7488 23572 7540
rect 23624 7528 23630 7540
rect 23753 7531 23811 7537
rect 23753 7528 23765 7531
rect 23624 7500 23765 7528
rect 23624 7488 23630 7500
rect 23753 7497 23765 7500
rect 23799 7497 23811 7531
rect 23753 7491 23811 7497
rect 25961 7531 26019 7537
rect 25961 7497 25973 7531
rect 26007 7528 26019 7531
rect 27154 7528 27160 7540
rect 26007 7500 27160 7528
rect 26007 7497 26019 7500
rect 25961 7491 26019 7497
rect 27154 7488 27160 7500
rect 27212 7488 27218 7540
rect 27338 7488 27344 7540
rect 27396 7528 27402 7540
rect 28074 7528 28080 7540
rect 27396 7500 28080 7528
rect 27396 7488 27402 7500
rect 28074 7488 28080 7500
rect 28132 7488 28138 7540
rect 28258 7488 28264 7540
rect 28316 7528 28322 7540
rect 30466 7528 30472 7540
rect 28316 7500 30472 7528
rect 28316 7488 28322 7500
rect 19797 7463 19855 7469
rect 19797 7429 19809 7463
rect 19843 7429 19855 7463
rect 20714 7460 20720 7472
rect 19797 7423 19855 7429
rect 20272 7432 20720 7460
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 11790 7392 11796 7404
rect 11747 7364 11796 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 9398 7324 9404 7336
rect 7616 7296 9076 7324
rect 9359 7296 9404 7324
rect 7616 7284 7622 7296
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7324 9735 7327
rect 11054 7324 11060 7336
rect 9723 7296 11060 7324
rect 9723 7293 9735 7296
rect 9677 7287 9735 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 12342 7324 12348 7336
rect 12303 7296 12348 7324
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 13740 7324 13768 7378
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14332 7364 14841 7392
rect 14332 7352 14338 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 16022 7352 16028 7404
rect 16080 7392 16086 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16080 7364 16957 7392
rect 16080 7352 16086 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20272 7401 20300 7432
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 22278 7460 22284 7472
rect 22239 7432 22284 7460
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 22554 7420 22560 7472
rect 22612 7460 22618 7472
rect 22612 7432 22770 7460
rect 22612 7420 22618 7432
rect 25222 7420 25228 7472
rect 25280 7420 25286 7472
rect 27430 7420 27436 7472
rect 27488 7460 27494 7472
rect 28902 7460 28908 7472
rect 27488 7432 27533 7460
rect 28658 7432 28908 7460
rect 27488 7420 27494 7432
rect 28902 7420 28908 7432
rect 28960 7420 28966 7472
rect 29656 7469 29684 7500
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 31570 7488 31576 7540
rect 31628 7528 31634 7540
rect 31665 7531 31723 7537
rect 31665 7528 31677 7531
rect 31628 7500 31677 7528
rect 31628 7488 31634 7500
rect 31665 7497 31677 7500
rect 31711 7497 31723 7531
rect 31665 7491 31723 7497
rect 32416 7500 32812 7528
rect 29641 7463 29699 7469
rect 29641 7429 29653 7463
rect 29687 7429 29699 7463
rect 32030 7460 32036 7472
rect 30866 7432 32036 7460
rect 29641 7423 29699 7429
rect 32030 7420 32036 7432
rect 32088 7420 32094 7472
rect 32416 7469 32444 7500
rect 32401 7463 32459 7469
rect 32401 7429 32413 7463
rect 32447 7429 32459 7463
rect 32401 7423 32459 7429
rect 32493 7463 32551 7469
rect 32493 7429 32505 7463
rect 32539 7460 32551 7463
rect 32582 7460 32588 7472
rect 32539 7432 32588 7460
rect 32539 7429 32551 7432
rect 32493 7423 32551 7429
rect 32582 7420 32588 7432
rect 32640 7420 32646 7472
rect 32784 7460 32812 7500
rect 34054 7488 34060 7540
rect 34112 7528 34118 7540
rect 34149 7531 34207 7537
rect 34149 7528 34161 7531
rect 34112 7500 34161 7528
rect 34112 7488 34118 7500
rect 34149 7497 34161 7500
rect 34195 7497 34207 7531
rect 34149 7491 34207 7497
rect 35618 7488 35624 7540
rect 35676 7528 35682 7540
rect 36814 7528 36820 7540
rect 35676 7500 36820 7528
rect 35676 7488 35682 7500
rect 36814 7488 36820 7500
rect 36872 7488 36878 7540
rect 36998 7488 37004 7540
rect 37056 7528 37062 7540
rect 37553 7531 37611 7537
rect 37553 7528 37565 7531
rect 37056 7500 37565 7528
rect 37056 7488 37062 7500
rect 37553 7497 37565 7500
rect 37599 7497 37611 7531
rect 37553 7491 37611 7497
rect 34698 7460 34704 7472
rect 32784 7432 34704 7460
rect 34698 7420 34704 7432
rect 34756 7420 34762 7472
rect 35250 7420 35256 7472
rect 35308 7460 35314 7472
rect 36173 7463 36231 7469
rect 36173 7460 36185 7463
rect 35308 7432 36185 7460
rect 35308 7420 35314 7432
rect 36173 7429 36185 7432
rect 36219 7429 36231 7463
rect 36173 7423 36231 7429
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20220 7364 20269 7392
rect 20220 7352 20226 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 20404 7364 21097 7392
rect 20404 7352 20410 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 21085 7355 21143 7361
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 26234 7352 26240 7404
rect 26292 7392 26298 7404
rect 26605 7395 26663 7401
rect 26605 7392 26617 7395
rect 26292 7364 26617 7392
rect 26292 7352 26298 7364
rect 26605 7361 26617 7364
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 26970 7352 26976 7404
rect 27028 7396 27034 7404
rect 27146 7396 27204 7401
rect 27028 7395 27204 7396
rect 27028 7368 27158 7395
rect 27028 7352 27034 7368
rect 27146 7361 27158 7368
rect 27192 7361 27204 7395
rect 29086 7392 29092 7404
rect 27146 7355 27204 7361
rect 28644 7364 29092 7392
rect 16758 7324 16764 7336
rect 13740 7296 16764 7324
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 16908 7296 17785 7324
rect 16908 7284 16914 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7324 18107 7327
rect 18506 7324 18512 7336
rect 18095 7296 18512 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18506 7284 18512 7296
rect 18564 7324 18570 7336
rect 20990 7324 20996 7336
rect 18564 7296 20996 7324
rect 18564 7284 18570 7296
rect 20990 7284 20996 7296
rect 21048 7284 21054 7336
rect 21542 7284 21548 7336
rect 21600 7324 21606 7336
rect 24026 7324 24032 7336
rect 21600 7296 24032 7324
rect 21600 7284 21606 7296
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 24210 7324 24216 7336
rect 24171 7296 24216 7324
rect 24210 7284 24216 7296
rect 24268 7284 24274 7336
rect 24489 7327 24547 7333
rect 24489 7293 24501 7327
rect 24535 7324 24547 7327
rect 26694 7324 26700 7336
rect 24535 7296 26700 7324
rect 24535 7293 24547 7296
rect 24489 7287 24547 7293
rect 26694 7284 26700 7296
rect 26752 7284 26758 7336
rect 27522 7284 27528 7336
rect 27580 7324 27586 7336
rect 28644 7324 28672 7364
rect 29086 7352 29092 7364
rect 29144 7352 29150 7404
rect 29362 7392 29368 7404
rect 29323 7364 29368 7392
rect 29362 7352 29368 7364
rect 29420 7352 29426 7404
rect 31573 7395 31631 7401
rect 31573 7361 31585 7395
rect 31619 7392 31631 7395
rect 31846 7392 31852 7404
rect 31619 7364 31852 7392
rect 31619 7361 31631 7364
rect 31573 7355 31631 7361
rect 31846 7352 31852 7364
rect 31904 7352 31910 7404
rect 33045 7395 33103 7401
rect 33045 7361 33057 7395
rect 33091 7392 33103 7395
rect 33134 7392 33140 7404
rect 33091 7364 33140 7392
rect 33091 7361 33103 7364
rect 33045 7355 33103 7361
rect 33134 7352 33140 7364
rect 33192 7352 33198 7404
rect 33502 7392 33508 7404
rect 33463 7364 33508 7392
rect 33502 7352 33508 7364
rect 33560 7352 33566 7404
rect 34793 7395 34851 7401
rect 33612 7390 34744 7392
rect 34793 7390 34805 7395
rect 33612 7364 34805 7390
rect 27580 7296 28672 7324
rect 27580 7284 27586 7296
rect 28902 7284 28908 7336
rect 28960 7324 28966 7336
rect 33612 7324 33640 7364
rect 34716 7362 34805 7364
rect 34793 7361 34805 7362
rect 34839 7361 34851 7395
rect 34793 7355 34851 7361
rect 36081 7395 36139 7401
rect 36081 7361 36093 7395
rect 36127 7361 36139 7395
rect 36081 7355 36139 7361
rect 36909 7395 36967 7401
rect 36909 7361 36921 7395
rect 36955 7392 36967 7395
rect 36998 7392 37004 7404
rect 36955 7364 37004 7392
rect 36955 7361 36967 7364
rect 36909 7355 36967 7361
rect 28960 7296 30696 7324
rect 28960 7284 28966 7296
rect 4632 7256 4660 7284
rect 5442 7256 5448 7268
rect 4632 7228 5448 7256
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 9030 7256 9036 7268
rect 5951 7228 9036 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 11149 7259 11207 7265
rect 11149 7225 11161 7259
rect 11195 7256 11207 7259
rect 12250 7256 12256 7268
rect 11195 7228 12256 7256
rect 11195 7225 11207 7228
rect 11149 7219 11207 7225
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 16390 7256 16396 7268
rect 13780 7228 16396 7256
rect 13780 7216 13786 7228
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 17037 7259 17095 7265
rect 17037 7225 17049 7259
rect 17083 7256 17095 7259
rect 17083 7228 17908 7256
rect 17083 7225 17095 7228
rect 17037 7219 17095 7225
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 2682 7188 2688 7200
rect 2639 7160 2688 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3510 7188 3516 7200
rect 3375 7160 3516 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 11790 7188 11796 7200
rect 6604 7160 11796 7188
rect 6604 7148 6610 7160
rect 11790 7148 11796 7160
rect 11848 7188 11854 7200
rect 14734 7188 14740 7200
rect 11848 7160 14740 7188
rect 11848 7148 11854 7160
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16942 7188 16948 7200
rect 16264 7160 16948 7188
rect 16264 7148 16270 7160
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 17494 7188 17500 7200
rect 17184 7160 17500 7188
rect 17184 7148 17190 7160
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 17880 7188 17908 7228
rect 19426 7216 19432 7268
rect 19484 7256 19490 7268
rect 20622 7256 20628 7268
rect 19484 7228 20628 7256
rect 19484 7216 19490 7228
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 26421 7259 26479 7265
rect 26421 7225 26433 7259
rect 26467 7256 26479 7259
rect 26602 7256 26608 7268
rect 26467 7228 26608 7256
rect 26467 7225 26479 7228
rect 26421 7219 26479 7225
rect 26602 7216 26608 7228
rect 26660 7216 26666 7268
rect 30668 7256 30696 7296
rect 32232 7296 33640 7324
rect 32232 7256 32260 7296
rect 33686 7284 33692 7336
rect 33744 7324 33750 7336
rect 35437 7327 35495 7333
rect 35437 7324 35449 7327
rect 33744 7296 35449 7324
rect 33744 7284 33750 7296
rect 35437 7293 35449 7296
rect 35483 7293 35495 7327
rect 35437 7287 35495 7293
rect 35710 7284 35716 7336
rect 35768 7324 35774 7336
rect 36096 7324 36124 7355
rect 36998 7352 37004 7364
rect 37056 7352 37062 7404
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7392 37519 7395
rect 37918 7392 37924 7404
rect 37507 7364 37924 7392
rect 37507 7361 37519 7364
rect 37461 7355 37519 7361
rect 37918 7352 37924 7364
rect 37976 7352 37982 7404
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 35768 7296 36124 7324
rect 35768 7284 35774 7296
rect 30668 7228 32260 7256
rect 32858 7216 32864 7268
rect 32916 7256 32922 7268
rect 34885 7259 34943 7265
rect 34885 7256 34897 7259
rect 32916 7228 34897 7256
rect 32916 7216 32922 7228
rect 34885 7225 34897 7228
rect 34931 7225 34943 7259
rect 34885 7219 34943 7225
rect 20162 7188 20168 7200
rect 17880 7160 20168 7188
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 20349 7191 20407 7197
rect 20349 7157 20361 7191
rect 20395 7188 20407 7191
rect 20806 7188 20812 7200
rect 20395 7160 20812 7188
rect 20395 7157 20407 7160
rect 20349 7151 20407 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 28534 7188 28540 7200
rect 25924 7160 28540 7188
rect 25924 7148 25930 7160
rect 28534 7148 28540 7160
rect 28592 7148 28598 7200
rect 28810 7148 28816 7200
rect 28868 7188 28874 7200
rect 28905 7191 28963 7197
rect 28905 7188 28917 7191
rect 28868 7160 28917 7188
rect 28868 7148 28874 7160
rect 28905 7157 28917 7160
rect 28951 7157 28963 7191
rect 28905 7151 28963 7157
rect 31113 7191 31171 7197
rect 31113 7157 31125 7191
rect 31159 7188 31171 7191
rect 31294 7188 31300 7200
rect 31159 7160 31300 7188
rect 31159 7157 31171 7160
rect 31113 7151 31171 7157
rect 31294 7148 31300 7160
rect 31352 7148 31358 7200
rect 32030 7148 32036 7200
rect 32088 7188 32094 7200
rect 32214 7188 32220 7200
rect 32088 7160 32220 7188
rect 32088 7148 32094 7160
rect 32214 7148 32220 7160
rect 32272 7148 32278 7200
rect 33318 7148 33324 7200
rect 33376 7188 33382 7200
rect 33597 7191 33655 7197
rect 33597 7188 33609 7191
rect 33376 7160 33609 7188
rect 33376 7148 33382 7160
rect 33597 7157 33609 7160
rect 33643 7157 33655 7191
rect 33597 7151 33655 7157
rect 34146 7148 34152 7200
rect 34204 7188 34210 7200
rect 35618 7188 35624 7200
rect 34204 7160 35624 7188
rect 34204 7148 34210 7160
rect 35618 7148 35624 7160
rect 35676 7148 35682 7200
rect 36630 7148 36636 7200
rect 36688 7188 36694 7200
rect 36725 7191 36783 7197
rect 36725 7188 36737 7191
rect 36688 7160 36737 7188
rect 36688 7148 36694 7160
rect 36725 7157 36737 7160
rect 36771 7157 36783 7191
rect 38102 7188 38108 7200
rect 38063 7160 38108 7188
rect 36725 7151 36783 7157
rect 38102 7148 38108 7160
rect 38160 7148 38166 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 4154 6984 4160 6996
rect 3660 6956 4160 6984
rect 3660 6944 3666 6956
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6984 4399 6987
rect 5074 6984 5080 6996
rect 4387 6956 5080 6984
rect 4387 6953 4399 6956
rect 4341 6947 4399 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 7088 6987 7146 6993
rect 7088 6953 7100 6987
rect 7134 6984 7146 6987
rect 11882 6984 11888 6996
rect 7134 6956 11888 6984
rect 7134 6953 7146 6956
rect 7088 6947 7146 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12124 6956 12388 6984
rect 12124 6944 12130 6956
rect 2958 6876 2964 6928
rect 3016 6916 3022 6928
rect 12360 6916 12388 6956
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13722 6984 13728 6996
rect 12492 6956 13728 6984
rect 12492 6944 12498 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 16466 6987 16524 6993
rect 16466 6984 16478 6987
rect 14516 6956 16478 6984
rect 14516 6944 14522 6956
rect 16466 6953 16478 6956
rect 16512 6953 16524 6987
rect 16466 6947 16524 6953
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 20346 6984 20352 6996
rect 17000 6956 20352 6984
rect 17000 6944 17006 6956
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 20980 6987 21038 6993
rect 20980 6953 20992 6987
rect 21026 6984 21038 6987
rect 21542 6984 21548 6996
rect 21026 6956 21548 6984
rect 21026 6953 21038 6956
rect 20980 6947 21038 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 21634 6944 21640 6996
rect 21692 6984 21698 6996
rect 21692 6956 22094 6984
rect 21692 6944 21698 6956
rect 15378 6916 15384 6928
rect 3016 6888 6960 6916
rect 12360 6888 15384 6916
rect 3016 6876 3022 6888
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 4798 6848 4804 6860
rect 2731 6820 4804 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 6932 6848 6960 6888
rect 15378 6876 15384 6888
rect 15436 6916 15442 6928
rect 16114 6916 16120 6928
rect 15436 6888 16120 6916
rect 15436 6876 15442 6888
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 17494 6876 17500 6928
rect 17552 6916 17558 6928
rect 20622 6916 20628 6928
rect 17552 6888 20628 6916
rect 17552 6876 17558 6888
rect 20622 6876 20628 6888
rect 20680 6876 20686 6928
rect 22066 6916 22094 6956
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22830 6984 22836 6996
rect 22336 6956 22836 6984
rect 22336 6944 22342 6956
rect 22830 6944 22836 6956
rect 22888 6944 22894 6996
rect 24026 6944 24032 6996
rect 24084 6984 24090 6996
rect 26326 6984 26332 6996
rect 24084 6956 26332 6984
rect 24084 6944 24090 6956
rect 26326 6944 26332 6956
rect 26384 6944 26390 6996
rect 26500 6987 26558 6993
rect 26500 6953 26512 6987
rect 26546 6984 26558 6987
rect 28258 6984 28264 6996
rect 26546 6956 28264 6984
rect 26546 6953 26558 6956
rect 26500 6947 26558 6953
rect 28258 6944 28264 6956
rect 28316 6944 28322 6996
rect 28721 6987 28779 6993
rect 28721 6953 28733 6987
rect 28767 6984 28779 6987
rect 29822 6984 29828 6996
rect 28767 6956 29828 6984
rect 28767 6953 28779 6956
rect 28721 6947 28779 6953
rect 29822 6944 29828 6956
rect 29880 6944 29886 6996
rect 30006 6993 30012 6996
rect 29996 6987 30012 6993
rect 29996 6953 30008 6987
rect 29996 6947 30012 6953
rect 30006 6944 30012 6947
rect 30064 6944 30070 6996
rect 33686 6984 33692 6996
rect 32232 6956 33692 6984
rect 22066 6888 23428 6916
rect 7558 6848 7564 6860
rect 6932 6820 7564 6848
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9306 6848 9312 6860
rect 9263 6820 9312 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 9456 6820 11069 6848
rect 9456 6808 9462 6820
rect 11057 6817 11069 6820
rect 11103 6848 11115 6851
rect 11698 6848 11704 6860
rect 11103 6820 11704 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 11698 6808 11704 6820
rect 11756 6848 11762 6860
rect 12342 6848 12348 6860
rect 11756 6820 12348 6848
rect 11756 6808 11762 6820
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 12400 6820 15025 6848
rect 12400 6808 12406 6820
rect 15013 6817 15025 6820
rect 15059 6817 15071 6851
rect 15013 6811 15071 6817
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6848 16267 6851
rect 16850 6848 16856 6860
rect 16255 6820 16856 6848
rect 16255 6817 16267 6820
rect 16209 6811 16267 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 23293 6851 23351 6857
rect 23293 6848 23305 6851
rect 17092 6820 23305 6848
rect 17092 6808 17098 6820
rect 23293 6817 23305 6820
rect 23339 6817 23351 6851
rect 23400 6848 23428 6888
rect 27586 6888 29408 6916
rect 26142 6848 26148 6860
rect 23400 6820 26148 6848
rect 23293 6811 23351 6817
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2130 6780 2136 6792
rect 1995 6752 2136 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2590 6780 2596 6792
rect 2551 6752 2596 6780
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3970 6780 3976 6792
rect 3283 6752 3976 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4246 6780 4252 6792
rect 4207 6752 4252 6780
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 5074 6780 5080 6792
rect 5035 6752 5080 6780
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 6178 6780 6184 6792
rect 5583 6752 6184 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6822 6780 6828 6792
rect 6783 6752 6828 6780
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 3329 6715 3387 6721
rect 3329 6681 3341 6715
rect 3375 6712 3387 6715
rect 3375 6684 7512 6712
rect 3375 6681 3387 6684
rect 3329 6675 3387 6681
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5350 6644 5356 6656
rect 4939 6616 5356 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5592 6616 5641 6644
rect 5592 6604 5598 6616
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 5629 6607 5687 6613
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7484 6644 7512 6684
rect 7834 6672 7840 6724
rect 7892 6672 7898 6724
rect 9324 6712 9352 6808
rect 10962 6780 10968 6792
rect 10428 6752 10968 6780
rect 9585 6715 9643 6721
rect 9585 6712 9597 6715
rect 9324 6684 9597 6712
rect 9585 6681 9597 6684
rect 9631 6681 9643 6715
rect 9585 6675 9643 6681
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 9732 6684 9777 6712
rect 9732 6672 9738 6684
rect 9858 6672 9864 6724
rect 9916 6712 9922 6724
rect 10428 6712 10456 6752
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 13078 6780 13084 6792
rect 13039 6752 13084 6780
rect 13078 6740 13084 6752
rect 13136 6780 13142 6792
rect 13354 6780 13360 6792
rect 13136 6752 13360 6780
rect 13136 6740 13142 6752
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 18782 6780 18788 6792
rect 13679 6752 16252 6780
rect 17618 6752 18788 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 10594 6712 10600 6724
rect 9916 6684 10456 6712
rect 10555 6684 10600 6712
rect 9916 6672 9922 6684
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 11333 6715 11391 6721
rect 11333 6712 11345 6715
rect 10744 6684 11345 6712
rect 10744 6672 10750 6684
rect 11333 6681 11345 6684
rect 11379 6681 11391 6715
rect 11333 6675 11391 6681
rect 11974 6672 11980 6724
rect 12032 6672 12038 6724
rect 14274 6712 14280 6724
rect 14235 6684 14280 6712
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 15102 6712 15108 6724
rect 14568 6684 15108 6712
rect 8386 6644 8392 6656
rect 7484 6616 8392 6644
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 8573 6647 8631 6653
rect 8573 6644 8585 6647
rect 8536 6616 8585 6644
rect 8536 6604 8542 6616
rect 8573 6613 8585 6616
rect 8619 6644 8631 6647
rect 11606 6644 11612 6656
rect 8619 6616 11612 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 14090 6644 14096 6656
rect 12124 6616 14096 6644
rect 12124 6604 12130 6616
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14182 6604 14188 6656
rect 14240 6644 14246 6656
rect 14568 6644 14596 6684
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 16224 6712 16252 6752
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 18877 6783 18935 6789
rect 18877 6749 18889 6783
rect 18923 6749 18935 6783
rect 18877 6743 18935 6749
rect 16758 6712 16764 6724
rect 16224 6684 16764 6712
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 18233 6715 18291 6721
rect 18233 6712 18245 6715
rect 18012 6684 18245 6712
rect 18012 6672 18018 6684
rect 18233 6681 18245 6684
rect 18279 6681 18291 6715
rect 18892 6712 18920 6743
rect 19150 6740 19156 6792
rect 19208 6782 19214 6792
rect 19429 6783 19487 6789
rect 19208 6780 19334 6782
rect 19429 6780 19441 6783
rect 19208 6754 19441 6780
rect 19208 6740 19214 6754
rect 19306 6752 19441 6754
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 20714 6780 20720 6792
rect 20675 6752 20720 6780
rect 19429 6743 19487 6749
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 22738 6780 22744 6792
rect 22699 6752 22744 6780
rect 22738 6740 22744 6752
rect 22796 6740 22802 6792
rect 22830 6740 22836 6792
rect 22888 6780 22894 6792
rect 24596 6789 24624 6820
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26970 6848 26976 6860
rect 26283 6820 26976 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26970 6808 26976 6820
rect 27028 6848 27034 6860
rect 27154 6848 27160 6860
rect 27028 6820 27160 6848
rect 27028 6808 27034 6820
rect 27154 6808 27160 6820
rect 27212 6848 27218 6860
rect 27586 6848 27614 6888
rect 29380 6860 29408 6888
rect 27212 6820 27614 6848
rect 27212 6808 27218 6820
rect 27706 6808 27712 6860
rect 27764 6848 27770 6860
rect 28261 6851 28319 6857
rect 28261 6848 28273 6851
rect 27764 6820 28273 6848
rect 27764 6808 27770 6820
rect 28261 6817 28273 6820
rect 28307 6817 28319 6851
rect 28261 6811 28319 6817
rect 29362 6808 29368 6860
rect 29420 6848 29426 6860
rect 29733 6851 29791 6857
rect 29733 6848 29745 6851
rect 29420 6820 29745 6848
rect 29420 6808 29426 6820
rect 29733 6817 29745 6820
rect 29779 6817 29791 6851
rect 29733 6811 29791 6817
rect 32033 6851 32091 6857
rect 32033 6817 32045 6851
rect 32079 6848 32091 6851
rect 32232 6848 32260 6956
rect 33686 6944 33692 6956
rect 33744 6944 33750 6996
rect 34054 6944 34060 6996
rect 34112 6984 34118 6996
rect 36262 6984 36268 6996
rect 34112 6956 36268 6984
rect 34112 6944 34118 6956
rect 36262 6944 36268 6956
rect 36320 6944 36326 6996
rect 34422 6916 34428 6928
rect 32416 6888 34428 6916
rect 32416 6860 32444 6888
rect 34422 6876 34428 6888
rect 34480 6876 34486 6928
rect 36078 6916 36084 6928
rect 34532 6888 36084 6916
rect 32398 6848 32404 6860
rect 32079 6820 32260 6848
rect 32359 6820 32404 6848
rect 32079 6817 32091 6820
rect 32033 6811 32091 6817
rect 32398 6808 32404 6820
rect 32456 6808 32462 6860
rect 34532 6848 34560 6888
rect 36078 6876 36084 6888
rect 36136 6876 36142 6928
rect 34164 6820 34560 6848
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 22888 6752 23213 6780
rect 22888 6740 22894 6752
rect 23201 6749 23213 6752
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 25222 6780 25228 6792
rect 25183 6752 25228 6780
rect 24581 6743 24639 6749
rect 20438 6712 20444 6724
rect 18892 6684 20444 6712
rect 18233 6675 18291 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 23658 6712 23664 6724
rect 22218 6684 23664 6712
rect 23658 6672 23664 6684
rect 23716 6672 23722 6724
rect 23860 6712 23888 6743
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 27798 6740 27804 6792
rect 27856 6780 27862 6792
rect 28905 6783 28963 6789
rect 28905 6780 28917 6783
rect 27856 6752 28917 6780
rect 27856 6740 27862 6752
rect 28905 6749 28917 6752
rect 28951 6749 28963 6783
rect 31662 6780 31668 6792
rect 31142 6752 31668 6780
rect 28905 6743 28963 6749
rect 31662 6740 31668 6752
rect 31720 6740 31726 6792
rect 32950 6740 32956 6792
rect 33008 6780 33014 6792
rect 33505 6783 33563 6789
rect 33505 6780 33517 6783
rect 33008 6752 33517 6780
rect 33008 6740 33014 6752
rect 33505 6749 33517 6752
rect 33551 6749 33563 6783
rect 33505 6743 33563 6749
rect 33597 6783 33655 6789
rect 33597 6749 33609 6783
rect 33643 6780 33655 6783
rect 33778 6780 33784 6792
rect 33643 6752 33784 6780
rect 33643 6749 33655 6752
rect 33597 6743 33655 6749
rect 33778 6740 33784 6752
rect 33836 6740 33842 6792
rect 34164 6789 34192 6820
rect 34698 6808 34704 6860
rect 34756 6848 34762 6860
rect 34885 6851 34943 6857
rect 34885 6848 34897 6851
rect 34756 6820 34897 6848
rect 34756 6808 34762 6820
rect 34885 6817 34897 6820
rect 34931 6817 34943 6851
rect 35710 6848 35716 6860
rect 34885 6811 34943 6817
rect 34992 6820 35716 6848
rect 34149 6783 34207 6789
rect 34149 6749 34161 6783
rect 34195 6749 34207 6783
rect 34149 6743 34207 6749
rect 34330 6740 34336 6792
rect 34388 6780 34394 6792
rect 34992 6780 35020 6820
rect 35710 6808 35716 6820
rect 35768 6808 35774 6860
rect 34388 6752 35020 6780
rect 35529 6783 35587 6789
rect 34388 6740 34394 6752
rect 35529 6749 35541 6783
rect 35575 6780 35587 6783
rect 35618 6780 35624 6792
rect 35575 6752 35624 6780
rect 35575 6749 35587 6752
rect 35529 6743 35587 6749
rect 35618 6740 35624 6752
rect 35676 6740 35682 6792
rect 36170 6780 36176 6792
rect 36131 6752 36176 6780
rect 36170 6740 36176 6752
rect 36228 6740 36234 6792
rect 36722 6740 36728 6792
rect 36780 6780 36786 6792
rect 36817 6783 36875 6789
rect 36817 6780 36829 6783
rect 36780 6752 36829 6780
rect 36780 6740 36786 6752
rect 36817 6749 36829 6752
rect 36863 6749 36875 6783
rect 36817 6743 36875 6749
rect 37458 6740 37464 6792
rect 37516 6780 37522 6792
rect 38013 6783 38071 6789
rect 38013 6780 38025 6783
rect 37516 6752 38025 6780
rect 37516 6740 37522 6752
rect 38013 6749 38025 6752
rect 38059 6749 38071 6783
rect 38013 6743 38071 6749
rect 30282 6712 30288 6724
rect 23860 6684 26924 6712
rect 27738 6684 30288 6712
rect 14240 6616 14596 6644
rect 14240 6604 14246 6616
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18693 6647 18751 6653
rect 18693 6644 18705 6647
rect 18564 6616 18705 6644
rect 18564 6604 18570 6616
rect 18693 6613 18705 6616
rect 18739 6613 18751 6647
rect 18693 6607 18751 6613
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 19392 6616 19625 6644
rect 19392 6604 19398 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 20990 6604 20996 6656
rect 21048 6644 21054 6656
rect 21358 6644 21364 6656
rect 21048 6616 21364 6644
rect 21048 6604 21054 6616
rect 21358 6604 21364 6616
rect 21416 6604 21422 6656
rect 22370 6604 22376 6656
rect 22428 6644 22434 6656
rect 23474 6644 23480 6656
rect 22428 6616 23480 6644
rect 22428 6604 22434 6616
rect 23474 6604 23480 6616
rect 23532 6604 23538 6656
rect 23937 6647 23995 6653
rect 23937 6613 23949 6647
rect 23983 6644 23995 6647
rect 24302 6644 24308 6656
rect 23983 6616 24308 6644
rect 23983 6613 23995 6616
rect 23937 6607 23995 6613
rect 24302 6604 24308 6616
rect 24360 6604 24366 6656
rect 24673 6647 24731 6653
rect 24673 6613 24685 6647
rect 24719 6644 24731 6647
rect 25130 6644 25136 6656
rect 24719 6616 25136 6644
rect 24719 6613 24731 6616
rect 24673 6607 24731 6613
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 25317 6647 25375 6653
rect 25317 6613 25329 6647
rect 25363 6644 25375 6647
rect 26510 6644 26516 6656
rect 25363 6616 26516 6644
rect 25363 6613 25375 6616
rect 25317 6607 25375 6613
rect 26510 6604 26516 6616
rect 26568 6604 26574 6656
rect 26896 6644 26924 6684
rect 30282 6672 30288 6684
rect 30340 6672 30346 6724
rect 32125 6715 32183 6721
rect 31404 6684 31708 6712
rect 31404 6644 31432 6684
rect 26896 6616 31432 6644
rect 31481 6647 31539 6653
rect 31481 6613 31493 6647
rect 31527 6644 31539 6647
rect 31570 6644 31576 6656
rect 31527 6616 31576 6644
rect 31527 6613 31539 6616
rect 31481 6607 31539 6613
rect 31570 6604 31576 6616
rect 31628 6604 31634 6656
rect 31680 6644 31708 6684
rect 32125 6681 32137 6715
rect 32171 6712 32183 6715
rect 32858 6712 32864 6724
rect 32171 6684 32864 6712
rect 32171 6681 32183 6684
rect 32125 6675 32183 6681
rect 32858 6672 32864 6684
rect 32916 6672 32922 6724
rect 36630 6712 36636 6724
rect 32968 6684 36636 6712
rect 32968 6644 32996 6684
rect 36630 6672 36636 6684
rect 36688 6672 36694 6724
rect 31680 6616 32996 6644
rect 33778 6604 33784 6656
rect 33836 6644 33842 6656
rect 34054 6644 34060 6656
rect 33836 6616 34060 6644
rect 33836 6604 33842 6616
rect 34054 6604 34060 6616
rect 34112 6604 34118 6656
rect 34238 6644 34244 6656
rect 34199 6616 34244 6644
rect 34238 6604 34244 6616
rect 34296 6604 34302 6656
rect 34698 6604 34704 6656
rect 34756 6644 34762 6656
rect 35434 6644 35440 6656
rect 34756 6616 35440 6644
rect 34756 6604 34762 6616
rect 35434 6604 35440 6616
rect 35492 6604 35498 6656
rect 35618 6644 35624 6656
rect 35579 6616 35624 6644
rect 35618 6604 35624 6616
rect 35676 6604 35682 6656
rect 35710 6604 35716 6656
rect 35768 6644 35774 6656
rect 36265 6647 36323 6653
rect 36265 6644 36277 6647
rect 35768 6616 36277 6644
rect 35768 6604 35774 6616
rect 36265 6613 36277 6616
rect 36311 6613 36323 6647
rect 36265 6607 36323 6613
rect 36446 6604 36452 6656
rect 36504 6644 36510 6656
rect 36909 6647 36967 6653
rect 36909 6644 36921 6647
rect 36504 6616 36921 6644
rect 36504 6604 36510 6616
rect 36909 6613 36921 6616
rect 36955 6613 36967 6647
rect 36909 6607 36967 6613
rect 38197 6647 38255 6653
rect 38197 6613 38209 6647
rect 38243 6644 38255 6647
rect 38286 6644 38292 6656
rect 38243 6616 38292 6644
rect 38243 6613 38255 6616
rect 38197 6607 38255 6613
rect 38286 6604 38292 6616
rect 38344 6604 38350 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 6454 6440 6460 6452
rect 3743 6412 6460 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 9398 6440 9404 6452
rect 7208 6412 9404 6440
rect 3050 6372 3056 6384
rect 2608 6344 3056 6372
rect 2608 6316 2636 6344
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 3326 6332 3332 6384
rect 3384 6372 3390 6384
rect 5077 6375 5135 6381
rect 5077 6372 5089 6375
rect 3384 6344 5089 6372
rect 3384 6332 3390 6344
rect 5077 6341 5089 6344
rect 5123 6341 5135 6375
rect 5077 6335 5135 6341
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 5997 6375 6055 6381
rect 5997 6372 6009 6375
rect 5960 6344 6009 6372
rect 5960 6332 5966 6344
rect 5997 6341 6009 6344
rect 6043 6341 6055 6375
rect 5997 6335 6055 6341
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1544 6276 1593 6304
rect 1544 6264 1550 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2590 6304 2596 6316
rect 2363 6276 2596 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3142 6304 3148 6316
rect 3007 6276 3148 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6304 3663 6307
rect 4062 6304 4068 6316
rect 3651 6276 4068 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4246 6304 4252 6316
rect 4207 6276 4252 6304
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 6546 6304 6552 6316
rect 6507 6276 6552 6304
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7208 6313 7236 6412
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 11146 6440 11152 6452
rect 9548 6412 11008 6440
rect 11107 6412 11152 6440
rect 9548 6400 9554 6412
rect 7469 6375 7527 6381
rect 7469 6341 7481 6375
rect 7515 6372 7527 6375
rect 7742 6372 7748 6384
rect 7515 6344 7748 6372
rect 7515 6341 7527 6344
rect 7469 6335 7527 6341
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 8754 6372 8760 6384
rect 8694 6344 8760 6372
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 9416 6313 9444 6400
rect 9677 6375 9735 6381
rect 9677 6341 9689 6375
rect 9723 6372 9735 6375
rect 9950 6372 9956 6384
rect 9723 6344 9956 6372
rect 9723 6341 9735 6344
rect 9677 6335 9735 6341
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 10318 6332 10324 6384
rect 10376 6332 10382 6384
rect 10980 6372 11008 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 13814 6440 13820 6452
rect 12544 6412 13820 6440
rect 11422 6372 11428 6384
rect 10980 6344 11428 6372
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 12066 6372 12072 6384
rect 11624 6344 12072 6372
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6880 6276 7205 6304
rect 6880 6264 6886 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11624 6304 11652 6344
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 12544 6381 12572 6412
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 14274 6400 14280 6452
rect 14332 6440 14338 6452
rect 19794 6440 19800 6452
rect 14332 6412 19800 6440
rect 14332 6400 14338 6412
rect 12529 6375 12587 6381
rect 12529 6341 12541 6375
rect 12575 6341 12587 6375
rect 14826 6372 14832 6384
rect 13754 6344 14832 6372
rect 12529 6335 12587 6341
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 15396 6381 15424 6412
rect 19794 6400 19800 6412
rect 19852 6400 19858 6452
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 22278 6440 22284 6452
rect 20496 6412 22284 6440
rect 20496 6400 20502 6412
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 22922 6440 22928 6452
rect 22480 6412 22928 6440
rect 15381 6375 15439 6381
rect 15381 6341 15393 6375
rect 15427 6341 15439 6375
rect 16482 6372 16488 6384
rect 15381 6335 15439 6341
rect 16040 6344 16488 6372
rect 11020 6276 11652 6304
rect 11020 6264 11026 6276
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 11756 6276 12265 6304
rect 11756 6264 11762 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 14734 6304 14740 6316
rect 14695 6276 14740 6304
rect 12253 6267 12311 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 16040 6304 16068 6344
rect 16482 6332 16488 6344
rect 16540 6332 16546 6384
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 16632 6344 17141 6372
rect 16632 6332 16638 6344
rect 17129 6341 17141 6344
rect 17175 6341 17187 6375
rect 18874 6372 18880 6384
rect 17129 6335 17187 6341
rect 17880 6344 18880 6372
rect 15068 6276 16068 6304
rect 16132 6276 16896 6304
rect 15068 6264 15074 6276
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4798 6236 4804 6248
rect 4387 6208 4804 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 6730 6236 6736 6248
rect 5031 6208 5948 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 2409 6171 2467 6177
rect 2409 6137 2421 6171
rect 2455 6168 2467 6171
rect 5442 6168 5448 6180
rect 2455 6140 5448 6168
rect 2455 6137 2467 6140
rect 2409 6131 2467 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5920 6168 5948 6208
rect 6104 6208 6736 6236
rect 6104 6168 6132 6208
rect 6730 6196 6736 6208
rect 6788 6236 6794 6248
rect 6788 6208 13584 6236
rect 6788 6196 6794 6208
rect 5920 6140 6132 6168
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6168 6699 6171
rect 6822 6168 6828 6180
rect 6687 6140 6828 6168
rect 6687 6137 6699 6140
rect 6641 6131 6699 6137
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 8864 6140 9536 6168
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6100 3111 6103
rect 3602 6100 3608 6112
rect 3099 6072 3608 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 4982 6100 4988 6112
rect 4488 6072 4988 6100
rect 4488 6060 4494 6072
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 8864 6100 8892 6140
rect 5408 6072 8892 6100
rect 8941 6103 8999 6109
rect 5408 6060 5414 6072
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9122 6100 9128 6112
rect 8987 6072 9128 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9508 6100 9536 6140
rect 10686 6128 10692 6180
rect 10744 6168 10750 6180
rect 13556 6168 13584 6208
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 14148 6208 14289 6236
rect 14148 6196 14154 6208
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 16132 6236 16160 6276
rect 14277 6199 14335 6205
rect 14384 6208 16160 6236
rect 16209 6239 16267 6245
rect 14384 6168 14412 6208
rect 16209 6205 16221 6239
rect 16255 6236 16267 6239
rect 16298 6236 16304 6248
rect 16255 6208 16304 6236
rect 16255 6205 16267 6208
rect 16209 6199 16267 6205
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 16868 6236 16896 6276
rect 17034 6236 17040 6248
rect 16868 6208 17040 6236
rect 17034 6196 17040 6208
rect 17092 6196 17098 6248
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 17184 6208 17325 6236
rect 17184 6196 17190 6208
rect 17313 6205 17325 6208
rect 17359 6236 17371 6239
rect 17586 6236 17592 6248
rect 17359 6208 17592 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 17880 6168 17908 6344
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 20070 6372 20076 6384
rect 20010 6344 20076 6372
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 22480 6372 22508 6412
rect 22922 6400 22928 6412
rect 22980 6400 22986 6452
rect 23014 6400 23020 6452
rect 23072 6440 23078 6452
rect 23753 6443 23811 6449
rect 23753 6440 23765 6443
rect 23072 6412 23765 6440
rect 23072 6400 23078 6412
rect 23753 6409 23765 6412
rect 23799 6409 23811 6443
rect 23753 6403 23811 6409
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 26602 6440 26608 6452
rect 25280 6412 26608 6440
rect 25280 6400 25286 6412
rect 26602 6400 26608 6412
rect 26660 6400 26666 6452
rect 28258 6400 28264 6452
rect 28316 6440 28322 6452
rect 28902 6440 28908 6452
rect 28316 6412 28908 6440
rect 28316 6400 28322 6412
rect 28902 6400 28908 6412
rect 28960 6400 28966 6452
rect 29178 6400 29184 6452
rect 29236 6440 29242 6452
rect 29822 6440 29828 6452
rect 29236 6412 29828 6440
rect 29236 6400 29242 6412
rect 29822 6400 29828 6412
rect 29880 6400 29886 6452
rect 36173 6443 36231 6449
rect 36173 6440 36185 6443
rect 30024 6412 36185 6440
rect 24486 6372 24492 6384
rect 21008 6344 22508 6372
rect 23506 6344 24492 6372
rect 20346 6264 20352 6316
rect 20404 6304 20410 6316
rect 21008 6313 21036 6344
rect 24486 6332 24492 6344
rect 24544 6332 24550 6384
rect 27430 6372 27436 6384
rect 26988 6344 27436 6372
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 20404 6276 21005 6304
rect 20404 6264 20410 6276
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 25590 6264 25596 6316
rect 25648 6264 25654 6316
rect 26142 6264 26148 6316
rect 26200 6304 26206 6316
rect 26421 6307 26479 6313
rect 26421 6304 26433 6307
rect 26200 6276 26433 6304
rect 26200 6264 26206 6276
rect 26421 6273 26433 6276
rect 26467 6273 26479 6307
rect 26421 6267 26479 6273
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18782 6236 18788 6248
rect 18555 6208 18644 6236
rect 18743 6208 18788 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 10744 6140 11468 6168
rect 13556 6140 14412 6168
rect 14752 6140 17908 6168
rect 10744 6128 10750 6140
rect 11330 6100 11336 6112
rect 9508 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 11440 6100 11468 6140
rect 14752 6100 14780 6140
rect 11440 6072 14780 6100
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 14884 6072 14929 6100
rect 14884 6060 14890 6072
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 17954 6100 17960 6112
rect 15160 6072 17960 6100
rect 15160 6060 15166 6072
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 18616 6100 18644 6208
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 20530 6236 20536 6248
rect 18932 6208 19840 6236
rect 20491 6208 20536 6236
rect 18932 6196 18938 6208
rect 19812 6168 19840 6208
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 22002 6236 22008 6248
rect 20680 6208 21864 6236
rect 21963 6208 22008 6236
rect 20680 6196 20686 6208
rect 21726 6168 21732 6180
rect 19812 6140 21732 6168
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 21836 6168 21864 6208
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 22281 6239 22339 6245
rect 22281 6236 22293 6239
rect 22112 6208 22293 6236
rect 22112 6168 22140 6208
rect 22281 6205 22293 6208
rect 22327 6205 22339 6239
rect 22281 6199 22339 6205
rect 22370 6196 22376 6248
rect 22428 6236 22434 6248
rect 23658 6236 23664 6248
rect 22428 6208 23664 6236
rect 22428 6196 22434 6208
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 24210 6236 24216 6248
rect 24171 6208 24216 6236
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 24320 6208 24501 6236
rect 24320 6168 24348 6208
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 26988 6236 27016 6344
rect 27430 6332 27436 6344
rect 27488 6332 27494 6384
rect 30024 6372 30052 6412
rect 36173 6409 36185 6412
rect 36219 6409 36231 6443
rect 36173 6403 36231 6409
rect 36538 6400 36544 6452
rect 36596 6440 36602 6452
rect 36817 6443 36875 6449
rect 36817 6440 36829 6443
rect 36596 6412 36829 6440
rect 36596 6400 36602 6412
rect 36817 6409 36829 6412
rect 36863 6409 36875 6443
rect 36817 6403 36875 6409
rect 32030 6372 32036 6384
rect 28658 6344 30052 6372
rect 30866 6344 32036 6372
rect 32030 6332 32036 6344
rect 32088 6332 32094 6384
rect 32306 6372 32312 6384
rect 32267 6344 32312 6372
rect 32306 6332 32312 6344
rect 32364 6332 32370 6384
rect 34034 6375 34092 6381
rect 34034 6372 34046 6375
rect 33796 6344 34046 6372
rect 33796 6316 33824 6344
rect 34034 6341 34046 6344
rect 34080 6341 34092 6375
rect 34034 6335 34092 6341
rect 34422 6332 34428 6384
rect 34480 6372 34486 6384
rect 34480 6344 36768 6372
rect 34480 6332 34486 6344
rect 27154 6304 27160 6316
rect 27115 6276 27160 6304
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 29362 6304 29368 6316
rect 29323 6276 29368 6304
rect 29362 6264 29368 6276
rect 29420 6264 29426 6316
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 31938 6304 31944 6316
rect 31803 6276 31944 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 31938 6264 31944 6276
rect 31996 6264 32002 6316
rect 33502 6304 33508 6316
rect 33463 6276 33508 6304
rect 33502 6264 33508 6276
rect 33560 6264 33566 6316
rect 33778 6264 33784 6316
rect 33836 6264 33842 6316
rect 36078 6304 36084 6316
rect 36039 6276 36084 6304
rect 36078 6264 36084 6276
rect 36136 6264 36142 6316
rect 36740 6313 36768 6344
rect 36725 6307 36783 6313
rect 36725 6273 36737 6307
rect 36771 6273 36783 6307
rect 36725 6267 36783 6273
rect 38105 6307 38163 6313
rect 38105 6273 38117 6307
rect 38151 6273 38163 6307
rect 38105 6267 38163 6273
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 25188 6208 27016 6236
rect 27080 6208 27445 6236
rect 25188 6196 25194 6208
rect 21836 6140 22140 6168
rect 23308 6140 24348 6168
rect 20714 6100 20720 6112
rect 18616 6072 20720 6100
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 21085 6103 21143 6109
rect 21085 6069 21097 6103
rect 21131 6100 21143 6103
rect 22094 6100 22100 6112
rect 21131 6072 22100 6100
rect 21131 6069 21143 6072
rect 21085 6063 21143 6069
rect 22094 6060 22100 6072
rect 22152 6060 22158 6112
rect 22278 6060 22284 6112
rect 22336 6100 22342 6112
rect 23308 6100 23336 6140
rect 26142 6128 26148 6180
rect 26200 6168 26206 6180
rect 27080 6168 27108 6208
rect 27433 6205 27445 6208
rect 27479 6205 27491 6239
rect 27433 6199 27491 6205
rect 27522 6196 27528 6248
rect 27580 6236 27586 6248
rect 29178 6236 29184 6248
rect 27580 6208 29184 6236
rect 27580 6196 27586 6208
rect 29178 6196 29184 6208
rect 29236 6196 29242 6248
rect 29641 6239 29699 6245
rect 29641 6205 29653 6239
rect 29687 6236 29699 6239
rect 31294 6236 31300 6248
rect 29687 6208 31300 6236
rect 29687 6205 29699 6208
rect 29641 6199 29699 6205
rect 31294 6196 31300 6208
rect 31352 6196 31358 6248
rect 32214 6236 32220 6248
rect 32127 6208 32220 6236
rect 32214 6196 32220 6208
rect 32272 6196 32278 6248
rect 32490 6236 32496 6248
rect 32451 6208 32496 6236
rect 32490 6196 32496 6208
rect 32548 6196 32554 6248
rect 33520 6236 33548 6264
rect 33965 6239 34023 6245
rect 33965 6236 33977 6239
rect 33520 6208 33977 6236
rect 33965 6205 33977 6208
rect 34011 6236 34023 6239
rect 34146 6236 34152 6248
rect 34011 6208 34152 6236
rect 34011 6205 34023 6208
rect 33965 6199 34023 6205
rect 34146 6196 34152 6208
rect 34204 6196 34210 6248
rect 34241 6239 34299 6245
rect 34241 6205 34253 6239
rect 34287 6205 34299 6239
rect 35434 6236 35440 6248
rect 35395 6208 35440 6236
rect 34241 6199 34299 6205
rect 26200 6140 27108 6168
rect 26200 6128 26206 6140
rect 30650 6128 30656 6180
rect 30708 6168 30714 6180
rect 32232 6168 32260 6196
rect 34256 6168 34284 6199
rect 35434 6196 35440 6208
rect 35492 6196 35498 6248
rect 35710 6196 35716 6248
rect 35768 6236 35774 6248
rect 38120 6236 38148 6267
rect 35768 6208 38148 6236
rect 35768 6196 35774 6208
rect 30708 6140 31156 6168
rect 32232 6140 34284 6168
rect 30708 6128 30714 6140
rect 22336 6072 23336 6100
rect 22336 6060 22342 6072
rect 23474 6060 23480 6112
rect 23532 6100 23538 6112
rect 25961 6103 26019 6109
rect 25961 6100 25973 6103
rect 23532 6072 25973 6100
rect 23532 6060 23538 6072
rect 25961 6069 25973 6072
rect 26007 6069 26019 6103
rect 25961 6063 26019 6069
rect 26513 6103 26571 6109
rect 26513 6069 26525 6103
rect 26559 6100 26571 6103
rect 30098 6100 30104 6112
rect 26559 6072 30104 6100
rect 26559 6069 26571 6072
rect 26513 6063 26571 6069
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 31128 6109 31156 6140
rect 31113 6103 31171 6109
rect 31113 6069 31125 6103
rect 31159 6069 31171 6103
rect 31570 6100 31576 6112
rect 31531 6072 31576 6100
rect 31113 6063 31171 6069
rect 31570 6060 31576 6072
rect 31628 6060 31634 6112
rect 31754 6060 31760 6112
rect 31812 6100 31818 6112
rect 35618 6100 35624 6112
rect 31812 6072 35624 6100
rect 31812 6060 31818 6072
rect 35618 6060 35624 6072
rect 35676 6060 35682 6112
rect 38194 6100 38200 6112
rect 38155 6072 38200 6100
rect 38194 6060 38200 6072
rect 38252 6060 38258 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 4246 5896 4252 5908
rect 2648 5868 4252 5896
rect 2648 5856 2654 5868
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 7088 5899 7146 5905
rect 7088 5896 7100 5899
rect 4488 5868 7100 5896
rect 4488 5856 4494 5868
rect 7088 5865 7100 5868
rect 7134 5896 7146 5899
rect 7834 5896 7840 5908
rect 7134 5868 7840 5896
rect 7134 5865 7146 5868
rect 7088 5859 7146 5865
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 8128 5868 19748 5896
rect 1854 5828 1860 5840
rect 1815 5800 1860 5828
rect 1854 5788 1860 5800
rect 1912 5788 1918 5840
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5828 3387 5831
rect 3878 5828 3884 5840
rect 3375 5800 3884 5828
rect 3375 5797 3387 5800
rect 3329 5791 3387 5797
rect 3878 5788 3884 5800
rect 3936 5788 3942 5840
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 5810 5828 5816 5840
rect 4856 5800 5816 5828
rect 4856 5788 4862 5800
rect 5810 5788 5816 5800
rect 5868 5828 5874 5840
rect 6546 5828 6552 5840
rect 5868 5800 6552 5828
rect 5868 5788 5874 5800
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 8128 5760 8156 5868
rect 8573 5831 8631 5837
rect 8573 5797 8585 5831
rect 8619 5828 8631 5831
rect 8662 5828 8668 5840
rect 8619 5800 8668 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 11241 5831 11299 5837
rect 11241 5797 11253 5831
rect 11287 5828 11299 5831
rect 11422 5828 11428 5840
rect 11287 5800 11428 5828
rect 11287 5797 11299 5800
rect 11241 5791 11299 5797
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 11606 5788 11612 5840
rect 11664 5828 11670 5840
rect 16390 5828 16396 5840
rect 11664 5800 11836 5828
rect 16351 5800 16396 5828
rect 11664 5788 11670 5800
rect 2740 5732 8156 5760
rect 2740 5720 2746 5732
rect 8294 5720 8300 5772
rect 8352 5720 8358 5772
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 9456 5732 9505 5760
rect 9456 5720 9462 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 11698 5760 11704 5772
rect 9824 5732 9869 5760
rect 11659 5732 11704 5760
rect 9824 5720 9830 5732
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 11808 5760 11836 5800
rect 16390 5788 16396 5800
rect 16448 5788 16454 5840
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 11808 5732 11989 5760
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 16298 5760 16304 5772
rect 14691 5732 16304 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 16298 5720 16304 5732
rect 16356 5760 16362 5772
rect 16850 5760 16856 5772
rect 16356 5732 16856 5760
rect 16356 5720 16362 5732
rect 16850 5720 16856 5732
rect 16908 5760 16914 5772
rect 17126 5760 17132 5772
rect 16908 5732 17132 5760
rect 16908 5720 16914 5732
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 18782 5760 18788 5772
rect 17276 5732 18788 5760
rect 17276 5720 17282 5732
rect 18782 5720 18788 5732
rect 18840 5720 18846 5772
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 1360 5664 2329 5692
rect 1360 5652 1366 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 2317 5655 2375 5661
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 4246 5692 4252 5704
rect 4207 5664 4252 5692
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6788 5664 6837 5692
rect 6788 5652 6794 5664
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8312 5692 8340 5720
rect 16574 5692 16580 5704
rect 8312 5664 9536 5692
rect 16054 5664 16580 5692
rect 1670 5624 1676 5636
rect 1631 5596 1676 5624
rect 1670 5584 1676 5596
rect 1728 5584 1734 5636
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 5350 5624 5356 5636
rect 4212 5596 5356 5624
rect 4212 5584 4218 5596
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 6362 5624 6368 5636
rect 5500 5596 5545 5624
rect 6323 5596 6368 5624
rect 5500 5584 5506 5596
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 7374 5624 7380 5636
rect 6604 5596 7380 5624
rect 6604 5584 6610 5596
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 9508 5624 9536 5664
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 19720 5701 19748 5868
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 22646 5896 22652 5908
rect 20588 5868 22652 5896
rect 20588 5856 20594 5868
rect 22646 5856 22652 5868
rect 22704 5856 22710 5908
rect 22830 5856 22836 5908
rect 22888 5896 22894 5908
rect 22888 5868 31064 5896
rect 22888 5856 22894 5868
rect 21726 5788 21732 5840
rect 21784 5828 21790 5840
rect 28629 5831 28687 5837
rect 21784 5800 25176 5828
rect 21784 5788 21790 5800
rect 20441 5763 20499 5769
rect 20441 5729 20453 5763
rect 20487 5760 20499 5763
rect 20714 5760 20720 5772
rect 20487 5732 20720 5760
rect 20487 5729 20499 5732
rect 20441 5723 20499 5729
rect 20714 5720 20720 5732
rect 20772 5760 20778 5772
rect 22002 5760 22008 5772
rect 20772 5732 22008 5760
rect 20772 5720 20778 5732
rect 22002 5720 22008 5732
rect 22060 5760 22066 5772
rect 23661 5763 23719 5769
rect 23661 5760 23673 5763
rect 22060 5732 23673 5760
rect 22060 5720 22066 5732
rect 23661 5729 23673 5732
rect 23707 5760 23719 5763
rect 24210 5760 24216 5772
rect 23707 5732 24216 5760
rect 23707 5729 23719 5732
rect 23661 5723 23719 5729
rect 24210 5720 24216 5732
rect 24268 5720 24274 5772
rect 25148 5769 25176 5800
rect 28629 5797 28641 5831
rect 28675 5828 28687 5831
rect 31036 5828 31064 5868
rect 32306 5856 32312 5908
rect 32364 5896 32370 5908
rect 35621 5899 35679 5905
rect 35621 5896 35633 5899
rect 32364 5868 35633 5896
rect 32364 5856 32370 5868
rect 35621 5865 35633 5868
rect 35667 5865 35679 5899
rect 35621 5859 35679 5865
rect 31754 5828 31760 5840
rect 28675 5800 29868 5828
rect 31036 5800 31760 5828
rect 28675 5797 28687 5800
rect 28629 5791 28687 5797
rect 25133 5763 25191 5769
rect 25133 5729 25145 5763
rect 25179 5729 25191 5763
rect 25133 5723 25191 5729
rect 26145 5763 26203 5769
rect 26145 5729 26157 5763
rect 26191 5760 26203 5763
rect 27154 5760 27160 5772
rect 26191 5732 27160 5760
rect 26191 5729 26203 5732
rect 26145 5723 26203 5729
rect 27154 5720 27160 5732
rect 27212 5720 27218 5772
rect 27430 5720 27436 5772
rect 27488 5760 27494 5772
rect 27488 5732 29316 5760
rect 27488 5720 27494 5732
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 20346 5692 20352 5704
rect 19705 5655 19763 5661
rect 19812 5664 20352 5692
rect 9508 5596 10180 5624
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 1544 5528 2513 5556
rect 1544 5516 1550 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 2501 5519 2559 5525
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 7742 5556 7748 5568
rect 4387 5528 7748 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 9674 5556 9680 5568
rect 7892 5528 9680 5556
rect 7892 5516 7898 5528
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 10152 5556 10180 5596
rect 10226 5584 10232 5636
rect 10284 5584 10290 5636
rect 12710 5584 12716 5636
rect 12768 5584 12774 5636
rect 13725 5627 13783 5633
rect 13725 5593 13737 5627
rect 13771 5624 13783 5627
rect 14090 5624 14096 5636
rect 13771 5596 14096 5624
rect 13771 5593 13783 5596
rect 13725 5587 13783 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 14921 5627 14979 5633
rect 14921 5593 14933 5627
rect 14967 5624 14979 5627
rect 15010 5624 15016 5636
rect 14967 5596 15016 5624
rect 14967 5593 14979 5596
rect 14921 5587 14979 5593
rect 15010 5584 15016 5596
rect 15068 5584 15074 5636
rect 17129 5627 17187 5633
rect 17129 5593 17141 5627
rect 17175 5624 17187 5627
rect 17218 5624 17224 5636
rect 17175 5596 17224 5624
rect 17175 5593 17187 5596
rect 17129 5587 17187 5593
rect 17218 5584 17224 5596
rect 17276 5624 17282 5636
rect 17402 5624 17408 5636
rect 17276 5596 17408 5624
rect 17276 5584 17282 5596
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 18138 5584 18144 5636
rect 18196 5584 18202 5636
rect 18874 5624 18880 5636
rect 18835 5596 18880 5624
rect 18874 5584 18880 5596
rect 18932 5584 18938 5636
rect 11054 5556 11060 5568
rect 10152 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 19812 5556 19840 5664
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 22830 5692 22836 5704
rect 21850 5664 22836 5692
rect 22830 5652 22836 5664
rect 22888 5652 22894 5704
rect 22925 5695 22983 5701
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 24762 5692 24768 5704
rect 22971 5664 24768 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 20438 5624 20444 5636
rect 19904 5596 20444 5624
rect 19904 5565 19932 5596
rect 20438 5584 20444 5596
rect 20496 5584 20502 5636
rect 20717 5627 20775 5633
rect 20717 5593 20729 5627
rect 20763 5624 20775 5627
rect 20990 5624 20996 5636
rect 20763 5596 20996 5624
rect 20763 5593 20775 5596
rect 20717 5587 20775 5593
rect 20990 5584 20996 5596
rect 21048 5584 21054 5636
rect 22186 5584 22192 5636
rect 22244 5624 22250 5636
rect 22465 5627 22523 5633
rect 22465 5624 22477 5627
rect 22244 5596 22477 5624
rect 22244 5584 22250 5596
rect 22465 5593 22477 5596
rect 22511 5593 22523 5627
rect 22465 5587 22523 5593
rect 14792 5528 19840 5556
rect 19889 5559 19947 5565
rect 14792 5516 14798 5528
rect 19889 5525 19901 5559
rect 19935 5525 19947 5559
rect 19889 5519 19947 5525
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 22940 5556 22968 5655
rect 24762 5652 24768 5664
rect 24820 5652 24826 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 24872 5624 24900 5655
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 28813 5695 28871 5701
rect 28813 5692 28825 5695
rect 27764 5664 28825 5692
rect 27764 5652 27770 5664
rect 28813 5661 28825 5664
rect 28859 5661 28871 5695
rect 29288 5692 29316 5732
rect 29362 5720 29368 5772
rect 29420 5760 29426 5772
rect 29733 5763 29791 5769
rect 29733 5760 29745 5763
rect 29420 5732 29745 5760
rect 29420 5720 29426 5732
rect 29733 5729 29745 5732
rect 29779 5729 29791 5763
rect 29840 5760 29868 5800
rect 31754 5788 31760 5800
rect 31812 5788 31818 5840
rect 33042 5828 33048 5840
rect 31864 5800 33048 5828
rect 31864 5760 31892 5800
rect 33042 5788 33048 5800
rect 33100 5788 33106 5840
rect 33134 5788 33140 5840
rect 33192 5828 33198 5840
rect 33778 5828 33784 5840
rect 33192 5800 33784 5828
rect 33192 5788 33198 5800
rect 33778 5788 33784 5800
rect 33836 5828 33842 5840
rect 34149 5831 34207 5837
rect 34149 5828 34161 5831
rect 33836 5800 34161 5828
rect 33836 5788 33842 5800
rect 34149 5797 34161 5800
rect 34195 5797 34207 5831
rect 34149 5791 34207 5797
rect 34698 5788 34704 5840
rect 34756 5828 34762 5840
rect 34977 5831 35035 5837
rect 34977 5828 34989 5831
rect 34756 5800 34989 5828
rect 34756 5788 34762 5800
rect 34977 5797 34989 5800
rect 35023 5797 35035 5831
rect 34977 5791 35035 5797
rect 35066 5788 35072 5840
rect 35124 5828 35130 5840
rect 36265 5831 36323 5837
rect 36265 5828 36277 5831
rect 35124 5800 36277 5828
rect 35124 5788 35130 5800
rect 36265 5797 36277 5800
rect 36311 5797 36323 5831
rect 36265 5791 36323 5797
rect 29840 5732 31892 5760
rect 32033 5763 32091 5769
rect 29733 5723 29791 5729
rect 32033 5729 32045 5763
rect 32079 5760 32091 5763
rect 35434 5760 35440 5772
rect 32079 5732 35440 5760
rect 32079 5729 32091 5732
rect 32033 5723 32091 5729
rect 35434 5720 35440 5732
rect 35492 5720 35498 5772
rect 29638 5692 29644 5704
rect 29288 5664 29644 5692
rect 28813 5655 28871 5661
rect 29638 5652 29644 5664
rect 29696 5652 29702 5704
rect 31110 5652 31116 5704
rect 31168 5652 31174 5704
rect 34514 5652 34520 5704
rect 34572 5692 34578 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34572 5664 34897 5692
rect 34572 5652 34578 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35529 5695 35587 5701
rect 35529 5661 35541 5695
rect 35575 5661 35587 5695
rect 35529 5655 35587 5661
rect 26326 5624 26332 5636
rect 24872 5596 26332 5624
rect 26326 5584 26332 5596
rect 26384 5584 26390 5636
rect 26421 5627 26479 5633
rect 26421 5593 26433 5627
rect 26467 5624 26479 5627
rect 26694 5624 26700 5636
rect 26467 5596 26700 5624
rect 26467 5593 26479 5596
rect 26421 5587 26479 5593
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 28074 5624 28080 5636
rect 27646 5596 28080 5624
rect 28074 5584 28080 5596
rect 28132 5584 28138 5636
rect 28169 5627 28227 5633
rect 28169 5593 28181 5627
rect 28215 5624 28227 5627
rect 28258 5624 28264 5636
rect 28215 5596 28264 5624
rect 28215 5593 28227 5596
rect 28169 5587 28227 5593
rect 28258 5584 28264 5596
rect 28316 5584 28322 5636
rect 30009 5627 30067 5633
rect 30009 5593 30021 5627
rect 30055 5624 30067 5627
rect 30282 5624 30288 5636
rect 30055 5596 30288 5624
rect 30055 5593 30067 5596
rect 30009 5587 30067 5593
rect 30282 5584 30288 5596
rect 30340 5584 30346 5636
rect 32125 5627 32183 5633
rect 32125 5624 32137 5627
rect 31312 5596 32137 5624
rect 20036 5528 22968 5556
rect 20036 5516 20042 5528
rect 23934 5516 23940 5568
rect 23992 5556 23998 5568
rect 26142 5556 26148 5568
rect 23992 5528 26148 5556
rect 23992 5516 23998 5528
rect 26142 5516 26148 5528
rect 26200 5516 26206 5568
rect 26510 5516 26516 5568
rect 26568 5556 26574 5568
rect 31312 5556 31340 5596
rect 32125 5593 32137 5596
rect 32171 5593 32183 5627
rect 32125 5587 32183 5593
rect 33045 5627 33103 5633
rect 33045 5593 33057 5627
rect 33091 5593 33103 5627
rect 33045 5587 33103 5593
rect 33597 5627 33655 5633
rect 33597 5593 33609 5627
rect 33643 5593 33655 5627
rect 33597 5587 33655 5593
rect 33689 5627 33747 5633
rect 33689 5593 33701 5627
rect 33735 5624 33747 5627
rect 35342 5624 35348 5636
rect 33735 5596 35348 5624
rect 33735 5593 33747 5596
rect 33689 5587 33747 5593
rect 26568 5528 31340 5556
rect 26568 5516 26574 5528
rect 31386 5516 31392 5568
rect 31444 5556 31450 5568
rect 31481 5559 31539 5565
rect 31481 5556 31493 5559
rect 31444 5528 31493 5556
rect 31444 5516 31450 5528
rect 31481 5525 31493 5528
rect 31527 5525 31539 5559
rect 31481 5519 31539 5525
rect 31570 5516 31576 5568
rect 31628 5556 31634 5568
rect 32490 5556 32496 5568
rect 31628 5528 32496 5556
rect 31628 5516 31634 5528
rect 32490 5516 32496 5528
rect 32548 5556 32554 5568
rect 33060 5556 33088 5587
rect 32548 5528 33088 5556
rect 33612 5556 33640 5587
rect 35342 5584 35348 5596
rect 35400 5584 35406 5636
rect 35544 5568 35572 5655
rect 35618 5652 35624 5704
rect 35676 5692 35682 5704
rect 36173 5695 36231 5701
rect 36173 5692 36185 5695
rect 35676 5664 36185 5692
rect 35676 5652 35682 5664
rect 36173 5661 36185 5664
rect 36219 5661 36231 5695
rect 37274 5692 37280 5704
rect 37235 5664 37280 5692
rect 36173 5655 36231 5661
rect 37274 5652 37280 5664
rect 37332 5652 37338 5704
rect 37366 5652 37372 5704
rect 37424 5692 37430 5704
rect 38013 5695 38071 5701
rect 38013 5692 38025 5695
rect 37424 5664 38025 5692
rect 37424 5652 37430 5664
rect 38013 5661 38025 5664
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 34698 5556 34704 5568
rect 33612 5528 34704 5556
rect 32548 5516 32554 5528
rect 34698 5516 34704 5528
rect 34756 5516 34762 5568
rect 35526 5516 35532 5568
rect 35584 5516 35590 5568
rect 37458 5556 37464 5568
rect 37419 5528 37464 5556
rect 37458 5516 37464 5528
rect 37516 5516 37522 5568
rect 38010 5516 38016 5568
rect 38068 5556 38074 5568
rect 38197 5559 38255 5565
rect 38197 5556 38209 5559
rect 38068 5528 38209 5556
rect 38068 5516 38074 5528
rect 38197 5525 38209 5528
rect 38243 5525 38255 5559
rect 38197 5519 38255 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 6822 5352 6828 5364
rect 3384 5324 6828 5352
rect 3384 5312 3390 5324
rect 3510 5284 3516 5296
rect 3471 5256 3516 5284
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 5000 5293 5028 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7374 5312 7380 5364
rect 7432 5352 7438 5364
rect 8294 5352 8300 5364
rect 7432 5324 8300 5352
rect 7432 5312 7438 5324
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 18874 5352 18880 5364
rect 8444 5324 10088 5352
rect 8444 5312 8450 5324
rect 4985 5287 5043 5293
rect 4985 5253 4997 5287
rect 5031 5253 5043 5287
rect 4985 5247 5043 5253
rect 5077 5287 5135 5293
rect 5077 5253 5089 5287
rect 5123 5284 5135 5287
rect 5166 5284 5172 5296
rect 5123 5256 5172 5284
rect 5123 5253 5135 5256
rect 5077 5247 5135 5253
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 6917 5287 6975 5293
rect 5684 5256 5856 5284
rect 5684 5244 5690 5256
rect 1118 5176 1124 5228
rect 1176 5216 1182 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1176 5188 1593 5216
rect 1176 5176 1182 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 1581 5179 1639 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 5828 5216 5856 5256
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 9030 5284 9036 5296
rect 6963 5256 9036 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 9030 5244 9036 5256
rect 9088 5244 9094 5296
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 10060 5293 10088 5324
rect 15120 5324 18880 5352
rect 15120 5296 15148 5324
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19153 5355 19211 5361
rect 19153 5321 19165 5355
rect 19199 5352 19211 5355
rect 21082 5352 21088 5364
rect 19199 5324 21088 5352
rect 19199 5321 19211 5324
rect 19153 5315 19211 5321
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 26142 5312 26148 5364
rect 26200 5352 26206 5364
rect 29178 5352 29184 5364
rect 26200 5324 29184 5352
rect 26200 5312 26206 5324
rect 29178 5312 29184 5324
rect 29236 5312 29242 5364
rect 30742 5312 30748 5364
rect 30800 5352 30806 5364
rect 31570 5352 31576 5364
rect 30800 5324 31576 5352
rect 30800 5312 30806 5324
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 32122 5312 32128 5364
rect 32180 5352 32186 5364
rect 32180 5324 32996 5352
rect 32180 5312 32186 5324
rect 9953 5287 10011 5293
rect 9953 5284 9965 5287
rect 9180 5256 9965 5284
rect 9180 5244 9186 5256
rect 9953 5253 9965 5256
rect 9999 5253 10011 5287
rect 9953 5247 10011 5253
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5253 10103 5287
rect 10045 5247 10103 5253
rect 12618 5244 12624 5296
rect 12676 5244 12682 5296
rect 13262 5244 13268 5296
rect 13320 5284 13326 5296
rect 14550 5284 14556 5296
rect 13320 5256 14556 5284
rect 13320 5244 13326 5256
rect 14550 5244 14556 5256
rect 14608 5244 14614 5296
rect 14829 5287 14887 5293
rect 14829 5253 14841 5287
rect 14875 5284 14887 5287
rect 15102 5284 15108 5296
rect 14875 5256 15108 5284
rect 14875 5253 14887 5256
rect 14829 5247 14887 5253
rect 15102 5244 15108 5256
rect 15160 5244 15166 5296
rect 16114 5284 16120 5296
rect 16054 5256 16120 5284
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 18046 5244 18052 5296
rect 18104 5244 18110 5296
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5284 18843 5287
rect 19058 5284 19064 5296
rect 18831 5256 19064 5284
rect 18831 5253 18843 5256
rect 18785 5247 18843 5253
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 21100 5284 21128 5312
rect 20930 5256 21128 5284
rect 24486 5244 24492 5296
rect 24544 5284 24550 5296
rect 24581 5287 24639 5293
rect 24581 5284 24593 5287
rect 24544 5256 24593 5284
rect 24544 5244 24550 5256
rect 24581 5253 24593 5256
rect 24627 5253 24639 5287
rect 26050 5284 26056 5296
rect 25806 5256 26056 5284
rect 24581 5247 24639 5253
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 26418 5244 26424 5296
rect 26476 5284 26482 5296
rect 27433 5287 27491 5293
rect 27433 5284 27445 5287
rect 26476 5256 27445 5284
rect 26476 5244 26482 5256
rect 27433 5253 27445 5256
rect 27479 5253 27491 5287
rect 27433 5247 27491 5253
rect 28166 5244 28172 5296
rect 28224 5244 28230 5296
rect 30190 5284 30196 5296
rect 28736 5256 30196 5284
rect 6178 5216 6184 5228
rect 5828 5188 6184 5216
rect 6178 5176 6184 5188
rect 6236 5216 6242 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6236 5188 7573 5216
rect 6236 5176 6242 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 7561 5179 7619 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 3418 5148 3424 5160
rect 3379 5120 3424 5148
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 4448 5080 4476 5111
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4672 5120 5273 5148
rect 4672 5108 4678 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 7006 5148 7012 5160
rect 5408 5120 7012 5148
rect 5408 5108 5414 5120
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 7248 5132 7696 5148
rect 7745 5135 7803 5141
rect 7745 5132 7757 5135
rect 7248 5120 7757 5132
rect 7248 5108 7254 5120
rect 7668 5104 7757 5120
rect 7745 5101 7757 5104
rect 7791 5101 7803 5135
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 9214 5148 9220 5160
rect 8352 5120 9220 5148
rect 8352 5108 8358 5120
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9398 5148 9404 5160
rect 9359 5120 9404 5148
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 10962 5148 10968 5160
rect 10923 5120 10968 5148
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 13630 5148 13636 5160
rect 12023 5120 13636 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 13814 5148 13820 5160
rect 13771 5120 13820 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14332 5120 14565 5148
rect 14332 5108 14338 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 16758 5148 16764 5160
rect 14553 5111 14611 5117
rect 14660 5120 16436 5148
rect 16719 5120 16764 5148
rect 7745 5095 7803 5101
rect 5626 5080 5632 5092
rect 4448 5052 5632 5080
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 7834 5040 7840 5092
rect 7892 5080 7898 5092
rect 11514 5080 11520 5092
rect 7892 5052 11520 5080
rect 7892 5040 7898 5052
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 14090 5040 14096 5092
rect 14148 5080 14154 5092
rect 14660 5080 14688 5120
rect 16298 5080 16304 5092
rect 14148 5052 14688 5080
rect 16259 5052 16304 5080
rect 14148 5040 14154 5052
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 1302 4972 1308 5024
rect 1360 5012 1366 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 1360 4984 1777 5012
rect 1360 4972 1366 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 2498 5012 2504 5024
rect 2459 4984 2504 5012
rect 1765 4975 1823 4981
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 9858 5012 9864 5024
rect 4028 4984 9864 5012
rect 4028 4972 4034 4984
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 16206 5012 16212 5024
rect 11112 4984 16212 5012
rect 11112 4972 11118 4984
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 16408 5012 16436 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 17126 5108 17132 5160
rect 17184 5148 17190 5160
rect 19444 5148 19472 5179
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 21453 5219 21511 5225
rect 21453 5216 21465 5219
rect 21324 5188 21465 5216
rect 21324 5176 21330 5188
rect 21453 5185 21465 5188
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 23382 5176 23388 5228
rect 23440 5176 23446 5228
rect 17184 5120 19472 5148
rect 19705 5151 19763 5157
rect 17184 5108 17190 5120
rect 19705 5117 19717 5151
rect 19751 5148 19763 5151
rect 20990 5148 20996 5160
rect 19751 5120 20996 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 22002 5148 22008 5160
rect 21963 5120 22008 5148
rect 22002 5108 22008 5120
rect 22060 5108 22066 5160
rect 22281 5151 22339 5157
rect 22281 5117 22293 5151
rect 22327 5148 22339 5151
rect 24302 5148 24308 5160
rect 22327 5120 24164 5148
rect 24263 5120 24308 5148
rect 22327 5117 22339 5120
rect 22281 5111 22339 5117
rect 23753 5083 23811 5089
rect 23753 5049 23765 5083
rect 23799 5080 23811 5083
rect 23934 5080 23940 5092
rect 23799 5052 23940 5080
rect 23799 5049 23811 5052
rect 23753 5043 23811 5049
rect 23934 5040 23940 5052
rect 23992 5040 23998 5092
rect 17024 5015 17082 5021
rect 17024 5012 17036 5015
rect 16408 4984 17036 5012
rect 17024 4981 17036 4984
rect 17070 5012 17082 5015
rect 19426 5012 19432 5024
rect 17070 4984 19432 5012
rect 17070 4981 17082 4984
rect 17024 4975 17082 4981
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 21174 4972 21180 5024
rect 21232 5012 21238 5024
rect 22738 5012 22744 5024
rect 21232 4984 22744 5012
rect 21232 4972 21238 4984
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 24136 5012 24164 5120
rect 24302 5108 24308 5120
rect 24360 5108 24366 5160
rect 25222 5108 25228 5160
rect 25280 5148 25286 5160
rect 26329 5151 26387 5157
rect 26329 5148 26341 5151
rect 25280 5120 26341 5148
rect 25280 5108 25286 5120
rect 26329 5117 26341 5120
rect 26375 5117 26387 5151
rect 27154 5148 27160 5160
rect 27115 5120 27160 5148
rect 26329 5111 26387 5117
rect 27154 5108 27160 5120
rect 27212 5108 27218 5160
rect 28736 5148 28764 5256
rect 30190 5244 30196 5256
rect 30248 5244 30254 5296
rect 31846 5284 31852 5296
rect 31142 5256 31852 5284
rect 31846 5244 31852 5256
rect 31904 5244 31910 5296
rect 31938 5244 31944 5296
rect 31996 5284 32002 5296
rect 32309 5287 32367 5293
rect 32309 5284 32321 5287
rect 31996 5256 32321 5284
rect 31996 5244 32002 5256
rect 32309 5253 32321 5256
rect 32355 5253 32367 5287
rect 32968 5284 32996 5324
rect 33042 5312 33048 5364
rect 33100 5352 33106 5364
rect 33100 5324 35480 5352
rect 33100 5312 33106 5324
rect 33505 5287 33563 5293
rect 33505 5284 33517 5287
rect 32968 5256 33517 5284
rect 32309 5247 32367 5253
rect 33505 5253 33517 5256
rect 33551 5284 33563 5287
rect 33965 5287 34023 5293
rect 33965 5284 33977 5287
rect 33551 5256 33977 5284
rect 33551 5253 33563 5256
rect 33505 5247 33563 5253
rect 33965 5253 33977 5256
rect 34011 5253 34023 5287
rect 33965 5247 34023 5253
rect 34057 5287 34115 5293
rect 34057 5253 34069 5287
rect 34103 5284 34115 5287
rect 35066 5284 35072 5296
rect 34103 5256 35072 5284
rect 34103 5253 34115 5256
rect 34057 5247 34115 5253
rect 35066 5244 35072 5256
rect 35124 5244 35130 5296
rect 29178 5216 29184 5228
rect 29139 5188 29184 5216
rect 29178 5176 29184 5188
rect 29236 5176 29242 5228
rect 35452 5225 35480 5324
rect 35437 5219 35495 5225
rect 34808 5188 35112 5216
rect 29638 5148 29644 5160
rect 27264 5120 28764 5148
rect 29599 5120 29644 5148
rect 26510 5040 26516 5092
rect 26568 5080 26574 5092
rect 27264 5080 27292 5120
rect 29638 5108 29644 5120
rect 29696 5108 29702 5160
rect 29917 5151 29975 5157
rect 29917 5117 29929 5151
rect 29963 5148 29975 5151
rect 31386 5148 31392 5160
rect 29963 5120 31392 5148
rect 29963 5117 29975 5120
rect 29917 5111 29975 5117
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 31726 5120 32168 5148
rect 26568 5052 27292 5080
rect 26568 5040 26574 5052
rect 30926 5040 30932 5092
rect 30984 5080 30990 5092
rect 31726 5080 31754 5120
rect 30984 5052 31754 5080
rect 30984 5040 30990 5052
rect 25774 5012 25780 5024
rect 24136 4984 25780 5012
rect 25774 4972 25780 4984
rect 25832 4972 25838 5024
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 31389 5015 31447 5021
rect 31389 5012 31401 5015
rect 26752 4984 31401 5012
rect 26752 4972 26758 4984
rect 31389 4981 31401 4984
rect 31435 5012 31447 5015
rect 31754 5012 31760 5024
rect 31435 4984 31760 5012
rect 31435 4981 31447 4984
rect 31389 4975 31447 4981
rect 31754 4972 31760 4984
rect 31812 4972 31818 5024
rect 32140 5012 32168 5120
rect 32214 5108 32220 5160
rect 32272 5148 32278 5160
rect 32490 5148 32496 5160
rect 32272 5120 32317 5148
rect 32451 5120 32496 5148
rect 32272 5108 32278 5120
rect 32490 5108 32496 5120
rect 32548 5108 32554 5160
rect 32582 5108 32588 5160
rect 32640 5148 32646 5160
rect 34808 5148 34836 5188
rect 32640 5120 34836 5148
rect 32640 5108 32646 5120
rect 34882 5108 34888 5160
rect 34940 5148 34946 5160
rect 35084 5148 35112 5188
rect 35437 5185 35449 5219
rect 35483 5185 35495 5219
rect 35437 5179 35495 5185
rect 36633 5219 36691 5225
rect 36633 5185 36645 5219
rect 36679 5216 36691 5219
rect 38102 5216 38108 5228
rect 36679 5188 38108 5216
rect 36679 5185 36691 5188
rect 36633 5179 36691 5185
rect 38102 5176 38108 5188
rect 38160 5176 38166 5228
rect 37461 5151 37519 5157
rect 37461 5148 37473 5151
rect 34940 5120 34985 5148
rect 35084 5120 37473 5148
rect 34940 5108 34946 5120
rect 37461 5117 37473 5120
rect 37507 5117 37519 5151
rect 37461 5111 37519 5117
rect 37737 5151 37795 5157
rect 37737 5117 37749 5151
rect 37783 5148 37795 5151
rect 38562 5148 38568 5160
rect 37783 5120 38568 5148
rect 37783 5117 37795 5120
rect 37737 5111 37795 5117
rect 38562 5108 38568 5120
rect 38620 5108 38626 5160
rect 32306 5040 32312 5092
rect 32364 5080 32370 5092
rect 35529 5083 35587 5089
rect 35529 5080 35541 5083
rect 32364 5052 35541 5080
rect 32364 5040 32370 5052
rect 35529 5049 35541 5052
rect 35575 5049 35587 5083
rect 35529 5043 35587 5049
rect 35618 5012 35624 5024
rect 32140 4984 35624 5012
rect 35618 4972 35624 4984
rect 35676 4972 35682 5024
rect 36814 5012 36820 5024
rect 36775 4984 36820 5012
rect 36814 4972 36820 4984
rect 36872 4972 36878 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 842 4768 848 4820
rect 900 4808 906 4820
rect 1765 4811 1823 4817
rect 1765 4808 1777 4811
rect 900 4780 1777 4808
rect 900 4768 906 4780
rect 1765 4777 1777 4780
rect 1811 4777 1823 4811
rect 1765 4771 1823 4777
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 2501 4811 2559 4817
rect 2501 4808 2513 4811
rect 2280 4780 2513 4808
rect 2280 4768 2286 4780
rect 2501 4777 2513 4780
rect 2547 4777 2559 4811
rect 2501 4771 2559 4777
rect 4065 4811 4123 4817
rect 4065 4777 4077 4811
rect 4111 4808 4123 4811
rect 8202 4808 8208 4820
rect 4111 4780 8208 4808
rect 4111 4777 4123 4780
rect 4065 4771 4123 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 9766 4808 9772 4820
rect 8619 4780 9772 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 9916 4780 16160 4808
rect 9916 4768 9922 4780
rect 6365 4743 6423 4749
rect 6365 4709 6377 4743
rect 6411 4740 6423 4743
rect 6638 4740 6644 4752
rect 6411 4712 6644 4740
rect 6411 4709 6423 4712
rect 6365 4703 6423 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 16132 4740 16160 4780
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 16264 4780 16313 4808
rect 16264 4768 16270 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 17218 4808 17224 4820
rect 16301 4771 16359 4777
rect 16684 4780 17224 4808
rect 16574 4740 16580 4752
rect 16132 4712 16580 4740
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4663 4644 6776 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 6748 4616 6776 4644
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 7800 4644 8432 4672
rect 7800 4632 7806 4644
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 3050 4604 3056 4616
rect 2004 4576 2544 4604
rect 3011 4576 3056 4604
rect 2004 4564 2010 4576
rect 1670 4536 1676 4548
rect 1631 4508 1676 4536
rect 1670 4496 1676 4508
rect 1728 4496 1734 4548
rect 1854 4496 1860 4548
rect 1912 4536 1918 4548
rect 2409 4539 2467 4545
rect 2409 4536 2421 4539
rect 1912 4508 2421 4536
rect 1912 4496 1918 4508
rect 2409 4505 2421 4508
rect 2455 4505 2467 4539
rect 2516 4536 2544 4576
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4522 4604 4528 4616
rect 4019 4576 4528 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6788 4576 6837 4604
rect 6788 4564 6794 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 2516 4508 4200 4536
rect 2409 4499 2467 4505
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4172 4468 4200 4508
rect 4798 4496 4804 4548
rect 4856 4536 4862 4548
rect 4893 4539 4951 4545
rect 4893 4536 4905 4539
rect 4856 4508 4905 4536
rect 4856 4496 4862 4508
rect 4893 4505 4905 4508
rect 4939 4505 4951 4539
rect 7101 4539 7159 4545
rect 4893 4499 4951 4505
rect 5000 4508 5382 4536
rect 5000 4468 5028 4508
rect 7101 4505 7113 4539
rect 7147 4505 7159 4539
rect 7101 4499 7159 4505
rect 4172 4440 5028 4468
rect 7116 4468 7144 4499
rect 7558 4496 7564 4548
rect 7616 4496 7622 4548
rect 8404 4536 8432 4644
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9493 4675 9551 4681
rect 9493 4672 9505 4675
rect 8996 4644 9505 4672
rect 8996 4632 9002 4644
rect 9493 4641 9505 4644
rect 9539 4641 9551 4675
rect 9493 4635 9551 4641
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 9732 4644 13768 4672
rect 9732 4632 9738 4644
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11112 4576 11253 4604
rect 11112 4564 11118 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 13740 4604 13768 4644
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 16684 4672 16712 4780
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 21174 4808 21180 4820
rect 17368 4780 21180 4808
rect 17368 4768 17374 4780
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 21266 4768 21272 4820
rect 21324 4808 21330 4820
rect 22186 4808 22192 4820
rect 21324 4780 22192 4808
rect 21324 4768 21330 4780
rect 22186 4768 22192 4780
rect 22244 4768 22250 4820
rect 25958 4768 25964 4820
rect 26016 4808 26022 4820
rect 33778 4808 33784 4820
rect 26016 4780 29040 4808
rect 26016 4768 26022 4780
rect 24578 4740 24584 4752
rect 18156 4712 18736 4740
rect 13872 4644 16712 4672
rect 16853 4675 16911 4681
rect 13872 4632 13878 4644
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 17126 4672 17132 4684
rect 16899 4644 17132 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 17218 4632 17224 4684
rect 17276 4672 17282 4684
rect 18156 4672 18184 4712
rect 18322 4672 18328 4684
rect 17276 4644 18184 4672
rect 18248 4644 18328 4672
rect 17276 4632 17282 4644
rect 14090 4604 14096 4616
rect 13740 4576 14096 4604
rect 11241 4567 11299 4573
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14332 4576 14565 4604
rect 14332 4564 14338 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 18248 4590 18276 4644
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18708 4616 18736 4712
rect 22204 4712 24584 4740
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 21177 4675 21235 4681
rect 18932 4644 20760 4672
rect 18932 4632 18938 4644
rect 14553 4567 14611 4573
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 19242 4604 19248 4616
rect 18748 4576 19248 4604
rect 18748 4564 18754 4576
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 19978 4604 19984 4616
rect 19475 4576 19984 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 9214 4536 9220 4548
rect 8404 4508 9076 4536
rect 9175 4508 9220 4536
rect 8662 4468 8668 4480
rect 7116 4440 8668 4468
rect 8662 4428 8668 4440
rect 8720 4428 8726 4480
rect 9048 4468 9076 4508
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 9309 4539 9367 4545
rect 9309 4505 9321 4539
rect 9355 4505 9367 4539
rect 11514 4536 11520 4548
rect 11475 4508 11520 4536
rect 9309 4499 9367 4505
rect 9324 4468 9352 4499
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 12802 4536 12808 4548
rect 12742 4508 12808 4536
rect 12802 4496 12808 4508
rect 12860 4496 12866 4548
rect 13265 4539 13323 4545
rect 13265 4505 13277 4539
rect 13311 4536 13323 4539
rect 14829 4539 14887 4545
rect 13311 4508 14596 4536
rect 13311 4505 13323 4508
rect 13265 4499 13323 4505
rect 9048 4440 9352 4468
rect 11606 4428 11612 4480
rect 11664 4468 11670 4480
rect 13538 4468 13544 4480
rect 11664 4440 13544 4468
rect 11664 4428 11670 4440
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 14568 4468 14596 4508
rect 14829 4505 14841 4539
rect 14875 4536 14887 4539
rect 15102 4536 15108 4548
rect 14875 4508 15108 4536
rect 14875 4505 14887 4508
rect 14829 4499 14887 4505
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 15838 4496 15844 4548
rect 15896 4496 15902 4548
rect 17034 4536 17040 4548
rect 16132 4508 17040 4536
rect 16132 4468 16160 4508
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 17129 4539 17187 4545
rect 17129 4505 17141 4539
rect 17175 4536 17187 4539
rect 17402 4536 17408 4548
rect 17175 4508 17408 4536
rect 17175 4505 17187 4508
rect 17129 4499 17187 4505
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 18877 4539 18935 4545
rect 18877 4505 18889 4539
rect 18923 4505 18935 4539
rect 20162 4536 20168 4548
rect 20123 4508 20168 4536
rect 18877 4499 18935 4505
rect 14568 4440 16160 4468
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 18892 4468 18920 4499
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 20732 4536 20760 4644
rect 21177 4641 21189 4675
rect 21223 4672 21235 4675
rect 22204 4672 22232 4712
rect 24578 4700 24584 4712
rect 24636 4700 24642 4752
rect 23750 4672 23756 4684
rect 21223 4644 22232 4672
rect 22296 4644 23756 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 22296 4590 22324 4644
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 24302 4632 24308 4684
rect 24360 4672 24366 4684
rect 25317 4675 25375 4681
rect 25317 4672 25329 4675
rect 24360 4644 25329 4672
rect 24360 4632 24366 4644
rect 25317 4641 25329 4644
rect 25363 4641 25375 4675
rect 25317 4635 25375 4641
rect 25406 4632 25412 4684
rect 25464 4672 25470 4684
rect 25464 4644 27384 4672
rect 25464 4632 25470 4644
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 23256 4576 23397 4604
rect 23256 4564 23262 4576
rect 23385 4573 23397 4576
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 24762 4604 24768 4616
rect 24627 4576 24768 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4573 26019 4607
rect 27356 4590 27384 4644
rect 27614 4632 27620 4684
rect 27672 4672 27678 4684
rect 27985 4675 28043 4681
rect 27985 4672 27997 4675
rect 27672 4644 27997 4672
rect 27672 4632 27678 4644
rect 27985 4641 27997 4644
rect 28031 4641 28043 4675
rect 29012 4672 29040 4780
rect 29104 4780 33784 4808
rect 29104 4749 29132 4780
rect 33778 4768 33784 4780
rect 33836 4768 33842 4820
rect 29089 4743 29147 4749
rect 29089 4709 29101 4743
rect 29135 4709 29147 4743
rect 29089 4703 29147 4709
rect 29012 4644 29224 4672
rect 27985 4635 28043 4641
rect 25961 4567 26019 4573
rect 21266 4536 21272 4548
rect 20732 4508 21272 4536
rect 21266 4496 21272 4508
rect 21324 4496 21330 4548
rect 22925 4539 22983 4545
rect 22925 4505 22937 4539
rect 22971 4536 22983 4539
rect 24486 4536 24492 4548
rect 22971 4508 24492 4536
rect 22971 4505 22983 4508
rect 22925 4499 22983 4505
rect 24486 4496 24492 4508
rect 24544 4496 24550 4548
rect 21450 4468 21456 4480
rect 16632 4440 21456 4468
rect 16632 4428 16638 4440
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 21542 4428 21548 4480
rect 21600 4468 21606 4480
rect 23569 4471 23627 4477
rect 23569 4468 23581 4471
rect 21600 4440 23581 4468
rect 21600 4428 21606 4440
rect 23569 4437 23581 4440
rect 23615 4437 23627 4471
rect 23569 4431 23627 4437
rect 24210 4428 24216 4480
rect 24268 4468 24274 4480
rect 25682 4468 25688 4480
rect 24268 4440 25688 4468
rect 24268 4428 24274 4440
rect 25682 4428 25688 4440
rect 25740 4428 25746 4480
rect 25774 4428 25780 4480
rect 25832 4468 25838 4480
rect 25976 4468 26004 4567
rect 26237 4539 26295 4545
rect 26237 4505 26249 4539
rect 26283 4536 26295 4539
rect 26510 4536 26516 4548
rect 26283 4508 26516 4536
rect 26283 4505 26295 4508
rect 26237 4499 26295 4505
rect 26510 4496 26516 4508
rect 26568 4496 26574 4548
rect 28074 4496 28080 4548
rect 28132 4536 28138 4548
rect 28537 4539 28595 4545
rect 28537 4536 28549 4539
rect 28132 4508 28549 4536
rect 28132 4496 28138 4508
rect 28537 4505 28549 4508
rect 28583 4505 28595 4539
rect 28537 4499 28595 4505
rect 28629 4539 28687 4545
rect 28629 4505 28641 4539
rect 28675 4505 28687 4539
rect 29196 4536 29224 4644
rect 29638 4632 29644 4684
rect 29696 4672 29702 4684
rect 29733 4675 29791 4681
rect 29733 4672 29745 4675
rect 29696 4644 29745 4672
rect 29696 4632 29702 4644
rect 29733 4641 29745 4644
rect 29779 4672 29791 4675
rect 31941 4675 31999 4681
rect 31941 4672 31953 4675
rect 29779 4644 31953 4672
rect 29779 4641 29791 4644
rect 29733 4635 29791 4641
rect 31941 4641 31953 4644
rect 31987 4672 31999 4675
rect 32306 4672 32312 4684
rect 31987 4644 32312 4672
rect 31987 4641 31999 4644
rect 31941 4635 31999 4641
rect 32306 4632 32312 4644
rect 32364 4632 32370 4684
rect 32858 4632 32864 4684
rect 32916 4672 32922 4684
rect 32916 4644 34192 4672
rect 32916 4632 32922 4644
rect 33686 4604 33692 4616
rect 33350 4576 33692 4604
rect 33686 4564 33692 4576
rect 33744 4564 33750 4616
rect 34164 4613 34192 4644
rect 34330 4632 34336 4684
rect 34388 4672 34394 4684
rect 35161 4675 35219 4681
rect 35161 4672 35173 4675
rect 34388 4644 35173 4672
rect 34388 4632 34394 4644
rect 35161 4641 35173 4644
rect 35207 4641 35219 4675
rect 35161 4635 35219 4641
rect 37461 4675 37519 4681
rect 37461 4641 37473 4675
rect 37507 4672 37519 4675
rect 39298 4672 39304 4684
rect 37507 4644 39304 4672
rect 37507 4641 37519 4644
rect 37461 4635 37519 4641
rect 39298 4632 39304 4644
rect 39356 4632 39362 4684
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4573 34207 4607
rect 34149 4567 34207 4573
rect 34238 4564 34244 4616
rect 34296 4604 34302 4616
rect 34885 4607 34943 4613
rect 34296 4576 34341 4604
rect 34296 4564 34302 4576
rect 34885 4573 34897 4607
rect 34931 4573 34943 4607
rect 36722 4604 36728 4616
rect 36683 4576 36728 4604
rect 34885 4567 34943 4573
rect 30009 4539 30067 4545
rect 30009 4536 30021 4539
rect 29196 4508 30021 4536
rect 28629 4499 28687 4505
rect 30009 4505 30021 4508
rect 30055 4505 30067 4539
rect 30009 4499 30067 4505
rect 27154 4468 27160 4480
rect 25832 4440 27160 4468
rect 25832 4428 25838 4440
rect 27154 4428 27160 4440
rect 27212 4428 27218 4480
rect 28644 4468 28672 4499
rect 31018 4496 31024 4548
rect 31076 4496 31082 4548
rect 31846 4536 31852 4548
rect 31312 4508 31852 4536
rect 31312 4468 31340 4508
rect 31846 4496 31852 4508
rect 31904 4496 31910 4548
rect 32217 4539 32275 4545
rect 32217 4505 32229 4539
rect 32263 4536 32275 4539
rect 32490 4536 32496 4548
rect 32263 4508 32496 4536
rect 32263 4505 32275 4508
rect 32217 4499 32275 4505
rect 28644 4440 31340 4468
rect 31481 4471 31539 4477
rect 31481 4437 31493 4471
rect 31527 4468 31539 4471
rect 32232 4468 32260 4499
rect 32490 4496 32496 4508
rect 32548 4496 32554 4548
rect 33520 4508 33824 4536
rect 31527 4440 32260 4468
rect 31527 4437 31539 4440
rect 31481 4431 31539 4437
rect 32582 4428 32588 4480
rect 32640 4468 32646 4480
rect 33520 4468 33548 4508
rect 32640 4440 33548 4468
rect 32640 4428 32646 4440
rect 33594 4428 33600 4480
rect 33652 4468 33658 4480
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 33652 4440 33701 4468
rect 33652 4428 33658 4440
rect 33689 4437 33701 4440
rect 33735 4437 33747 4471
rect 33796 4468 33824 4508
rect 33870 4496 33876 4548
rect 33928 4536 33934 4548
rect 34900 4536 34928 4567
rect 36722 4564 36728 4576
rect 36780 4564 36786 4616
rect 37737 4607 37795 4613
rect 37737 4573 37749 4607
rect 37783 4604 37795 4607
rect 38838 4604 38844 4616
rect 37783 4576 38844 4604
rect 37783 4573 37795 4576
rect 37737 4567 37795 4573
rect 38838 4564 38844 4576
rect 38896 4564 38902 4616
rect 38654 4536 38660 4548
rect 33928 4508 34928 4536
rect 34992 4508 38660 4536
rect 33928 4496 33934 4508
rect 34992 4468 35020 4508
rect 38654 4496 38660 4508
rect 38712 4496 38718 4548
rect 33796 4440 35020 4468
rect 33689 4431 33747 4437
rect 35802 4428 35808 4480
rect 35860 4468 35866 4480
rect 36909 4471 36967 4477
rect 36909 4468 36921 4471
rect 35860 4440 36921 4468
rect 35860 4428 35866 4440
rect 36909 4437 36921 4440
rect 36955 4437 36967 4471
rect 36909 4431 36967 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 3752 4236 4660 4264
rect 3752 4224 3758 4236
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 2869 4199 2927 4205
rect 2869 4196 2881 4199
rect 2832 4168 2881 4196
rect 2832 4156 2838 4168
rect 2869 4165 2881 4168
rect 2915 4165 2927 4199
rect 4522 4196 4528 4208
rect 4483 4168 4528 4196
rect 2869 4159 2927 4165
rect 4522 4156 4528 4168
rect 4580 4156 4586 4208
rect 4632 4196 4660 4236
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 8570 4264 8576 4276
rect 4856 4236 8576 4264
rect 4856 4224 4862 4236
rect 8570 4224 8576 4236
rect 8628 4264 8634 4276
rect 14182 4264 14188 4276
rect 8628 4236 11652 4264
rect 8628 4224 8634 4236
rect 7009 4199 7067 4205
rect 7009 4196 7021 4199
rect 4632 4168 5014 4196
rect 6748 4168 7021 4196
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1452 4100 1593 4128
rect 1452 4088 1458 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6748 4128 6776 4168
rect 7009 4165 7021 4168
rect 7055 4165 7067 4199
rect 7009 4159 7067 4165
rect 7098 4156 7104 4208
rect 7156 4196 7162 4208
rect 7156 4168 7498 4196
rect 7156 4156 7162 4168
rect 8938 4128 8944 4140
rect 6052 4100 6776 4128
rect 8899 4100 8944 4128
rect 6052 4088 6058 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 11624 4128 11652 4236
rect 11716 4236 14188 4264
rect 11716 4205 11744 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 16298 4224 16304 4276
rect 16356 4264 16362 4276
rect 16356 4236 20944 4264
rect 16356 4224 16362 4236
rect 11701 4199 11759 4205
rect 11701 4165 11713 4199
rect 11747 4165 11759 4199
rect 13446 4196 13452 4208
rect 11701 4159 11759 4165
rect 11808 4168 13452 4196
rect 11808 4128 11836 4168
rect 13446 4156 13452 4168
rect 13504 4156 13510 4208
rect 14918 4196 14924 4208
rect 14582 4168 14924 4196
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 15102 4196 15108 4208
rect 15063 4168 15108 4196
rect 15102 4156 15108 4168
rect 15160 4156 15166 4208
rect 16117 4199 16175 4205
rect 16117 4165 16129 4199
rect 16163 4196 16175 4199
rect 17405 4199 17463 4205
rect 16163 4168 17356 4196
rect 16163 4165 16175 4168
rect 16117 4159 16175 4165
rect 11624 4100 11836 4128
rect 17328 4128 17356 4168
rect 17405 4165 17417 4199
rect 17451 4196 17463 4199
rect 18598 4196 18604 4208
rect 17451 4168 18604 4196
rect 17451 4165 17463 4168
rect 17405 4159 17463 4165
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 18782 4156 18788 4208
rect 18840 4156 18846 4208
rect 20916 4196 20944 4236
rect 20990 4224 20996 4276
rect 21048 4264 21054 4276
rect 24210 4264 24216 4276
rect 21048 4236 24216 4264
rect 21048 4224 21054 4236
rect 24210 4224 24216 4236
rect 24268 4224 24274 4276
rect 24302 4224 24308 4276
rect 24360 4224 24366 4276
rect 24486 4224 24492 4276
rect 24544 4264 24550 4276
rect 30282 4264 30288 4276
rect 24544 4236 30288 4264
rect 24544 4224 24550 4236
rect 30282 4224 30288 4236
rect 30340 4224 30346 4276
rect 30558 4224 30564 4276
rect 30616 4264 30622 4276
rect 31570 4264 31576 4276
rect 30616 4236 31576 4264
rect 30616 4224 30622 4236
rect 31570 4224 31576 4236
rect 31628 4224 31634 4276
rect 31846 4224 31852 4276
rect 31904 4264 31910 4276
rect 32582 4264 32588 4276
rect 31904 4236 32588 4264
rect 31904 4224 31910 4236
rect 32582 4224 32588 4236
rect 32640 4224 32646 4276
rect 32674 4224 32680 4276
rect 32732 4264 32738 4276
rect 33873 4267 33931 4273
rect 33873 4264 33885 4267
rect 32732 4236 33885 4264
rect 32732 4224 32738 4236
rect 33873 4233 33885 4236
rect 33919 4264 33931 4267
rect 33919 4236 36308 4264
rect 33919 4233 33931 4236
rect 33873 4227 33931 4233
rect 21818 4196 21824 4208
rect 20916 4168 21824 4196
rect 21818 4156 21824 4168
rect 21876 4156 21882 4208
rect 22186 4196 22192 4208
rect 22147 4168 22192 4196
rect 22186 4156 22192 4168
rect 22244 4156 22250 4208
rect 24320 4196 24348 4224
rect 23860 4168 24348 4196
rect 17954 4128 17960 4140
rect 17328 4100 17960 4128
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 20806 4128 20812 4140
rect 20767 4100 20812 4128
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 23860 4137 23888 4168
rect 25130 4156 25136 4208
rect 25188 4156 25194 4208
rect 25682 4156 25688 4208
rect 25740 4196 25746 4208
rect 27522 4196 27528 4208
rect 25740 4168 27528 4196
rect 25740 4156 25746 4168
rect 27522 4156 27528 4168
rect 27580 4156 27586 4208
rect 31202 4196 31208 4208
rect 31142 4168 31208 4196
rect 31202 4156 31208 4168
rect 31260 4156 31266 4208
rect 32306 4196 32312 4208
rect 32140 4168 32312 4196
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4097 23903 4131
rect 26329 4131 26387 4137
rect 26329 4128 26341 4131
rect 23845 4091 23903 4097
rect 25332 4100 26341 4128
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2958 4060 2964 4072
rect 2823 4032 2964 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4060 3847 4063
rect 3970 4060 3976 4072
rect 3835 4032 3976 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4212 4032 4261 4060
rect 4212 4020 4218 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 9125 4063 9183 4069
rect 6788 4032 6833 4060
rect 6788 4020 6794 4032
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 10778 4060 10784 4072
rect 10739 4032 10784 4060
rect 9125 4023 9183 4029
rect 658 3952 664 4004
rect 716 3992 722 4004
rect 3234 3992 3240 4004
rect 716 3964 3240 3992
rect 716 3952 722 3964
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 5994 3992 6000 4004
rect 5955 3964 6000 3992
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 9140 3992 9168 4023
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 11112 4032 12449 4060
rect 11112 4020 11118 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13354 4060 13360 4072
rect 13315 4032 13360 4060
rect 13081 4023 13139 4029
rect 8260 3964 9168 3992
rect 8260 3952 8266 3964
rect 1762 3924 1768 3936
rect 1723 3896 1768 3924
rect 1762 3884 1768 3896
rect 1820 3884 1826 3936
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 7558 3924 7564 3936
rect 2832 3896 7564 3924
rect 2832 3884 2838 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 8478 3924 8484 3936
rect 8439 3896 8484 3924
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 12986 3924 12992 3936
rect 8812 3896 12992 3924
rect 8812 3884 8818 3896
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13096 3924 13124 4023
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 16298 4060 16304 4072
rect 16259 4032 16304 4060
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18322 4060 18328 4072
rect 18283 4032 18328 4060
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 18472 4032 20085 4060
rect 18472 4020 18478 4032
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 20533 4063 20591 4069
rect 20533 4029 20545 4063
rect 20579 4029 20591 4063
rect 20533 4023 20591 4029
rect 20548 3992 20576 4023
rect 21818 4020 21824 4072
rect 21876 4060 21882 4072
rect 22097 4063 22155 4069
rect 22097 4060 22109 4063
rect 21876 4032 22109 4060
rect 21876 4020 21882 4032
rect 22097 4029 22109 4032
rect 22143 4029 22155 4063
rect 22097 4023 22155 4029
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 23109 4063 23167 4069
rect 23109 4060 23121 4063
rect 22428 4032 23121 4060
rect 22428 4020 22434 4032
rect 23109 4029 23121 4032
rect 23155 4060 23167 4063
rect 23474 4060 23480 4072
rect 23155 4032 23480 4060
rect 23155 4029 23167 4032
rect 23109 4023 23167 4029
rect 23474 4020 23480 4032
rect 23532 4020 23538 4072
rect 19352 3964 20576 3992
rect 14090 3924 14096 3936
rect 13096 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 17494 3924 17500 3936
rect 17455 3896 17500 3924
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 19352 3924 19380 3964
rect 20898 3952 20904 4004
rect 20956 3992 20962 4004
rect 23860 3992 23888 4091
rect 24121 4063 24179 4069
rect 24121 4029 24133 4063
rect 24167 4060 24179 4063
rect 24210 4060 24216 4072
rect 24167 4032 24216 4060
rect 24167 4029 24179 4032
rect 24121 4023 24179 4029
rect 24210 4020 24216 4032
rect 24268 4020 24274 4072
rect 24854 4020 24860 4072
rect 24912 4060 24918 4072
rect 25332 4060 25360 4100
rect 26329 4097 26341 4100
rect 26375 4097 26387 4131
rect 26329 4091 26387 4097
rect 28534 4088 28540 4140
rect 28592 4088 28598 4140
rect 29638 4128 29644 4140
rect 29599 4100 29644 4128
rect 29638 4088 29644 4100
rect 29696 4088 29702 4140
rect 32140 4137 32168 4168
rect 32306 4156 32312 4168
rect 32364 4156 32370 4208
rect 33410 4156 33416 4208
rect 33468 4156 33474 4208
rect 34609 4199 34667 4205
rect 34609 4196 34621 4199
rect 34440 4168 34621 4196
rect 32125 4131 32183 4137
rect 32125 4097 32137 4131
rect 32171 4097 32183 4131
rect 34146 4128 34152 4140
rect 34107 4100 34152 4128
rect 32125 4091 32183 4097
rect 34146 4088 34152 4100
rect 34204 4128 34210 4140
rect 34440 4128 34468 4168
rect 34609 4165 34621 4168
rect 34655 4165 34667 4199
rect 34609 4159 34667 4165
rect 34701 4199 34759 4205
rect 34701 4165 34713 4199
rect 34747 4196 34759 4199
rect 34747 4168 35480 4196
rect 34747 4165 34759 4168
rect 34701 4159 34759 4165
rect 34204 4100 34468 4128
rect 35452 4128 35480 4168
rect 35894 4128 35900 4140
rect 35452 4100 35900 4128
rect 34204 4088 34210 4100
rect 35894 4088 35900 4100
rect 35952 4088 35958 4140
rect 35986 4088 35992 4140
rect 36044 4128 36050 4140
rect 36173 4131 36231 4137
rect 36173 4128 36185 4131
rect 36044 4100 36185 4128
rect 36044 4088 36050 4100
rect 36173 4097 36185 4100
rect 36219 4097 36231 4131
rect 36280 4128 36308 4236
rect 37090 4128 37096 4140
rect 36280 4100 37096 4128
rect 36173 4091 36231 4097
rect 37090 4088 37096 4100
rect 37148 4088 37154 4140
rect 37550 4088 37556 4140
rect 37608 4128 37614 4140
rect 37737 4131 37795 4137
rect 37737 4128 37749 4131
rect 37608 4100 37749 4128
rect 37608 4088 37614 4100
rect 37737 4097 37749 4100
rect 37783 4097 37795 4131
rect 37737 4091 37795 4097
rect 24912 4032 25360 4060
rect 24912 4020 24918 4032
rect 25590 4020 25596 4072
rect 25648 4060 25654 4072
rect 25869 4063 25927 4069
rect 25869 4060 25881 4063
rect 25648 4032 25881 4060
rect 25648 4020 25654 4032
rect 25869 4029 25881 4032
rect 25915 4029 25927 4063
rect 27154 4060 27160 4072
rect 27115 4032 27160 4060
rect 25869 4023 25927 4029
rect 27154 4020 27160 4032
rect 27212 4020 27218 4072
rect 27264 4032 29132 4060
rect 20956 3964 23888 3992
rect 20956 3952 20962 3964
rect 25498 3952 25504 4004
rect 25556 3992 25562 4004
rect 26234 3992 26240 4004
rect 25556 3964 26240 3992
rect 25556 3952 25562 3964
rect 26234 3952 26240 3964
rect 26292 3952 26298 4004
rect 26421 3995 26479 4001
rect 26421 3961 26433 3995
rect 26467 3992 26479 3995
rect 27264 3992 27292 4032
rect 26467 3964 27292 3992
rect 26467 3961 26479 3964
rect 26421 3955 26479 3961
rect 17736 3896 19380 3924
rect 17736 3884 17742 3896
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 23014 3924 23020 3936
rect 20312 3896 23020 3924
rect 20312 3884 20318 3896
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23106 3884 23112 3936
rect 23164 3924 23170 3936
rect 27246 3924 27252 3936
rect 23164 3896 27252 3924
rect 23164 3884 23170 3896
rect 27246 3884 27252 3896
rect 27304 3884 27310 3936
rect 27420 3927 27478 3933
rect 27420 3893 27432 3927
rect 27466 3924 27478 3927
rect 27614 3924 27620 3936
rect 27466 3896 27620 3924
rect 27466 3893 27478 3896
rect 27420 3887 27478 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 29104 3924 29132 4032
rect 29178 4020 29184 4072
rect 29236 4060 29242 4072
rect 29236 4032 29281 4060
rect 29236 4020 29242 4032
rect 29454 4020 29460 4072
rect 29512 4060 29518 4072
rect 29914 4060 29920 4072
rect 29512 4032 29920 4060
rect 29512 4020 29518 4032
rect 29914 4020 29920 4032
rect 29972 4020 29978 4072
rect 30466 4020 30472 4072
rect 30524 4060 30530 4072
rect 31389 4063 31447 4069
rect 30524 4032 31340 4060
rect 30524 4020 30530 4032
rect 31312 3992 31340 4032
rect 31389 4029 31401 4063
rect 31435 4060 31447 4063
rect 32401 4063 32459 4069
rect 32401 4060 32413 4063
rect 31435 4032 32413 4060
rect 31435 4029 31447 4032
rect 31389 4023 31447 4029
rect 32401 4029 32413 4032
rect 32447 4060 32459 4063
rect 34422 4060 34428 4072
rect 32447 4032 34428 4060
rect 32447 4029 32459 4032
rect 32401 4023 32459 4029
rect 34422 4020 34428 4032
rect 34480 4020 34486 4072
rect 34698 4020 34704 4072
rect 34756 4060 34762 4072
rect 35434 4060 35440 4072
rect 34756 4032 35440 4060
rect 34756 4020 34762 4032
rect 35434 4020 35440 4032
rect 35492 4020 35498 4072
rect 35618 4060 35624 4072
rect 35579 4032 35624 4060
rect 35618 4020 35624 4032
rect 35676 4020 35682 4072
rect 37461 4063 37519 4069
rect 37461 4029 37473 4063
rect 37507 4060 37519 4063
rect 38654 4060 38660 4072
rect 37507 4032 38660 4060
rect 37507 4029 37519 4032
rect 37461 4023 37519 4029
rect 38654 4020 38660 4032
rect 38712 4020 38718 4072
rect 35342 3992 35348 4004
rect 31312 3964 31754 3992
rect 31294 3924 31300 3936
rect 29104 3896 31300 3924
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 31726 3924 31754 3964
rect 33428 3964 35348 3992
rect 33428 3924 33456 3964
rect 35342 3952 35348 3964
rect 35400 3952 35406 4004
rect 36262 3992 36268 4004
rect 36004 3964 36268 3992
rect 31726 3896 33456 3924
rect 33502 3884 33508 3936
rect 33560 3924 33566 3936
rect 33778 3924 33784 3936
rect 33560 3896 33784 3924
rect 33560 3884 33566 3896
rect 33778 3884 33784 3896
rect 33836 3884 33842 3936
rect 33962 3884 33968 3936
rect 34020 3924 34026 3936
rect 36004 3924 36032 3964
rect 36262 3952 36268 3964
rect 36320 3952 36326 4004
rect 34020 3896 36032 3924
rect 34020 3884 34026 3896
rect 36078 3884 36084 3936
rect 36136 3924 36142 3936
rect 36357 3927 36415 3933
rect 36357 3924 36369 3927
rect 36136 3896 36369 3924
rect 36136 3884 36142 3896
rect 36357 3893 36369 3896
rect 36403 3893 36415 3927
rect 36357 3887 36415 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 4706 3720 4712 3732
rect 3436 3692 4712 3720
rect 3326 3652 3332 3664
rect 3287 3624 3332 3652
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 2832 3556 2877 3584
rect 2832 3544 2838 3556
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 2869 3451 2927 3457
rect 2096 3420 2774 3448
rect 2096 3408 2102 3420
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3380 2191 3383
rect 2590 3380 2596 3392
rect 2179 3352 2596 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 2746 3380 2774 3420
rect 2869 3417 2881 3451
rect 2915 3448 2927 3451
rect 3436 3448 3464 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 5960 3692 6377 3720
rect 5960 3680 5966 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 18782 3720 18788 3732
rect 7616 3692 18788 3720
rect 7616 3680 7622 3692
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 28074 3720 28080 3732
rect 19484 3692 28080 3720
rect 19484 3680 19490 3692
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 10870 3652 10876 3664
rect 8168 3624 10876 3652
rect 8168 3612 8174 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 16574 3612 16580 3664
rect 16632 3652 16638 3664
rect 16632 3624 16988 3652
rect 16632 3612 16638 3624
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4304 3556 4629 3584
rect 4304 3544 4310 3556
rect 4617 3553 4629 3556
rect 4663 3584 4675 3587
rect 7101 3587 7159 3593
rect 4663 3556 6408 3584
rect 4663 3553 4675 3556
rect 4617 3547 4675 3553
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 6380 3516 6408 3556
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7190 3584 7196 3596
rect 7147 3556 7196 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7190 3544 7196 3556
rect 7248 3584 7254 3596
rect 8754 3584 8760 3596
rect 7248 3556 8760 3584
rect 7248 3544 7254 3556
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9214 3584 9220 3596
rect 9175 3556 9220 3584
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 10042 3584 10048 3596
rect 10003 3556 10048 3584
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 10152 3556 13093 3584
rect 6730 3516 6736 3528
rect 6380 3488 6736 3516
rect 6730 3476 6736 3488
rect 6788 3516 6794 3528
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 6788 3488 6837 3516
rect 6788 3476 6794 3488
rect 6825 3485 6837 3488
rect 6871 3485 6883 3519
rect 6825 3479 6883 3485
rect 2915 3420 3464 3448
rect 3528 3420 4844 3448
rect 2915 3417 2927 3420
rect 2869 3411 2927 3417
rect 3528 3380 3556 3420
rect 4062 3380 4068 3392
rect 2746 3352 3556 3380
rect 4023 3352 4068 3380
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4816 3380 4844 3420
rect 4890 3408 4896 3460
rect 4948 3448 4954 3460
rect 6270 3448 6276 3460
rect 4948 3420 4993 3448
rect 6118 3420 6276 3448
rect 4948 3408 4954 3420
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 7558 3408 7564 3460
rect 7616 3408 7622 3460
rect 8404 3420 8708 3448
rect 8404 3380 8432 3420
rect 8570 3380 8576 3392
rect 4816 3352 8432 3380
rect 8531 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 8680 3380 8708 3420
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 9364 3420 9409 3448
rect 9364 3408 9370 3420
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 10152 3448 10180 3556
rect 13081 3553 13093 3556
rect 13127 3553 13139 3587
rect 14274 3584 14280 3596
rect 14187 3556 14280 3584
rect 13081 3547 13139 3553
rect 14274 3544 14280 3556
rect 14332 3584 14338 3596
rect 16960 3584 16988 3624
rect 18322 3612 18328 3664
rect 18380 3652 18386 3664
rect 18690 3652 18696 3664
rect 18380 3624 18696 3652
rect 18380 3612 18386 3624
rect 18690 3612 18696 3624
rect 18748 3612 18754 3664
rect 22462 3612 22468 3664
rect 22520 3612 22526 3664
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 14332 3556 16804 3584
rect 16960 3556 17141 3584
rect 14332 3544 14338 3556
rect 16776 3528 16804 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 20254 3584 20260 3596
rect 20215 3556 20260 3584
rect 17129 3547 17187 3553
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 21726 3544 21732 3596
rect 21784 3584 21790 3596
rect 22005 3587 22063 3593
rect 22005 3584 22017 3587
rect 21784 3556 22017 3584
rect 21784 3544 21790 3556
rect 22005 3553 22017 3556
rect 22051 3553 22063 3587
rect 22480 3584 22508 3612
rect 22940 3593 22968 3692
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 38194 3720 38200 3732
rect 38155 3692 38200 3720
rect 38194 3680 38200 3692
rect 38252 3680 38258 3732
rect 23014 3612 23020 3664
rect 23072 3652 23078 3664
rect 23072 3624 24624 3652
rect 23072 3612 23078 3624
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 22480 3556 22569 3584
rect 22005 3547 22063 3553
rect 22557 3553 22569 3556
rect 22603 3553 22615 3587
rect 22557 3547 22615 3553
rect 22925 3587 22983 3593
rect 22925 3553 22937 3587
rect 22971 3553 22983 3587
rect 24596 3584 24624 3624
rect 24762 3612 24768 3664
rect 24820 3652 24826 3664
rect 24820 3624 25912 3652
rect 24820 3612 24826 3624
rect 25590 3584 25596 3596
rect 24596 3556 25596 3584
rect 22925 3547 22983 3553
rect 25590 3544 25596 3556
rect 25648 3544 25654 3596
rect 25774 3584 25780 3596
rect 25735 3556 25780 3584
rect 25774 3544 25780 3556
rect 25832 3544 25838 3596
rect 25884 3584 25912 3624
rect 27246 3612 27252 3664
rect 27304 3652 27310 3664
rect 30558 3652 30564 3664
rect 27304 3624 30564 3652
rect 27304 3612 27310 3624
rect 30558 3612 30564 3624
rect 30616 3612 30622 3664
rect 30668 3624 36584 3652
rect 30668 3584 30696 3624
rect 25884 3556 28304 3584
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13722 3516 13728 3528
rect 13587 3488 13728 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16816 3488 16865 3516
rect 16816 3476 16822 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 18230 3476 18236 3528
rect 18288 3476 18294 3528
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19981 3519 20039 3525
rect 19981 3516 19993 3519
rect 19300 3488 19993 3516
rect 19300 3476 19306 3488
rect 19981 3485 19993 3488
rect 20027 3485 20039 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 19981 3479 20039 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3516 27859 3519
rect 27890 3516 27896 3528
rect 27847 3488 27896 3516
rect 27847 3485 27859 3488
rect 27801 3479 27859 3485
rect 27890 3476 27896 3488
rect 27948 3476 27954 3528
rect 28276 3525 28304 3556
rect 28368 3556 30696 3584
rect 28261 3519 28319 3525
rect 28261 3485 28273 3519
rect 28307 3485 28319 3519
rect 28261 3479 28319 3485
rect 11330 3448 11336 3460
rect 9640 3420 10180 3448
rect 11291 3420 11336 3448
rect 9640 3408 9646 3420
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 14553 3451 14611 3457
rect 11440 3420 11822 3448
rect 11440 3380 11468 3420
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 14642 3448 14648 3460
rect 14599 3420 14648 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 15194 3408 15200 3460
rect 15252 3408 15258 3460
rect 16298 3448 16304 3460
rect 16211 3420 16304 3448
rect 16298 3408 16304 3420
rect 16356 3448 16362 3460
rect 17218 3448 17224 3460
rect 16356 3420 17224 3448
rect 16356 3408 16362 3420
rect 17218 3408 17224 3420
rect 17276 3408 17282 3460
rect 18877 3451 18935 3457
rect 18877 3417 18889 3451
rect 18923 3448 18935 3451
rect 18966 3448 18972 3460
rect 18923 3420 18972 3448
rect 18923 3417 18935 3420
rect 18877 3411 18935 3417
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 19058 3408 19064 3460
rect 19116 3448 19122 3460
rect 20530 3448 20536 3460
rect 19116 3420 20536 3448
rect 19116 3408 19122 3420
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 20714 3408 20720 3460
rect 20772 3408 20778 3460
rect 22646 3408 22652 3460
rect 22704 3448 22710 3460
rect 22704 3420 22749 3448
rect 22704 3408 22710 3420
rect 23934 3408 23940 3460
rect 23992 3448 23998 3460
rect 26053 3451 26111 3457
rect 23992 3420 24900 3448
rect 23992 3408 23998 3420
rect 8680 3352 11468 3380
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 14090 3380 14096 3392
rect 13679 3352 14096 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 21818 3380 21824 3392
rect 18840 3352 21824 3380
rect 18840 3340 18846 3352
rect 21818 3340 21824 3352
rect 21876 3380 21882 3392
rect 23106 3380 23112 3392
rect 21876 3352 23112 3380
rect 21876 3340 21882 3352
rect 23106 3340 23112 3352
rect 23164 3340 23170 3392
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 24765 3383 24823 3389
rect 24765 3380 24777 3383
rect 23256 3352 24777 3380
rect 23256 3340 23262 3352
rect 24765 3349 24777 3352
rect 24811 3349 24823 3383
rect 24872 3380 24900 3420
rect 26053 3417 26065 3451
rect 26099 3448 26111 3451
rect 26142 3448 26148 3460
rect 26099 3420 26148 3448
rect 26099 3417 26111 3420
rect 26053 3411 26111 3417
rect 26142 3408 26148 3420
rect 26200 3408 26206 3460
rect 27278 3420 27936 3448
rect 27706 3380 27712 3392
rect 24872 3352 27712 3380
rect 24765 3343 24823 3349
rect 27706 3340 27712 3352
rect 27764 3340 27770 3392
rect 27908 3380 27936 3420
rect 27982 3408 27988 3460
rect 28040 3448 28046 3460
rect 28368 3448 28396 3556
rect 30742 3544 30748 3596
rect 30800 3584 30806 3596
rect 30800 3556 30845 3584
rect 30800 3544 30806 3556
rect 30926 3544 30932 3596
rect 30984 3584 30990 3596
rect 32582 3584 32588 3596
rect 30984 3556 31029 3584
rect 32543 3556 32588 3584
rect 30984 3544 30990 3556
rect 32582 3544 32588 3556
rect 32640 3544 32646 3596
rect 33137 3587 33195 3593
rect 33137 3553 33149 3587
rect 33183 3584 33195 3587
rect 34330 3584 34336 3596
rect 33183 3556 34336 3584
rect 33183 3553 33195 3556
rect 33137 3547 33195 3553
rect 34330 3544 34336 3556
rect 34388 3544 34394 3596
rect 35250 3584 35256 3596
rect 35211 3556 35256 3584
rect 35250 3544 35256 3556
rect 35308 3544 35314 3596
rect 36556 3593 36584 3624
rect 36541 3587 36599 3593
rect 36541 3553 36553 3587
rect 36587 3553 36599 3587
rect 36541 3547 36599 3553
rect 37553 3587 37611 3593
rect 37553 3553 37565 3587
rect 37599 3584 37611 3587
rect 38470 3584 38476 3596
rect 37599 3556 38476 3584
rect 37599 3553 37611 3556
rect 37553 3547 37611 3553
rect 38470 3544 38476 3556
rect 38528 3544 38534 3596
rect 29730 3476 29736 3528
rect 29788 3516 29794 3528
rect 30009 3519 30067 3525
rect 30009 3516 30021 3519
rect 29788 3488 30021 3516
rect 29788 3476 29794 3488
rect 30009 3485 30021 3488
rect 30055 3485 30067 3519
rect 30009 3479 30067 3485
rect 32508 3488 32720 3516
rect 28040 3420 28396 3448
rect 29089 3451 29147 3457
rect 28040 3408 28046 3420
rect 29089 3417 29101 3451
rect 29135 3448 29147 3451
rect 29638 3448 29644 3460
rect 29135 3420 29644 3448
rect 29135 3417 29147 3420
rect 29089 3411 29147 3417
rect 29638 3408 29644 3420
rect 29696 3408 29702 3460
rect 32508 3448 32536 3488
rect 29748 3420 32536 3448
rect 32692 3448 32720 3488
rect 37918 3476 37924 3528
rect 37976 3516 37982 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 37976 3488 38117 3516
rect 37976 3476 37982 3488
rect 38105 3485 38117 3488
rect 38151 3485 38163 3519
rect 38105 3479 38163 3485
rect 33134 3448 33140 3460
rect 32692 3420 33140 3448
rect 29748 3380 29776 3420
rect 33134 3408 33140 3420
rect 33192 3408 33198 3460
rect 33229 3451 33287 3457
rect 33229 3417 33241 3451
rect 33275 3448 33287 3451
rect 33962 3448 33968 3460
rect 33275 3420 33968 3448
rect 33275 3417 33287 3420
rect 33229 3411 33287 3417
rect 33962 3408 33968 3420
rect 34020 3408 34026 3460
rect 34054 3408 34060 3460
rect 34112 3448 34118 3460
rect 34149 3451 34207 3457
rect 34149 3448 34161 3451
rect 34112 3420 34161 3448
rect 34112 3408 34118 3420
rect 34149 3417 34161 3420
rect 34195 3417 34207 3451
rect 34149 3411 34207 3417
rect 34977 3451 35035 3457
rect 34977 3417 34989 3451
rect 35023 3417 35035 3451
rect 34977 3411 35035 3417
rect 35069 3451 35127 3457
rect 35069 3417 35081 3451
rect 35115 3448 35127 3451
rect 35342 3448 35348 3460
rect 35115 3420 35348 3448
rect 35115 3417 35127 3420
rect 35069 3411 35127 3417
rect 27908 3352 29776 3380
rect 30193 3383 30251 3389
rect 30193 3349 30205 3383
rect 30239 3380 30251 3383
rect 30282 3380 30288 3392
rect 30239 3352 30288 3380
rect 30239 3349 30251 3352
rect 30193 3343 30251 3349
rect 30282 3340 30288 3352
rect 30340 3340 30346 3392
rect 30742 3340 30748 3392
rect 30800 3380 30806 3392
rect 34992 3380 35020 3411
rect 35342 3408 35348 3420
rect 35400 3408 35406 3460
rect 36630 3448 36636 3460
rect 36591 3420 36636 3448
rect 36630 3408 36636 3420
rect 36688 3408 36694 3460
rect 30800 3352 35020 3380
rect 30800 3340 30806 3352
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 5166 3176 5172 3188
rect 3436 3148 5172 3176
rect 2133 3111 2191 3117
rect 2133 3077 2145 3111
rect 2179 3108 2191 3111
rect 3234 3108 3240 3120
rect 2179 3080 3240 3108
rect 2179 3077 2191 3080
rect 2133 3071 2191 3077
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 3436 3040 3464 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 9306 3176 9312 3188
rect 6512 3148 9312 3176
rect 6512 3136 6518 3148
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 12894 3176 12900 3188
rect 9456 3148 12900 3176
rect 9456 3136 9462 3148
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 16298 3176 16304 3188
rect 13044 3148 16304 3176
rect 13044 3136 13050 3148
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 17770 3176 17776 3188
rect 16408 3148 17776 3176
rect 4525 3111 4583 3117
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 4798 3108 4804 3120
rect 4571 3080 4804 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 5534 3068 5540 3120
rect 5592 3068 5598 3120
rect 7364 3111 7422 3117
rect 7364 3077 7376 3111
rect 7410 3108 7422 3111
rect 7466 3108 7472 3120
rect 7410 3080 7472 3108
rect 7410 3077 7422 3080
rect 7364 3071 7422 3077
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 7834 3068 7840 3120
rect 7892 3068 7898 3120
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 8904 3080 10074 3108
rect 8904 3068 8910 3080
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 10928 3080 12558 3108
rect 10928 3068 10934 3080
rect 14826 3068 14832 3120
rect 14884 3108 14890 3120
rect 14884 3080 15042 3108
rect 14884 3068 14890 3080
rect 2823 3012 3464 3040
rect 3513 3043 3571 3049
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 4246 3040 4252 3052
rect 4207 3012 4252 3040
rect 3513 3003 3571 3009
rect 1026 2864 1032 2916
rect 1084 2904 1090 2916
rect 3528 2904 3556 3003
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 11112 3012 11805 3040
rect 11112 3000 11118 3012
rect 11793 3009 11805 3012
rect 11839 3009 11851 3043
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 11793 3003 11851 3009
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 16408 3040 16436 3148
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 19242 3176 19248 3188
rect 18104 3148 19248 3176
rect 18104 3136 18110 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 21818 3176 21824 3188
rect 19536 3148 21824 3176
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 17092 3080 17618 3108
rect 17092 3068 17098 3080
rect 19260 3049 19288 3136
rect 19536 3117 19564 3148
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 21910 3136 21916 3188
rect 21968 3176 21974 3188
rect 22554 3176 22560 3188
rect 21968 3148 22560 3176
rect 21968 3136 21974 3148
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 26513 3179 26571 3185
rect 26513 3176 26525 3179
rect 22664 3148 26525 3176
rect 19521 3111 19579 3117
rect 19521 3077 19533 3111
rect 19567 3077 19579 3111
rect 19521 3071 19579 3077
rect 20070 3068 20076 3120
rect 20128 3068 20134 3120
rect 21266 3108 21272 3120
rect 21227 3080 21272 3108
rect 21266 3068 21272 3080
rect 21324 3068 21330 3120
rect 22186 3068 22192 3120
rect 22244 3108 22250 3120
rect 22664 3108 22692 3148
rect 26513 3145 26525 3148
rect 26559 3145 26571 3179
rect 26513 3139 26571 3145
rect 27448 3148 31248 3176
rect 22244 3080 22692 3108
rect 22244 3068 22250 3080
rect 22922 3068 22928 3120
rect 22980 3068 22986 3120
rect 24486 3108 24492 3120
rect 24447 3080 24492 3108
rect 24486 3068 24492 3080
rect 24544 3068 24550 3120
rect 24946 3068 24952 3120
rect 25004 3068 25010 3120
rect 26326 3068 26332 3120
rect 26384 3108 26390 3120
rect 27062 3108 27068 3120
rect 26384 3080 27068 3108
rect 26384 3068 26390 3080
rect 27062 3068 27068 3080
rect 27120 3068 27126 3120
rect 27448 3117 27476 3148
rect 27433 3111 27491 3117
rect 27433 3077 27445 3111
rect 27479 3077 27491 3111
rect 27433 3071 27491 3077
rect 28718 3068 28724 3120
rect 28776 3108 28782 3120
rect 31220 3108 31248 3148
rect 31294 3136 31300 3188
rect 31352 3176 31358 3188
rect 31352 3148 34744 3176
rect 31352 3136 31358 3148
rect 32674 3108 32680 3120
rect 28776 3080 30406 3108
rect 31220 3080 32680 3108
rect 28776 3068 28782 3080
rect 32674 3068 32680 3080
rect 32732 3068 32738 3120
rect 34422 3108 34428 3120
rect 33810 3080 34428 3108
rect 34422 3068 34428 3080
rect 34480 3068 34486 3120
rect 34606 3108 34612 3120
rect 34567 3080 34612 3108
rect 34606 3068 34612 3080
rect 34664 3068 34670 3120
rect 34716 3117 34744 3148
rect 34701 3111 34759 3117
rect 34701 3077 34713 3111
rect 34747 3077 34759 3111
rect 34701 3071 34759 3077
rect 34790 3068 34796 3120
rect 34848 3108 34854 3120
rect 35621 3111 35679 3117
rect 35621 3108 35633 3111
rect 34848 3080 35633 3108
rect 34848 3068 34854 3080
rect 35621 3077 35633 3080
rect 35667 3077 35679 3111
rect 35621 3071 35679 3077
rect 16132 3012 16436 3040
rect 19245 3043 19303 3049
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 4948 2944 6009 2972
rect 4948 2932 4954 2944
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 6788 2944 7113 2972
rect 6788 2932 6794 2944
rect 7101 2941 7113 2944
rect 7147 2972 7159 2975
rect 9306 2972 9312 2984
rect 7147 2944 9312 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 9582 2972 9588 2984
rect 9543 2944 9588 2972
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 11020 2944 13829 2972
rect 11020 2932 11026 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 13817 2935 13875 2941
rect 14292 2944 14565 2972
rect 6914 2904 6920 2916
rect 1084 2876 3556 2904
rect 5920 2876 6920 2904
rect 1084 2864 1090 2876
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 2961 2839 3019 2845
rect 2961 2836 2973 2839
rect 992 2808 2973 2836
rect 992 2796 998 2808
rect 2961 2805 2973 2808
rect 3007 2805 3019 2839
rect 2961 2799 3019 2805
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 5920 2836 5948 2876
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 11606 2904 11612 2916
rect 10612 2876 11612 2904
rect 3743 2808 5948 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 6052 2808 8861 2836
rect 6052 2796 6058 2808
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 8849 2799 8907 2805
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 10612 2836 10640 2876
rect 11606 2864 11612 2876
rect 11664 2864 11670 2916
rect 13078 2864 13084 2916
rect 13136 2904 13142 2916
rect 14292 2904 14320 2944
rect 14553 2941 14565 2944
rect 14599 2972 14611 2975
rect 16132 2972 16160 3012
rect 19245 3009 19257 3043
rect 19291 3009 19303 3043
rect 21634 3040 21640 3052
rect 19245 3003 19303 3009
rect 20732 3012 21640 3040
rect 14599 2944 16160 2972
rect 16301 2975 16359 2981
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 16301 2941 16313 2975
rect 16347 2941 16359 2975
rect 16301 2935 16359 2941
rect 13136 2876 14320 2904
rect 13136 2864 13142 2876
rect 16022 2864 16028 2916
rect 16080 2904 16086 2916
rect 16316 2904 16344 2935
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16816 2944 16865 2972
rect 16816 2932 16822 2944
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 17126 2972 17132 2984
rect 17087 2944 17132 2972
rect 16853 2935 16911 2941
rect 17126 2932 17132 2944
rect 17184 2932 17190 2984
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 20732 2972 20760 3012
rect 21634 3000 21640 3012
rect 21692 3000 21698 3052
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 23842 3000 23848 3052
rect 23900 3040 23906 3052
rect 24210 3040 24216 3052
rect 23900 3012 24216 3040
rect 23900 3000 23906 3012
rect 24210 3000 24216 3012
rect 24268 3000 24274 3052
rect 26418 3040 26424 3052
rect 26379 3012 26424 3040
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 36354 3040 36360 3052
rect 17276 2944 20760 2972
rect 17276 2932 17282 2944
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 22278 2972 22284 2984
rect 20864 2944 21220 2972
rect 22239 2944 22284 2972
rect 20864 2932 20870 2944
rect 18966 2904 18972 2916
rect 16080 2876 16344 2904
rect 18156 2876 18972 2904
rect 16080 2864 16086 2876
rect 9456 2808 10640 2836
rect 11057 2839 11115 2845
rect 9456 2796 9462 2808
rect 11057 2805 11069 2839
rect 11103 2836 11115 2839
rect 11422 2836 11428 2848
rect 11103 2808 11428 2836
rect 11103 2805 11115 2808
rect 11057 2799 11115 2805
rect 11422 2796 11428 2808
rect 11480 2836 11486 2848
rect 12050 2839 12108 2845
rect 12050 2836 12062 2839
rect 11480 2808 12062 2836
rect 11480 2796 11486 2808
rect 12050 2805 12062 2808
rect 12096 2805 12108 2839
rect 12050 2799 12108 2805
rect 12250 2796 12256 2848
rect 12308 2836 12314 2848
rect 17678 2836 17684 2848
rect 12308 2808 17684 2836
rect 12308 2796 12314 2808
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 17770 2796 17776 2848
rect 17828 2836 17834 2848
rect 18156 2836 18184 2876
rect 18966 2864 18972 2876
rect 19024 2864 19030 2916
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 21082 2904 21088 2916
rect 20772 2876 21088 2904
rect 20772 2864 20778 2876
rect 21082 2864 21088 2876
rect 21140 2864 21146 2916
rect 21192 2904 21220 2944
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 25958 2972 25964 2984
rect 23532 2944 24256 2972
rect 25919 2944 25964 2972
rect 23532 2932 23538 2944
rect 24118 2904 24124 2916
rect 21192 2876 22094 2904
rect 17828 2808 18184 2836
rect 17828 2796 17834 2808
rect 18230 2796 18236 2848
rect 18288 2836 18294 2848
rect 18601 2839 18659 2845
rect 18601 2836 18613 2839
rect 18288 2808 18613 2836
rect 18288 2796 18294 2808
rect 18601 2805 18613 2808
rect 18647 2805 18659 2839
rect 18601 2799 18659 2805
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 20898 2836 20904 2848
rect 19300 2808 20904 2836
rect 19300 2796 19306 2808
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 22066 2836 22094 2876
rect 23308 2876 24124 2904
rect 23308 2836 23336 2876
rect 24118 2864 24124 2876
rect 24176 2864 24182 2916
rect 22066 2808 23336 2836
rect 23753 2839 23811 2845
rect 23753 2805 23765 2839
rect 23799 2836 23811 2839
rect 24026 2836 24032 2848
rect 23799 2808 24032 2836
rect 23799 2805 23811 2808
rect 23753 2799 23811 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 24228 2836 24256 2944
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 27154 2972 27160 2984
rect 27115 2944 27160 2972
rect 27154 2932 27160 2944
rect 27212 2932 27218 2984
rect 27430 2932 27436 2984
rect 27488 2972 27494 2984
rect 27982 2972 27988 2984
rect 27488 2944 27988 2972
rect 27488 2932 27494 2944
rect 27982 2932 27988 2944
rect 28040 2932 28046 2984
rect 28552 2904 28580 3026
rect 35452 3012 36216 3040
rect 36315 3012 36360 3040
rect 28626 2932 28632 2984
rect 28684 2972 28690 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 28684 2944 29193 2972
rect 28684 2932 28690 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29638 2972 29644 2984
rect 29599 2944 29644 2972
rect 29181 2935 29239 2941
rect 29638 2932 29644 2944
rect 29696 2932 29702 2984
rect 29914 2972 29920 2984
rect 29875 2944 29920 2972
rect 29914 2932 29920 2944
rect 29972 2932 29978 2984
rect 31389 2975 31447 2981
rect 31389 2941 31401 2975
rect 31435 2972 31447 2975
rect 31478 2972 31484 2984
rect 31435 2944 31484 2972
rect 31435 2941 31447 2944
rect 31389 2935 31447 2941
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 32306 2972 32312 2984
rect 32267 2944 32312 2972
rect 32306 2932 32312 2944
rect 32364 2932 32370 2984
rect 32585 2975 32643 2981
rect 32585 2941 32597 2975
rect 32631 2972 32643 2975
rect 33594 2972 33600 2984
rect 32631 2944 33600 2972
rect 32631 2941 32643 2944
rect 32585 2935 32643 2941
rect 33594 2932 33600 2944
rect 33652 2932 33658 2984
rect 35452 2972 35480 3012
rect 33888 2944 35480 2972
rect 36081 2975 36139 2981
rect 28552 2876 29776 2904
rect 26970 2836 26976 2848
rect 24228 2808 26976 2836
rect 26970 2796 26976 2808
rect 27028 2796 27034 2848
rect 27154 2796 27160 2848
rect 27212 2836 27218 2848
rect 29638 2836 29644 2848
rect 27212 2808 29644 2836
rect 27212 2796 27218 2808
rect 29638 2796 29644 2808
rect 29696 2796 29702 2848
rect 29748 2836 29776 2876
rect 30374 2836 30380 2848
rect 29748 2808 30380 2836
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 31570 2796 31576 2848
rect 31628 2836 31634 2848
rect 33888 2836 33916 2944
rect 36081 2941 36093 2975
rect 36127 2941 36139 2975
rect 36188 2972 36216 3012
rect 36354 3000 36360 3012
rect 36412 3000 36418 3052
rect 37734 3040 37740 3052
rect 37695 3012 37740 3040
rect 37734 3000 37740 3012
rect 37792 3000 37798 3052
rect 37461 2975 37519 2981
rect 37461 2972 37473 2975
rect 36188 2944 37473 2972
rect 36081 2935 36139 2941
rect 37461 2941 37473 2944
rect 37507 2941 37519 2975
rect 37461 2935 37519 2941
rect 34146 2864 34152 2916
rect 34204 2904 34210 2916
rect 36096 2904 36124 2935
rect 34204 2876 36124 2904
rect 34204 2864 34210 2876
rect 34054 2836 34060 2848
rect 31628 2808 33916 2836
rect 34015 2808 34060 2836
rect 31628 2796 31634 2808
rect 34054 2796 34060 2808
rect 34112 2796 34118 2848
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 37458 2836 37464 2848
rect 34848 2808 37464 2836
rect 34848 2796 34854 2808
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 4522 2632 4528 2644
rect 1903 2604 4528 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 6178 2632 6184 2644
rect 5040 2604 6184 2632
rect 5040 2592 5046 2604
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 9398 2632 9404 2644
rect 6886 2604 9404 2632
rect 2314 2564 2320 2576
rect 2275 2536 2320 2564
rect 2314 2524 2320 2536
rect 2372 2524 2378 2576
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2533 2651 2567
rect 2593 2527 2651 2533
rect 4341 2567 4399 2573
rect 4341 2533 4353 2567
rect 4387 2564 4399 2567
rect 6886 2564 6914 2604
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 11698 2592 11704 2644
rect 11756 2632 11762 2644
rect 16574 2632 16580 2644
rect 11756 2604 16580 2632
rect 11756 2592 11762 2604
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 16666 2592 16672 2644
rect 16724 2592 16730 2644
rect 28905 2635 28963 2641
rect 16776 2604 28856 2632
rect 4387 2536 6914 2564
rect 11149 2567 11207 2573
rect 4387 2533 4399 2536
rect 4341 2527 4399 2533
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 15933 2567 15991 2573
rect 11195 2536 11836 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 2332 2496 2360 2524
rect 1688 2468 2360 2496
rect 2608 2496 2636 2527
rect 5810 2496 5816 2508
rect 2608 2468 5816 2496
rect 1688 2437 1716 2468
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 6362 2496 6368 2508
rect 6043 2468 6368 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6788 2468 6837 2496
rect 6788 2456 6794 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 7101 2499 7159 2505
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 7190 2496 7196 2508
rect 7147 2468 7196 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 7524 2468 8585 2496
rect 7524 2456 7530 2468
rect 8573 2465 8585 2468
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 9306 2456 9312 2508
rect 9364 2496 9370 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 9364 2468 9413 2496
rect 9364 2456 9370 2468
rect 9401 2465 9413 2468
rect 9447 2496 9459 2499
rect 11054 2496 11060 2508
rect 9447 2468 11060 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 11054 2456 11060 2468
rect 11112 2496 11118 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11112 2468 11713 2496
rect 11112 2456 11118 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11808 2496 11836 2536
rect 13188 2536 14320 2564
rect 13188 2496 13216 2536
rect 14182 2496 14188 2508
rect 11808 2468 13216 2496
rect 14143 2468 14188 2496
rect 11701 2459 11759 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14292 2496 14320 2536
rect 15933 2533 15945 2567
rect 15979 2564 15991 2567
rect 16684 2564 16712 2592
rect 15979 2536 16712 2564
rect 15979 2533 15991 2536
rect 15933 2527 15991 2533
rect 15194 2496 15200 2508
rect 14292 2468 15200 2496
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 1673 2391 1731 2397
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 4154 2428 4160 2440
rect 4115 2400 4160 2428
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11204 2400 11744 2428
rect 11204 2388 11210 2400
rect 4982 2360 4988 2372
rect 4943 2332 4988 2360
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 5132 2332 5177 2360
rect 5132 2320 5138 2332
rect 5350 2320 5356 2372
rect 5408 2360 5414 2372
rect 5408 2332 7052 2360
rect 5408 2320 5414 2332
rect 3329 2295 3387 2301
rect 3329 2261 3341 2295
rect 3375 2292 3387 2295
rect 6914 2292 6920 2304
rect 3375 2264 6920 2292
rect 3375 2261 3387 2264
rect 3329 2255 3387 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7024 2292 7052 2332
rect 7208 2332 7590 2360
rect 7208 2292 7236 2332
rect 9582 2320 9588 2372
rect 9640 2360 9646 2372
rect 9677 2363 9735 2369
rect 9677 2360 9689 2363
rect 9640 2332 9689 2360
rect 9640 2320 9646 2332
rect 9677 2329 9689 2332
rect 9723 2329 9735 2363
rect 11716 2360 11744 2400
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 10902 2332 11284 2360
rect 11716 2332 11989 2360
rect 9677 2323 9735 2329
rect 7024 2264 7236 2292
rect 11256 2292 11284 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 12526 2320 12532 2372
rect 12584 2320 12590 2372
rect 13722 2360 13728 2372
rect 13683 2332 13728 2360
rect 13722 2320 13728 2332
rect 13780 2320 13786 2372
rect 14458 2360 14464 2372
rect 14419 2332 14464 2360
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 16776 2360 16804 2604
rect 28828 2564 28856 2604
rect 28905 2601 28917 2635
rect 28951 2632 28963 2635
rect 29454 2632 29460 2644
rect 28951 2604 29460 2632
rect 28951 2601 28963 2604
rect 28905 2595 28963 2601
rect 29454 2592 29460 2604
rect 29512 2592 29518 2644
rect 34238 2632 34244 2644
rect 29564 2604 34244 2632
rect 29564 2564 29592 2604
rect 34238 2592 34244 2604
rect 34296 2592 34302 2644
rect 28828 2536 29592 2564
rect 34057 2567 34115 2573
rect 34057 2533 34069 2567
rect 34103 2564 34115 2567
rect 34103 2536 35020 2564
rect 34103 2533 34115 2536
rect 34057 2527 34115 2533
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 16908 2468 19441 2496
rect 16908 2456 16914 2468
rect 19429 2465 19441 2468
rect 19475 2496 19487 2499
rect 20162 2496 20168 2508
rect 19475 2468 20168 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 20162 2456 20168 2468
rect 20220 2456 20226 2508
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 22005 2499 22063 2505
rect 22005 2496 22017 2499
rect 20956 2468 22017 2496
rect 20956 2456 20962 2468
rect 22005 2465 22017 2468
rect 22051 2465 22063 2499
rect 22005 2459 22063 2465
rect 22281 2499 22339 2505
rect 22281 2465 22293 2499
rect 22327 2496 22339 2499
rect 23566 2496 23572 2508
rect 22327 2468 23572 2496
rect 22327 2465 22339 2468
rect 22281 2459 22339 2465
rect 23566 2456 23572 2468
rect 23624 2456 23630 2508
rect 23842 2456 23848 2508
rect 23900 2496 23906 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23900 2468 24593 2496
rect 23900 2456 23906 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 24627 2468 27169 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 27157 2459 27215 2465
rect 29638 2456 29644 2508
rect 29696 2496 29702 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29696 2468 29745 2496
rect 29696 2456 29702 2468
rect 29733 2465 29745 2468
rect 29779 2496 29791 2499
rect 32306 2496 32312 2508
rect 29779 2468 32312 2496
rect 29779 2465 29791 2468
rect 29733 2459 29791 2465
rect 32306 2456 32312 2468
rect 32364 2496 32370 2508
rect 34885 2499 34943 2505
rect 34885 2496 34897 2499
rect 32364 2468 34897 2496
rect 32364 2456 32370 2468
rect 34885 2465 34897 2468
rect 34931 2465 34943 2499
rect 34992 2496 35020 2536
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 34992 2468 35173 2496
rect 34885 2459 34943 2465
rect 35161 2465 35173 2468
rect 35207 2496 35219 2499
rect 35526 2496 35532 2508
rect 35207 2468 35532 2496
rect 35207 2465 35219 2468
rect 35161 2459 35219 2465
rect 35526 2456 35532 2468
rect 35584 2456 35590 2508
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 37642 2456 37648 2508
rect 37700 2496 37706 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 37700 2468 37749 2496
rect 37700 2456 37706 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 15686 2332 16804 2360
rect 17129 2363 17187 2369
rect 17129 2329 17141 2363
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 12066 2292 12072 2304
rect 11256 2264 12072 2292
rect 12066 2252 12072 2264
rect 12124 2252 12130 2304
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2292 16359 2295
rect 17144 2292 17172 2323
rect 17586 2320 17592 2372
rect 17644 2320 17650 2372
rect 18874 2360 18880 2372
rect 18835 2332 18880 2360
rect 18874 2320 18880 2332
rect 18932 2320 18938 2372
rect 19705 2363 19763 2369
rect 19705 2329 19717 2363
rect 19751 2329 19763 2363
rect 21358 2360 21364 2372
rect 20930 2332 21364 2360
rect 19705 2323 19763 2329
rect 17218 2292 17224 2304
rect 16347 2264 17224 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 19720 2292 19748 2323
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 21453 2363 21511 2369
rect 21453 2329 21465 2363
rect 21499 2360 21511 2363
rect 22278 2360 22284 2372
rect 21499 2332 22284 2360
rect 21499 2329 21511 2332
rect 21453 2323 21511 2329
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 23290 2320 23296 2372
rect 23348 2320 23354 2372
rect 23658 2320 23664 2372
rect 23716 2360 23722 2372
rect 23716 2332 23888 2360
rect 23716 2320 23722 2332
rect 20714 2292 20720 2304
rect 19720 2264 20720 2292
rect 20714 2252 20720 2264
rect 20772 2252 20778 2304
rect 23750 2292 23756 2304
rect 23711 2264 23756 2292
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 23860 2292 23888 2332
rect 24118 2320 24124 2372
rect 24176 2360 24182 2372
rect 24854 2360 24860 2372
rect 24176 2332 24860 2360
rect 24176 2320 24182 2332
rect 24854 2320 24860 2332
rect 24912 2320 24918 2372
rect 27430 2360 27436 2372
rect 24964 2332 25346 2360
rect 26344 2332 27436 2360
rect 24964 2292 24992 2332
rect 26344 2301 26372 2332
rect 27430 2320 27436 2332
rect 27488 2320 27494 2372
rect 29914 2360 29920 2372
rect 28658 2332 29920 2360
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 30006 2320 30012 2372
rect 30064 2360 30070 2372
rect 31294 2360 31300 2372
rect 30064 2332 30109 2360
rect 31234 2332 31300 2360
rect 30064 2320 30070 2332
rect 31294 2320 31300 2332
rect 31352 2320 31358 2372
rect 32585 2363 32643 2369
rect 32585 2329 32597 2363
rect 32631 2329 32643 2363
rect 34698 2360 34704 2372
rect 33810 2332 34704 2360
rect 32585 2323 32643 2329
rect 23860 2264 24992 2292
rect 26329 2295 26387 2301
rect 26329 2261 26341 2295
rect 26375 2261 26387 2295
rect 26329 2255 26387 2261
rect 28350 2252 28356 2304
rect 28408 2292 28414 2304
rect 31481 2295 31539 2301
rect 31481 2292 31493 2295
rect 28408 2264 31493 2292
rect 28408 2252 28414 2264
rect 31481 2261 31493 2264
rect 31527 2292 31539 2295
rect 32600 2292 32628 2323
rect 34698 2320 34704 2332
rect 34756 2320 34762 2372
rect 36446 2360 36452 2372
rect 36386 2332 36452 2360
rect 36446 2320 36452 2332
rect 36504 2320 36510 2372
rect 36630 2292 36636 2304
rect 31527 2264 32628 2292
rect 36591 2264 36636 2292
rect 31527 2261 31539 2264
rect 31481 2255 31539 2261
rect 36630 2252 36636 2264
rect 36688 2252 36694 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 22646 2088 22652 2100
rect 4120 2060 22652 2088
rect 4120 2048 4126 2060
rect 22646 2048 22652 2060
rect 22704 2048 22710 2100
rect 23750 2048 23756 2100
rect 23808 2088 23814 2100
rect 24762 2088 24768 2100
rect 23808 2060 24768 2088
rect 23808 2048 23814 2060
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
rect 29914 2048 29920 2100
rect 29972 2088 29978 2100
rect 32766 2088 32772 2100
rect 29972 2060 32772 2088
rect 29972 2048 29978 2060
rect 32766 2048 32772 2060
rect 32824 2048 32830 2100
rect 36630 2088 36636 2100
rect 35866 2060 36636 2088
rect 2682 1980 2688 2032
rect 2740 2020 2746 2032
rect 5074 2020 5080 2032
rect 2740 1992 5080 2020
rect 2740 1980 2746 1992
rect 5074 1980 5080 1992
rect 5132 1980 5138 2032
rect 6914 1980 6920 2032
rect 6972 2020 6978 2032
rect 10318 2020 10324 2032
rect 6972 1992 10324 2020
rect 6972 1980 6978 1992
rect 10318 1980 10324 1992
rect 10376 1980 10382 2032
rect 10686 1980 10692 2032
rect 10744 2020 10750 2032
rect 13722 2020 13728 2032
rect 10744 1992 13728 2020
rect 10744 1980 10750 1992
rect 13722 1980 13728 1992
rect 13780 2020 13786 2032
rect 17126 2020 17132 2032
rect 13780 1992 17132 2020
rect 13780 1980 13786 1992
rect 17126 1980 17132 1992
rect 17184 1980 17190 2032
rect 17218 1980 17224 2032
rect 17276 2020 17282 2032
rect 26694 2020 26700 2032
rect 17276 1992 26700 2020
rect 17276 1980 17282 1992
rect 26694 1980 26700 1992
rect 26752 2020 26758 2032
rect 34054 2020 34060 2032
rect 26752 1992 34060 2020
rect 26752 1980 26758 1992
rect 34054 1980 34060 1992
rect 34112 1980 34118 2032
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 11698 1952 11704 1964
rect 3844 1924 11704 1952
rect 3844 1912 3850 1924
rect 11698 1912 11704 1924
rect 11756 1912 11762 1964
rect 14458 1912 14464 1964
rect 14516 1952 14522 1964
rect 16574 1952 16580 1964
rect 14516 1924 16580 1952
rect 14516 1912 14522 1924
rect 16574 1912 16580 1924
rect 16632 1912 16638 1964
rect 16666 1912 16672 1964
rect 16724 1952 16730 1964
rect 16724 1924 17724 1952
rect 16724 1912 16730 1924
rect 14090 1844 14096 1896
rect 14148 1884 14154 1896
rect 17586 1884 17592 1896
rect 14148 1856 17592 1884
rect 14148 1844 14154 1856
rect 17586 1844 17592 1856
rect 17644 1844 17650 1896
rect 17696 1884 17724 1924
rect 21358 1912 21364 1964
rect 21416 1952 21422 1964
rect 21416 1924 26234 1952
rect 21416 1912 21422 1924
rect 22278 1884 22284 1896
rect 17696 1856 22284 1884
rect 22278 1844 22284 1856
rect 22336 1844 22342 1896
rect 9582 1776 9588 1828
rect 9640 1816 9646 1828
rect 18230 1816 18236 1828
rect 9640 1788 18236 1816
rect 9640 1776 9646 1788
rect 18230 1776 18236 1788
rect 18288 1776 18294 1828
rect 26206 1816 26234 1924
rect 27614 1912 27620 1964
rect 27672 1952 27678 1964
rect 28442 1952 28448 1964
rect 27672 1924 28448 1952
rect 27672 1912 27678 1924
rect 28442 1912 28448 1924
rect 28500 1952 28506 1964
rect 35866 1952 35894 2060
rect 36630 2048 36636 2060
rect 36688 2048 36694 2100
rect 28500 1924 35894 1952
rect 28500 1912 28506 1924
rect 39022 1816 39028 1828
rect 26206 1788 39028 1816
rect 39022 1776 39028 1788
rect 39080 1776 39086 1828
rect 3142 1708 3148 1760
rect 3200 1748 3206 1760
rect 18506 1748 18512 1760
rect 3200 1720 18512 1748
rect 3200 1708 3206 1720
rect 18506 1708 18512 1720
rect 18564 1708 18570 1760
rect 11330 1640 11336 1692
rect 11388 1680 11394 1692
rect 18874 1680 18880 1692
rect 11388 1652 18880 1680
rect 11388 1640 11394 1652
rect 18874 1640 18880 1652
rect 18932 1640 18938 1692
rect 16574 1572 16580 1624
rect 16632 1612 16638 1624
rect 23750 1612 23756 1624
rect 16632 1584 23756 1612
rect 16632 1572 16638 1584
rect 23750 1572 23756 1584
rect 23808 1572 23814 1624
rect 29638 1572 29644 1624
rect 29696 1612 29702 1624
rect 36998 1612 37004 1624
rect 29696 1584 37004 1612
rect 29696 1572 29702 1584
rect 36998 1572 37004 1584
rect 37056 1572 37062 1624
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 2498 1340 2504 1352
rect 72 1312 2504 1340
rect 72 1300 78 1312
rect 2498 1300 2504 1312
rect 2556 1300 2562 1352
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20 37272 72 37324
rect 2964 37272 3016 37324
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 15476 37315 15528 37324
rect 15476 37281 15485 37315
rect 15485 37281 15519 37315
rect 15519 37281 15528 37315
rect 15476 37272 15528 37281
rect 16856 37272 16908 37324
rect 19432 37272 19484 37324
rect 23848 37272 23900 37324
rect 26516 37272 26568 37324
rect 31576 37272 31628 37324
rect 38016 37272 38068 37324
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 3056 37204 3108 37256
rect 3240 37204 3292 37256
rect 5080 37204 5132 37256
rect 5172 37204 5224 37256
rect 6552 37247 6604 37256
rect 6552 37213 6561 37247
rect 6561 37213 6595 37247
rect 6595 37213 6604 37247
rect 6552 37204 6604 37213
rect 7840 37247 7892 37256
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 9680 37204 9732 37256
rect 12164 37204 12216 37256
rect 12992 37204 13044 37256
rect 15752 37247 15804 37256
rect 15752 37213 15761 37247
rect 15761 37213 15795 37247
rect 15795 37213 15804 37247
rect 15752 37204 15804 37213
rect 16120 37204 16172 37256
rect 18052 37204 18104 37256
rect 18604 37247 18656 37256
rect 18604 37213 18613 37247
rect 18613 37213 18647 37247
rect 18647 37213 18656 37247
rect 18604 37204 18656 37213
rect 19984 37247 20036 37256
rect 19984 37213 19993 37247
rect 19993 37213 20027 37247
rect 20027 37213 20036 37247
rect 19984 37204 20036 37213
rect 21180 37204 21232 37256
rect 21272 37204 21324 37256
rect 22468 37204 22520 37256
rect 23204 37204 23256 37256
rect 24032 37204 24084 37256
rect 10508 37136 10560 37188
rect 10692 37136 10744 37188
rect 13360 37136 13412 37188
rect 2780 37068 2832 37120
rect 3976 37111 4028 37120
rect 3976 37077 3985 37111
rect 3985 37077 4019 37111
rect 4019 37077 4028 37111
rect 3976 37068 4028 37077
rect 4620 37068 4672 37120
rect 5356 37111 5408 37120
rect 5356 37077 5365 37111
rect 5365 37077 5399 37111
rect 5399 37077 5408 37111
rect 5356 37068 5408 37077
rect 5816 37068 5868 37120
rect 7748 37068 7800 37120
rect 10968 37068 11020 37120
rect 12440 37068 12492 37120
rect 13544 37068 13596 37120
rect 18696 37068 18748 37120
rect 20076 37068 20128 37120
rect 20720 37068 20772 37120
rect 24400 37136 24452 37188
rect 25780 37204 25832 37256
rect 27528 37204 27580 37256
rect 27712 37204 27764 37256
rect 29000 37204 29052 37256
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 30380 37204 30432 37256
rect 30748 37204 30800 37256
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 34796 37204 34848 37256
rect 34980 37204 35032 37256
rect 36268 37204 36320 37256
rect 22560 37068 22612 37120
rect 22928 37068 22980 37120
rect 26056 37136 26108 37188
rect 24584 37068 24636 37120
rect 25136 37068 25188 37120
rect 27068 37068 27120 37120
rect 28908 37136 28960 37188
rect 29000 37111 29052 37120
rect 29000 37077 29009 37111
rect 29009 37077 29043 37111
rect 29043 37077 29052 37111
rect 29000 37068 29052 37077
rect 29644 37068 29696 37120
rect 30472 37111 30524 37120
rect 30472 37077 30481 37111
rect 30481 37077 30515 37111
rect 30515 37077 30524 37111
rect 30472 37068 30524 37077
rect 33508 37068 33560 37120
rect 34520 37068 34572 37120
rect 35440 37068 35492 37120
rect 36084 37068 36136 37120
rect 37096 37068 37148 37120
rect 39304 37068 39356 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1308 36864 1360 36916
rect 2872 36864 2924 36916
rect 3056 36864 3108 36916
rect 3148 36864 3200 36916
rect 5448 36796 5500 36848
rect 2320 36771 2372 36780
rect 2320 36737 2329 36771
rect 2329 36737 2363 36771
rect 2363 36737 2372 36771
rect 2320 36728 2372 36737
rect 10692 36864 10744 36916
rect 11612 36864 11664 36916
rect 19984 36864 20036 36916
rect 22468 36907 22520 36916
rect 7840 36796 7892 36848
rect 22468 36873 22477 36907
rect 22477 36873 22511 36907
rect 22511 36873 22520 36907
rect 22468 36864 22520 36873
rect 24032 36907 24084 36916
rect 24032 36873 24041 36907
rect 24041 36873 24075 36907
rect 24075 36873 24084 36907
rect 24032 36864 24084 36873
rect 32220 36864 32272 36916
rect 36176 36864 36228 36916
rect 36728 36864 36780 36916
rect 2412 36660 2464 36712
rect 3976 36660 4028 36712
rect 6920 36660 6972 36712
rect 9036 36728 9088 36780
rect 10324 36728 10376 36780
rect 14188 36728 14240 36780
rect 16764 36728 16816 36780
rect 18880 36771 18932 36780
rect 18880 36737 18889 36771
rect 18889 36737 18923 36771
rect 18923 36737 18932 36771
rect 18880 36728 18932 36737
rect 28908 36796 28960 36848
rect 30288 36796 30340 36848
rect 23572 36771 23624 36780
rect 12900 36660 12952 36712
rect 23572 36737 23581 36771
rect 23581 36737 23615 36771
rect 23615 36737 23624 36771
rect 23572 36728 23624 36737
rect 24216 36771 24268 36780
rect 24216 36737 24225 36771
rect 24225 36737 24259 36771
rect 24259 36737 24268 36771
rect 24216 36728 24268 36737
rect 23020 36660 23072 36712
rect 30748 36660 30800 36712
rect 5080 36592 5132 36644
rect 35532 36728 35584 36780
rect 36820 36728 36872 36780
rect 37372 36592 37424 36644
rect 5356 36524 5408 36576
rect 9036 36524 9088 36576
rect 9404 36524 9456 36576
rect 17040 36524 17092 36576
rect 35532 36567 35584 36576
rect 35532 36533 35541 36567
rect 35541 36533 35575 36567
rect 35575 36533 35584 36567
rect 35532 36524 35584 36533
rect 36820 36567 36872 36576
rect 36820 36533 36829 36567
rect 36829 36533 36863 36567
rect 36863 36533 36872 36567
rect 36820 36524 36872 36533
rect 37648 36567 37700 36576
rect 37648 36533 37657 36567
rect 37657 36533 37691 36567
rect 37691 36533 37700 36567
rect 37648 36524 37700 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 664 36320 716 36372
rect 15752 36320 15804 36372
rect 23572 36320 23624 36372
rect 38660 36320 38712 36372
rect 23480 36252 23532 36304
rect 36820 36252 36872 36304
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 2688 36116 2740 36168
rect 2964 36116 3016 36168
rect 7104 36116 7156 36168
rect 36544 36159 36596 36168
rect 36544 36125 36553 36159
rect 36553 36125 36587 36159
rect 36587 36125 36596 36159
rect 36544 36116 36596 36125
rect 37188 36116 37240 36168
rect 2228 36048 2280 36100
rect 5448 36048 5500 36100
rect 16120 36048 16172 36100
rect 37096 36048 37148 36100
rect 37556 36091 37608 36100
rect 37556 36057 37565 36091
rect 37565 36057 37599 36091
rect 37599 36057 37608 36091
rect 37556 36048 37608 36057
rect 5816 35980 5868 36032
rect 6460 35980 6512 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 2320 35819 2372 35828
rect 2320 35785 2329 35819
rect 2329 35785 2363 35819
rect 2363 35785 2372 35819
rect 2320 35776 2372 35785
rect 24216 35776 24268 35828
rect 38292 35776 38344 35828
rect 1860 35640 1912 35692
rect 20352 35708 20404 35760
rect 36728 35640 36780 35692
rect 23480 35572 23532 35624
rect 1768 35479 1820 35488
rect 1768 35445 1777 35479
rect 1777 35445 1811 35479
rect 1811 35445 1820 35479
rect 1768 35436 1820 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 37188 35275 37240 35284
rect 37188 35241 37197 35275
rect 37197 35241 37231 35275
rect 37231 35241 37240 35275
rect 37188 35232 37240 35241
rect 37372 35071 37424 35080
rect 37372 35037 37381 35071
rect 37381 35037 37415 35071
rect 37415 35037 37424 35071
rect 37372 35028 37424 35037
rect 37464 34892 37516 34944
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2596 34688 2648 34740
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 31760 34552 31812 34604
rect 37188 34484 37240 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17132 33804 17184 33856
rect 33600 33804 33652 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 36728 33600 36780 33652
rect 4620 33464 4672 33516
rect 5816 33507 5868 33516
rect 5816 33473 5825 33507
rect 5825 33473 5859 33507
rect 5859 33473 5868 33507
rect 5816 33464 5868 33473
rect 2044 33396 2096 33448
rect 34612 33464 34664 33516
rect 1768 33371 1820 33380
rect 1768 33337 1777 33371
rect 1777 33337 1811 33371
rect 1811 33337 1820 33371
rect 1768 33328 1820 33337
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 8944 33260 8996 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 26056 32895 26108 32904
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 19340 32716 19392 32768
rect 25228 32716 25280 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2688 32512 2740 32564
rect 33324 32512 33376 32564
rect 19340 32487 19392 32496
rect 19340 32453 19349 32487
rect 19349 32453 19383 32487
rect 19383 32453 19392 32487
rect 19340 32444 19392 32453
rect 19984 32444 20036 32496
rect 20352 32487 20404 32496
rect 20352 32453 20361 32487
rect 20361 32453 20395 32487
rect 20395 32453 20404 32487
rect 20352 32444 20404 32453
rect 29000 32376 29052 32428
rect 33140 32376 33192 32428
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 1860 32351 1912 32360
rect 1860 32317 1869 32351
rect 1869 32317 1903 32351
rect 1903 32317 1912 32351
rect 1860 32308 1912 32317
rect 37464 32351 37516 32360
rect 37464 32317 37473 32351
rect 37473 32317 37507 32351
rect 37507 32317 37516 32351
rect 37464 32308 37516 32317
rect 30748 32215 30800 32224
rect 30748 32181 30757 32215
rect 30757 32181 30791 32215
rect 30791 32181 30800 32215
rect 30748 32172 30800 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 9128 31900 9180 31952
rect 14464 31900 14516 31952
rect 38200 31943 38252 31952
rect 38200 31909 38209 31943
rect 38209 31909 38243 31943
rect 38243 31909 38252 31943
rect 38200 31900 38252 31909
rect 1676 31764 1728 31816
rect 6460 31832 6512 31884
rect 10968 31832 11020 31884
rect 6092 31764 6144 31816
rect 9036 31764 9088 31816
rect 9404 31764 9456 31816
rect 14740 31764 14792 31816
rect 38016 31807 38068 31816
rect 38016 31773 38025 31807
rect 38025 31773 38059 31807
rect 38059 31773 38068 31807
rect 38016 31764 38068 31773
rect 1768 31671 1820 31680
rect 1768 31637 1777 31671
rect 1777 31637 1811 31671
rect 1811 31637 1820 31671
rect 1768 31628 1820 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 38016 31424 38068 31476
rect 17132 31399 17184 31408
rect 17132 31365 17141 31399
rect 17141 31365 17175 31399
rect 17175 31365 17184 31399
rect 17132 31356 17184 31365
rect 6920 31288 6972 31340
rect 13820 31288 13872 31340
rect 16580 31288 16632 31340
rect 30472 31288 30524 31340
rect 35440 31288 35492 31340
rect 14464 31263 14516 31272
rect 14464 31229 14473 31263
rect 14473 31229 14507 31263
rect 14507 31229 14516 31263
rect 14464 31220 14516 31229
rect 14832 31220 14884 31272
rect 7380 31084 7432 31136
rect 14924 31127 14976 31136
rect 14924 31093 14933 31127
rect 14933 31093 14967 31127
rect 14967 31093 14976 31127
rect 14924 31084 14976 31093
rect 22100 31084 22152 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4620 30880 4672 30932
rect 12992 30923 13044 30932
rect 12992 30889 13001 30923
rect 13001 30889 13035 30923
rect 13035 30889 13044 30923
rect 12992 30880 13044 30889
rect 21180 30880 21232 30932
rect 14924 30812 14976 30864
rect 8944 30744 8996 30796
rect 12808 30744 12860 30796
rect 14832 30787 14884 30796
rect 14832 30753 14841 30787
rect 14841 30753 14875 30787
rect 14875 30753 14884 30787
rect 14832 30744 14884 30753
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 10692 30676 10744 30728
rect 11060 30651 11112 30660
rect 11060 30617 11069 30651
rect 11069 30617 11103 30651
rect 11103 30617 11112 30651
rect 11060 30608 11112 30617
rect 11612 30608 11664 30660
rect 15384 30676 15436 30728
rect 24400 30676 24452 30728
rect 25596 30608 25648 30660
rect 6736 30540 6788 30592
rect 29092 30540 29144 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 11060 30336 11112 30388
rect 21824 30336 21876 30388
rect 13820 30268 13872 30320
rect 14464 30311 14516 30320
rect 14464 30277 14473 30311
rect 14473 30277 14507 30311
rect 14507 30277 14516 30311
rect 14464 30268 14516 30277
rect 16028 30268 16080 30320
rect 12164 30200 12216 30252
rect 16120 30243 16172 30252
rect 15108 30132 15160 30184
rect 14924 30064 14976 30116
rect 16120 30209 16129 30243
rect 16129 30209 16163 30243
rect 16163 30209 16172 30243
rect 16120 30200 16172 30209
rect 15016 29996 15068 30048
rect 16304 30064 16356 30116
rect 18880 30268 18932 30320
rect 21916 30268 21968 30320
rect 23480 30200 23532 30252
rect 26700 30268 26752 30320
rect 26792 30268 26844 30320
rect 38108 30243 38160 30252
rect 22100 30175 22152 30184
rect 22100 30141 22109 30175
rect 22109 30141 22143 30175
rect 22143 30141 22152 30175
rect 23112 30175 23164 30184
rect 22100 30132 22152 30141
rect 23112 30141 23121 30175
rect 23121 30141 23155 30175
rect 23155 30141 23164 30175
rect 23112 30132 23164 30141
rect 25504 30132 25556 30184
rect 38108 30209 38117 30243
rect 38117 30209 38151 30243
rect 38151 30209 38160 30243
rect 38108 30200 38160 30209
rect 29092 30175 29144 30184
rect 29092 30141 29101 30175
rect 29101 30141 29135 30175
rect 29135 30141 29144 30175
rect 29092 30132 29144 30141
rect 35348 30132 35400 30184
rect 31116 30064 31168 30116
rect 38292 30107 38344 30116
rect 38292 30073 38301 30107
rect 38301 30073 38335 30107
rect 38335 30073 38344 30107
rect 38292 30064 38344 30073
rect 17316 29996 17368 30048
rect 23664 30039 23716 30048
rect 23664 30005 23673 30039
rect 23673 30005 23707 30039
rect 23707 30005 23716 30039
rect 23664 29996 23716 30005
rect 23756 29996 23808 30048
rect 24860 29996 24912 30048
rect 26884 29996 26936 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 10692 29835 10744 29844
rect 10692 29801 10701 29835
rect 10701 29801 10735 29835
rect 10735 29801 10744 29835
rect 10692 29792 10744 29801
rect 15384 29835 15436 29844
rect 9496 29724 9548 29776
rect 11152 29724 11204 29776
rect 2596 29656 2648 29708
rect 6368 29588 6420 29640
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 9312 29631 9364 29640
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 10968 29588 11020 29640
rect 13360 29631 13412 29640
rect 13360 29597 13369 29631
rect 13369 29597 13403 29631
rect 13403 29597 13412 29631
rect 13360 29588 13412 29597
rect 15384 29801 15393 29835
rect 15393 29801 15427 29835
rect 15427 29801 15436 29835
rect 15384 29792 15436 29801
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 18604 29792 18656 29844
rect 21916 29835 21968 29844
rect 21916 29801 21925 29835
rect 21925 29801 21959 29835
rect 21959 29801 21968 29835
rect 21916 29792 21968 29801
rect 26792 29835 26844 29844
rect 26792 29801 26801 29835
rect 26801 29801 26835 29835
rect 26835 29801 26844 29835
rect 26792 29792 26844 29801
rect 15108 29656 15160 29708
rect 23204 29656 23256 29708
rect 17040 29631 17092 29640
rect 13636 29520 13688 29572
rect 17040 29597 17049 29631
rect 17049 29597 17083 29631
rect 17083 29597 17092 29631
rect 17040 29588 17092 29597
rect 18236 29631 18288 29640
rect 18236 29597 18245 29631
rect 18245 29597 18279 29631
rect 18279 29597 18288 29631
rect 18236 29588 18288 29597
rect 21456 29588 21508 29640
rect 22744 29588 22796 29640
rect 23020 29631 23072 29640
rect 23020 29597 23029 29631
rect 23029 29597 23063 29631
rect 23063 29597 23072 29631
rect 23020 29588 23072 29597
rect 23572 29588 23624 29640
rect 16764 29520 16816 29572
rect 1768 29495 1820 29504
rect 1768 29461 1777 29495
rect 1777 29461 1811 29495
rect 1811 29461 1820 29495
rect 1768 29452 1820 29461
rect 9772 29495 9824 29504
rect 9772 29461 9781 29495
rect 9781 29461 9815 29495
rect 9815 29461 9824 29495
rect 9772 29452 9824 29461
rect 14004 29452 14056 29504
rect 15108 29452 15160 29504
rect 18696 29452 18748 29504
rect 23388 29452 23440 29504
rect 24032 29452 24084 29504
rect 25228 29699 25280 29708
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 26700 29631 26752 29640
rect 26700 29597 26709 29631
rect 26709 29597 26743 29631
rect 26743 29597 26752 29631
rect 26700 29588 26752 29597
rect 38016 29631 38068 29640
rect 38016 29597 38025 29631
rect 38025 29597 38059 29631
rect 38059 29597 38068 29631
rect 38016 29588 38068 29597
rect 25320 29563 25372 29572
rect 25320 29529 25329 29563
rect 25329 29529 25363 29563
rect 25363 29529 25372 29563
rect 25320 29520 25372 29529
rect 25504 29520 25556 29572
rect 29736 29452 29788 29504
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9312 29291 9364 29300
rect 9312 29257 9321 29291
rect 9321 29257 9355 29291
rect 9355 29257 9364 29291
rect 9312 29248 9364 29257
rect 14648 29248 14700 29300
rect 20628 29248 20680 29300
rect 25320 29291 25372 29300
rect 25320 29257 25329 29291
rect 25329 29257 25363 29291
rect 25363 29257 25372 29291
rect 25320 29248 25372 29257
rect 6644 29112 6696 29164
rect 11152 29112 11204 29164
rect 11336 29112 11388 29164
rect 9680 29044 9732 29096
rect 15016 29155 15068 29164
rect 15016 29121 15025 29155
rect 15025 29121 15059 29155
rect 15059 29121 15068 29155
rect 15016 29112 15068 29121
rect 14832 29087 14884 29096
rect 1768 29019 1820 29028
rect 1768 28985 1777 29019
rect 1777 28985 1811 29019
rect 1811 28985 1820 29019
rect 1768 28976 1820 28985
rect 12256 28976 12308 29028
rect 14832 29053 14841 29087
rect 14841 29053 14875 29087
rect 14875 29053 14884 29087
rect 14832 29044 14884 29053
rect 21824 29180 21876 29232
rect 15844 29112 15896 29164
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 23480 29180 23532 29232
rect 23756 29223 23808 29232
rect 23756 29189 23765 29223
rect 23765 29189 23799 29223
rect 23799 29189 23808 29223
rect 23756 29180 23808 29189
rect 23940 29180 23992 29232
rect 20904 29112 20956 29121
rect 20628 29044 20680 29096
rect 25228 29155 25280 29164
rect 25228 29121 25237 29155
rect 25237 29121 25271 29155
rect 25271 29121 25280 29155
rect 25228 29112 25280 29121
rect 27988 29180 28040 29232
rect 30748 29180 30800 29232
rect 31024 29223 31076 29232
rect 31024 29189 31033 29223
rect 31033 29189 31067 29223
rect 31067 29189 31076 29223
rect 31024 29180 31076 29189
rect 28908 29112 28960 29164
rect 23664 29087 23716 29096
rect 23664 29053 23673 29087
rect 23673 29053 23707 29087
rect 23707 29053 23716 29087
rect 23664 29044 23716 29053
rect 23756 29044 23808 29096
rect 15292 28976 15344 29028
rect 11520 28908 11572 28960
rect 11888 28908 11940 28960
rect 15660 28908 15712 28960
rect 16120 28908 16172 28960
rect 16396 28908 16448 28960
rect 20904 28908 20956 28960
rect 21272 28908 21324 28960
rect 22836 28976 22888 29028
rect 27252 29019 27304 29028
rect 27252 28985 27261 29019
rect 27261 28985 27295 29019
rect 27295 28985 27304 29019
rect 27252 28976 27304 28985
rect 31116 28976 31168 29028
rect 37188 29044 37240 29096
rect 37740 29087 37792 29096
rect 37740 29053 37749 29087
rect 37749 29053 37783 29087
rect 37783 29053 37792 29087
rect 37740 29044 37792 29053
rect 35532 28976 35584 29028
rect 23480 28908 23532 28960
rect 26148 28908 26200 28960
rect 26332 28951 26384 28960
rect 26332 28917 26341 28951
rect 26341 28917 26375 28951
rect 26375 28917 26384 28951
rect 26332 28908 26384 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6368 28747 6420 28756
rect 6368 28713 6377 28747
rect 6377 28713 6411 28747
rect 6411 28713 6420 28747
rect 6368 28704 6420 28713
rect 9772 28704 9824 28756
rect 10876 28704 10928 28756
rect 9128 28568 9180 28620
rect 6736 28500 6788 28552
rect 11060 28500 11112 28552
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 16028 28636 16080 28688
rect 14832 28568 14884 28620
rect 14556 28500 14608 28552
rect 7472 28364 7524 28416
rect 11428 28432 11480 28484
rect 11520 28475 11572 28484
rect 11520 28441 11529 28475
rect 11529 28441 11563 28475
rect 11563 28441 11572 28475
rect 11520 28432 11572 28441
rect 12440 28475 12492 28484
rect 12440 28441 12449 28475
rect 12449 28441 12483 28475
rect 12483 28441 12492 28475
rect 12440 28432 12492 28441
rect 14464 28432 14516 28484
rect 14740 28432 14792 28484
rect 15016 28475 15068 28484
rect 15016 28441 15025 28475
rect 15025 28441 15059 28475
rect 15059 28441 15068 28475
rect 15016 28432 15068 28441
rect 15108 28475 15160 28484
rect 15108 28441 15117 28475
rect 15117 28441 15151 28475
rect 15151 28441 15160 28475
rect 15108 28432 15160 28441
rect 15292 28432 15344 28484
rect 17316 28704 17368 28756
rect 16212 28568 16264 28620
rect 19432 28636 19484 28688
rect 20260 28636 20312 28688
rect 22008 28704 22060 28756
rect 31024 28636 31076 28688
rect 33140 28636 33192 28688
rect 16764 28543 16816 28552
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 20076 28611 20128 28620
rect 20076 28577 20085 28611
rect 20085 28577 20119 28611
rect 20119 28577 20128 28611
rect 20076 28568 20128 28577
rect 20352 28568 20404 28620
rect 21364 28568 21416 28620
rect 19340 28500 19392 28552
rect 22744 28500 22796 28552
rect 24216 28500 24268 28552
rect 25136 28500 25188 28552
rect 26148 28568 26200 28620
rect 37740 28568 37792 28620
rect 32128 28500 32180 28552
rect 12900 28364 12952 28416
rect 14188 28364 14240 28416
rect 14372 28407 14424 28416
rect 14372 28373 14381 28407
rect 14381 28373 14415 28407
rect 14415 28373 14424 28407
rect 14372 28364 14424 28373
rect 17776 28432 17828 28484
rect 15752 28364 15804 28416
rect 16028 28364 16080 28416
rect 16856 28407 16908 28416
rect 16856 28373 16865 28407
rect 16865 28373 16899 28407
rect 16899 28373 16908 28407
rect 16856 28364 16908 28373
rect 19432 28364 19484 28416
rect 21272 28475 21324 28484
rect 21272 28441 21281 28475
rect 21281 28441 21315 28475
rect 21315 28441 21324 28475
rect 21272 28432 21324 28441
rect 24032 28432 24084 28484
rect 25044 28432 25096 28484
rect 26332 28432 26384 28484
rect 26976 28475 27028 28484
rect 26976 28441 26985 28475
rect 26985 28441 27019 28475
rect 27019 28441 27028 28475
rect 26976 28432 27028 28441
rect 29184 28432 29236 28484
rect 21824 28364 21876 28416
rect 23112 28364 23164 28416
rect 23296 28364 23348 28416
rect 24768 28364 24820 28416
rect 24860 28364 24912 28416
rect 28632 28364 28684 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 6644 28203 6696 28212
rect 6644 28169 6653 28203
rect 6653 28169 6687 28203
rect 6687 28169 6696 28203
rect 6644 28160 6696 28169
rect 14832 28160 14884 28212
rect 1860 28092 1912 28144
rect 8300 28067 8352 28076
rect 8300 28033 8309 28067
rect 8309 28033 8343 28067
rect 8343 28033 8352 28067
rect 8300 28024 8352 28033
rect 9864 28092 9916 28144
rect 13820 28092 13872 28144
rect 11428 28024 11480 28076
rect 11704 28024 11756 28076
rect 12072 28067 12124 28076
rect 12072 28033 12081 28067
rect 12081 28033 12115 28067
rect 12115 28033 12124 28067
rect 12072 28024 12124 28033
rect 13912 28024 13964 28076
rect 9588 27956 9640 28008
rect 10692 27999 10744 28008
rect 10692 27965 10701 27999
rect 10701 27965 10735 27999
rect 10735 27965 10744 27999
rect 10692 27956 10744 27965
rect 12716 27999 12768 28008
rect 12716 27965 12725 27999
rect 12725 27965 12759 27999
rect 12759 27965 12768 27999
rect 12716 27956 12768 27965
rect 13176 27956 13228 28008
rect 13544 27999 13596 28008
rect 13544 27965 13553 27999
rect 13553 27965 13587 27999
rect 13587 27965 13596 27999
rect 13544 27956 13596 27965
rect 16856 28160 16908 28212
rect 22928 28160 22980 28212
rect 16304 28135 16356 28144
rect 16304 28101 16313 28135
rect 16313 28101 16347 28135
rect 16347 28101 16356 28135
rect 16304 28092 16356 28101
rect 17868 28135 17920 28144
rect 17868 28101 17877 28135
rect 17877 28101 17911 28135
rect 17911 28101 17920 28135
rect 17868 28092 17920 28101
rect 23756 28160 23808 28212
rect 29000 28160 29052 28212
rect 23296 28135 23348 28144
rect 23296 28101 23305 28135
rect 23305 28101 23339 28135
rect 23339 28101 23348 28135
rect 23296 28092 23348 28101
rect 24860 28135 24912 28144
rect 24860 28101 24869 28135
rect 24869 28101 24903 28135
rect 24903 28101 24912 28135
rect 24860 28092 24912 28101
rect 25780 28135 25832 28144
rect 25780 28101 25789 28135
rect 25789 28101 25823 28135
rect 25823 28101 25832 28135
rect 25780 28092 25832 28101
rect 28632 28135 28684 28144
rect 28632 28101 28641 28135
rect 28641 28101 28675 28135
rect 28675 28101 28684 28135
rect 28632 28092 28684 28101
rect 29092 28092 29144 28144
rect 30472 28092 30524 28144
rect 16948 28024 17000 28076
rect 18972 28024 19024 28076
rect 19340 28024 19392 28076
rect 20628 28024 20680 28076
rect 20996 28024 21048 28076
rect 21548 28024 21600 28076
rect 22008 28024 22060 28076
rect 26240 28067 26292 28076
rect 26240 28033 26249 28067
rect 26249 28033 26283 28067
rect 26283 28033 26292 28067
rect 26240 28024 26292 28033
rect 26516 28024 26568 28076
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 27712 28024 27764 28076
rect 15660 27999 15712 28008
rect 15660 27965 15669 27999
rect 15669 27965 15703 27999
rect 15703 27965 15712 27999
rect 15660 27956 15712 27965
rect 17776 27999 17828 28008
rect 17776 27965 17785 27999
rect 17785 27965 17819 27999
rect 17819 27965 17828 27999
rect 17776 27956 17828 27965
rect 23388 27956 23440 28008
rect 23756 27999 23808 28008
rect 23756 27965 23765 27999
rect 23765 27965 23799 27999
rect 23799 27965 23808 27999
rect 23756 27956 23808 27965
rect 24584 27956 24636 28008
rect 28080 27956 28132 28008
rect 29000 27999 29052 28008
rect 29000 27965 29009 27999
rect 29009 27965 29043 27999
rect 29043 27965 29052 27999
rect 29000 27956 29052 27965
rect 29552 27956 29604 28008
rect 33968 27956 34020 28008
rect 25504 27888 25556 27940
rect 11980 27820 12032 27872
rect 12164 27863 12216 27872
rect 12164 27829 12173 27863
rect 12173 27829 12207 27863
rect 12207 27829 12216 27863
rect 12164 27820 12216 27829
rect 15660 27820 15712 27872
rect 16948 27863 17000 27872
rect 16948 27829 16957 27863
rect 16957 27829 16991 27863
rect 16991 27829 17000 27863
rect 16948 27820 17000 27829
rect 19340 27863 19392 27872
rect 19340 27829 19349 27863
rect 19349 27829 19383 27863
rect 19383 27829 19392 27863
rect 19340 27820 19392 27829
rect 20444 27820 20496 27872
rect 22192 27863 22244 27872
rect 22192 27829 22201 27863
rect 22201 27829 22235 27863
rect 22235 27829 22244 27863
rect 22192 27820 22244 27829
rect 26424 27820 26476 27872
rect 27896 27863 27948 27872
rect 27896 27829 27905 27863
rect 27905 27829 27939 27863
rect 27939 27829 27948 27863
rect 27896 27820 27948 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 9772 27616 9824 27668
rect 7472 27523 7524 27532
rect 7472 27489 7481 27523
rect 7481 27489 7515 27523
rect 7515 27489 7524 27523
rect 7472 27480 7524 27489
rect 10968 27480 11020 27532
rect 4068 27412 4120 27464
rect 9772 27455 9824 27464
rect 7564 27387 7616 27396
rect 7564 27353 7573 27387
rect 7573 27353 7607 27387
rect 7607 27353 7616 27387
rect 7564 27344 7616 27353
rect 8484 27387 8536 27396
rect 8484 27353 8493 27387
rect 8493 27353 8527 27387
rect 8527 27353 8536 27387
rect 8484 27344 8536 27353
rect 9772 27421 9781 27455
rect 9781 27421 9815 27455
rect 9815 27421 9824 27455
rect 9772 27412 9824 27421
rect 10784 27344 10836 27396
rect 13544 27548 13596 27600
rect 13820 27616 13872 27668
rect 16856 27616 16908 27668
rect 17868 27616 17920 27668
rect 20720 27616 20772 27668
rect 23664 27616 23716 27668
rect 14556 27548 14608 27600
rect 15016 27548 15068 27600
rect 12256 27455 12308 27464
rect 12256 27421 12265 27455
rect 12265 27421 12299 27455
rect 12299 27421 12308 27455
rect 12256 27412 12308 27421
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 12532 27344 12584 27396
rect 13636 27480 13688 27532
rect 16304 27523 16356 27532
rect 16304 27489 16313 27523
rect 16313 27489 16347 27523
rect 16347 27489 16356 27523
rect 16304 27480 16356 27489
rect 11520 27276 11572 27328
rect 14096 27344 14148 27396
rect 14464 27387 14516 27396
rect 14464 27353 14473 27387
rect 14473 27353 14507 27387
rect 14507 27353 14516 27387
rect 14464 27344 14516 27353
rect 15752 27412 15804 27464
rect 16764 27412 16816 27464
rect 15660 27344 15712 27396
rect 15936 27387 15988 27396
rect 15936 27353 15945 27387
rect 15945 27353 15979 27387
rect 15979 27353 15988 27387
rect 15936 27344 15988 27353
rect 15476 27276 15528 27328
rect 16948 27344 17000 27396
rect 19248 27344 19300 27396
rect 21548 27548 21600 27600
rect 21824 27548 21876 27600
rect 26240 27616 26292 27668
rect 30472 27591 30524 27600
rect 20352 27480 20404 27532
rect 20812 27387 20864 27396
rect 19340 27276 19392 27328
rect 20812 27353 20821 27387
rect 20821 27353 20855 27387
rect 20855 27353 20864 27387
rect 20812 27344 20864 27353
rect 23480 27412 23532 27464
rect 23940 27412 23992 27464
rect 21824 27387 21876 27396
rect 21824 27353 21833 27387
rect 21833 27353 21867 27387
rect 21867 27353 21876 27387
rect 21824 27344 21876 27353
rect 22008 27344 22060 27396
rect 25780 27480 25832 27532
rect 30472 27557 30481 27591
rect 30481 27557 30515 27591
rect 30515 27557 30524 27591
rect 30472 27548 30524 27557
rect 33876 27548 33928 27600
rect 26700 27523 26752 27532
rect 26700 27489 26709 27523
rect 26709 27489 26743 27523
rect 26743 27489 26752 27523
rect 26700 27480 26752 27489
rect 27252 27480 27304 27532
rect 28172 27523 28224 27532
rect 28172 27489 28181 27523
rect 28181 27489 28215 27523
rect 28215 27489 28224 27523
rect 28172 27480 28224 27489
rect 27344 27412 27396 27464
rect 24676 27344 24728 27396
rect 24768 27387 24820 27396
rect 24768 27353 24777 27387
rect 24777 27353 24811 27387
rect 24811 27353 24820 27387
rect 24768 27344 24820 27353
rect 25320 27344 25372 27396
rect 26424 27344 26476 27396
rect 27896 27387 27948 27396
rect 27896 27353 27905 27387
rect 27905 27353 27939 27387
rect 27939 27353 27948 27387
rect 31760 27480 31812 27532
rect 29736 27455 29788 27464
rect 29736 27421 29745 27455
rect 29745 27421 29779 27455
rect 29779 27421 29788 27455
rect 29736 27412 29788 27421
rect 30380 27455 30432 27464
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 38292 27455 38344 27464
rect 38292 27421 38301 27455
rect 38301 27421 38335 27455
rect 38335 27421 38344 27455
rect 38292 27412 38344 27421
rect 27896 27344 27948 27353
rect 30472 27344 30524 27396
rect 24400 27276 24452 27328
rect 27712 27276 27764 27328
rect 28080 27276 28132 27328
rect 34520 27276 34572 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8300 27072 8352 27124
rect 9772 27115 9824 27124
rect 9772 27081 9781 27115
rect 9781 27081 9815 27115
rect 9815 27081 9824 27115
rect 9772 27072 9824 27081
rect 10692 27072 10744 27124
rect 11060 27115 11112 27124
rect 11060 27081 11069 27115
rect 11069 27081 11103 27115
rect 11103 27081 11112 27115
rect 11060 27072 11112 27081
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 9680 26979 9732 26988
rect 9680 26945 9689 26979
rect 9689 26945 9723 26979
rect 9723 26945 9732 26979
rect 9680 26936 9732 26945
rect 12256 27004 12308 27056
rect 12348 27004 12400 27056
rect 14556 27047 14608 27056
rect 14556 27013 14565 27047
rect 14565 27013 14599 27047
rect 14599 27013 14608 27047
rect 14556 27004 14608 27013
rect 15108 27072 15160 27124
rect 20352 27072 20404 27124
rect 10692 26936 10744 26988
rect 10876 26936 10928 26988
rect 7380 26868 7432 26920
rect 12164 26936 12216 26988
rect 14096 26936 14148 26988
rect 14280 26936 14332 26988
rect 15844 26936 15896 26988
rect 10784 26732 10836 26784
rect 14004 26868 14056 26920
rect 15016 26868 15068 26920
rect 15384 26868 15436 26920
rect 16948 27004 17000 27056
rect 17592 27004 17644 27056
rect 18788 27047 18840 27056
rect 18788 27013 18797 27047
rect 18797 27013 18831 27047
rect 18831 27013 18840 27047
rect 18788 27004 18840 27013
rect 20444 27004 20496 27056
rect 22376 26936 22428 26988
rect 11980 26800 12032 26852
rect 15936 26800 15988 26852
rect 18236 26868 18288 26920
rect 18696 26911 18748 26920
rect 18696 26877 18705 26911
rect 18705 26877 18739 26911
rect 18739 26877 18748 26911
rect 18696 26868 18748 26877
rect 20720 26868 20772 26920
rect 20904 26911 20956 26920
rect 20904 26877 20913 26911
rect 20913 26877 20947 26911
rect 20947 26877 20956 26911
rect 20904 26868 20956 26877
rect 26608 27072 26660 27124
rect 22836 27047 22888 27056
rect 22836 27013 22845 27047
rect 22845 27013 22879 27047
rect 22879 27013 22888 27047
rect 22836 27004 22888 27013
rect 24676 27047 24728 27056
rect 24676 27013 24685 27047
rect 24685 27013 24719 27047
rect 24719 27013 24728 27047
rect 24676 27004 24728 27013
rect 24768 27004 24820 27056
rect 26884 27004 26936 27056
rect 29736 27072 29788 27124
rect 33324 27115 33376 27124
rect 33324 27081 33333 27115
rect 33333 27081 33367 27115
rect 33367 27081 33376 27115
rect 33324 27072 33376 27081
rect 27344 27004 27396 27056
rect 26424 26936 26476 26988
rect 27436 26936 27488 26988
rect 24584 26911 24636 26920
rect 19064 26800 19116 26852
rect 19248 26843 19300 26852
rect 19248 26809 19257 26843
rect 19257 26809 19291 26843
rect 19291 26809 19300 26843
rect 19248 26800 19300 26809
rect 19524 26800 19576 26852
rect 24584 26877 24593 26911
rect 24593 26877 24627 26911
rect 24627 26877 24636 26911
rect 24584 26868 24636 26877
rect 24860 26911 24912 26920
rect 24860 26877 24869 26911
rect 24869 26877 24903 26911
rect 24903 26877 24912 26911
rect 24860 26868 24912 26877
rect 24492 26800 24544 26852
rect 27344 26868 27396 26920
rect 27160 26800 27212 26852
rect 29460 26936 29512 26988
rect 30380 26936 30432 26988
rect 28080 26911 28132 26920
rect 28080 26877 28089 26911
rect 28089 26877 28123 26911
rect 28123 26877 28132 26911
rect 28080 26868 28132 26877
rect 31944 26868 31996 26920
rect 33600 26936 33652 26988
rect 38292 26979 38344 26988
rect 38292 26945 38301 26979
rect 38301 26945 38335 26979
rect 38335 26945 38344 26979
rect 38292 26936 38344 26945
rect 34704 26868 34756 26920
rect 14832 26732 14884 26784
rect 15844 26732 15896 26784
rect 18052 26732 18104 26784
rect 21180 26732 21232 26784
rect 21364 26732 21416 26784
rect 24768 26732 24820 26784
rect 26792 26732 26844 26784
rect 35348 26800 35400 26852
rect 29368 26732 29420 26784
rect 31300 26732 31352 26784
rect 37280 26732 37332 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 7564 26528 7616 26580
rect 10784 26571 10836 26580
rect 10784 26537 10793 26571
rect 10793 26537 10827 26571
rect 10827 26537 10836 26571
rect 10784 26528 10836 26537
rect 14556 26528 14608 26580
rect 14924 26571 14976 26580
rect 14924 26537 14933 26571
rect 14933 26537 14967 26571
rect 14967 26537 14976 26571
rect 14924 26528 14976 26537
rect 18788 26571 18840 26580
rect 18788 26537 18797 26571
rect 18797 26537 18831 26571
rect 18831 26537 18840 26571
rect 18788 26528 18840 26537
rect 9680 26460 9732 26512
rect 10600 26460 10652 26512
rect 12348 26460 12400 26512
rect 13084 26460 13136 26512
rect 12716 26435 12768 26444
rect 12716 26401 12725 26435
rect 12725 26401 12759 26435
rect 12759 26401 12768 26435
rect 12716 26392 12768 26401
rect 12900 26392 12952 26444
rect 15384 26460 15436 26512
rect 15752 26460 15804 26512
rect 17408 26460 17460 26512
rect 19248 26460 19300 26512
rect 20168 26460 20220 26512
rect 10508 26324 10560 26376
rect 10784 26324 10836 26376
rect 11336 26367 11388 26376
rect 11336 26333 11345 26367
rect 11345 26333 11379 26367
rect 11379 26333 11388 26367
rect 11336 26324 11388 26333
rect 11796 26324 11848 26376
rect 8484 26256 8536 26308
rect 12808 26299 12860 26308
rect 12808 26265 12817 26299
rect 12817 26265 12851 26299
rect 12851 26265 12860 26299
rect 12808 26256 12860 26265
rect 14372 26392 14424 26444
rect 14556 26324 14608 26376
rect 15108 26324 15160 26376
rect 16028 26299 16080 26308
rect 16028 26265 16030 26299
rect 16030 26265 16064 26299
rect 16064 26265 16080 26299
rect 16948 26392 17000 26444
rect 19340 26392 19392 26444
rect 20076 26392 20128 26444
rect 24676 26528 24728 26580
rect 30472 26528 30524 26580
rect 31392 26528 31444 26580
rect 34612 26528 34664 26580
rect 24952 26460 25004 26512
rect 25320 26460 25372 26512
rect 26148 26460 26200 26512
rect 25780 26392 25832 26444
rect 27252 26460 27304 26512
rect 27344 26460 27396 26512
rect 26332 26392 26384 26444
rect 26700 26392 26752 26444
rect 27068 26392 27120 26444
rect 18604 26324 18656 26376
rect 16028 26256 16080 26265
rect 17224 26256 17276 26308
rect 17316 26299 17368 26308
rect 17316 26265 17325 26299
rect 17325 26265 17359 26299
rect 17359 26265 17368 26299
rect 17316 26256 17368 26265
rect 18052 26256 18104 26308
rect 18788 26256 18840 26308
rect 19524 26299 19576 26308
rect 19524 26265 19533 26299
rect 19533 26265 19567 26299
rect 19567 26265 19576 26299
rect 19524 26256 19576 26265
rect 20168 26256 20220 26308
rect 21364 26299 21416 26308
rect 21364 26265 21373 26299
rect 21373 26265 21407 26299
rect 21407 26265 21416 26299
rect 21364 26256 21416 26265
rect 22836 26256 22888 26308
rect 22928 26299 22980 26308
rect 22928 26265 22937 26299
rect 22937 26265 22971 26299
rect 22971 26265 22980 26299
rect 22928 26256 22980 26265
rect 24124 26256 24176 26308
rect 24492 26256 24544 26308
rect 24768 26299 24820 26308
rect 24768 26265 24777 26299
rect 24777 26265 24811 26299
rect 24811 26265 24820 26299
rect 24768 26256 24820 26265
rect 30472 26435 30524 26444
rect 30472 26401 30481 26435
rect 30481 26401 30515 26435
rect 30515 26401 30524 26435
rect 30472 26392 30524 26401
rect 31024 26392 31076 26444
rect 27712 26367 27764 26376
rect 27712 26333 27721 26367
rect 27721 26333 27755 26367
rect 27755 26333 27764 26367
rect 27712 26324 27764 26333
rect 27436 26256 27488 26308
rect 28540 26324 28592 26376
rect 31300 26367 31352 26376
rect 31300 26333 31309 26367
rect 31309 26333 31343 26367
rect 31343 26333 31352 26367
rect 31300 26324 31352 26333
rect 31944 26367 31996 26376
rect 31944 26333 31953 26367
rect 31953 26333 31987 26367
rect 31987 26333 31996 26367
rect 31944 26324 31996 26333
rect 29828 26299 29880 26308
rect 27160 26188 27212 26240
rect 29828 26265 29837 26299
rect 29837 26265 29871 26299
rect 29871 26265 29880 26299
rect 29828 26256 29880 26265
rect 31576 26188 31628 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 12624 25984 12676 26036
rect 12992 25984 13044 26036
rect 12532 25959 12584 25968
rect 12532 25925 12541 25959
rect 12541 25925 12575 25959
rect 12575 25925 12584 25959
rect 12532 25916 12584 25925
rect 15108 25959 15160 25968
rect 15108 25925 15117 25959
rect 15117 25925 15151 25959
rect 15151 25925 15160 25959
rect 15108 25916 15160 25925
rect 17316 25984 17368 26036
rect 17592 26027 17644 26036
rect 17592 25993 17601 26027
rect 17601 25993 17635 26027
rect 17635 25993 17644 26027
rect 17592 25984 17644 25993
rect 17684 25984 17736 26036
rect 13084 25891 13136 25900
rect 13084 25857 13093 25891
rect 13093 25857 13127 25891
rect 13127 25857 13136 25891
rect 13084 25848 13136 25857
rect 10968 25780 11020 25832
rect 11888 25823 11940 25832
rect 11888 25789 11897 25823
rect 11897 25789 11931 25823
rect 11931 25789 11940 25823
rect 11888 25780 11940 25789
rect 17408 25848 17460 25900
rect 20076 25916 20128 25968
rect 10876 25712 10928 25764
rect 14556 25780 14608 25832
rect 15016 25823 15068 25832
rect 15016 25789 15025 25823
rect 15025 25789 15059 25823
rect 15059 25789 15068 25823
rect 15016 25780 15068 25789
rect 15660 25823 15712 25832
rect 15660 25789 15669 25823
rect 15669 25789 15703 25823
rect 15703 25789 15712 25823
rect 15660 25780 15712 25789
rect 14464 25712 14516 25764
rect 17132 25712 17184 25764
rect 19248 25780 19300 25832
rect 20812 25984 20864 26036
rect 22008 25984 22060 26036
rect 20812 25780 20864 25832
rect 21824 25848 21876 25900
rect 23112 25959 23164 25968
rect 23112 25925 23121 25959
rect 23121 25925 23155 25959
rect 23155 25925 23164 25959
rect 23112 25916 23164 25925
rect 24584 25959 24636 25968
rect 24584 25925 24593 25959
rect 24593 25925 24627 25959
rect 24627 25925 24636 25959
rect 24584 25916 24636 25925
rect 26148 25916 26200 25968
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 27528 25984 27580 26036
rect 28908 25916 28960 25968
rect 38016 25984 38068 26036
rect 29736 25916 29788 25968
rect 30104 25916 30156 25968
rect 38200 25916 38252 25968
rect 23388 25780 23440 25832
rect 24032 25823 24084 25832
rect 24032 25789 24041 25823
rect 24041 25789 24075 25823
rect 24075 25789 24084 25823
rect 24032 25780 24084 25789
rect 24952 25823 25004 25832
rect 24952 25789 24961 25823
rect 24961 25789 24995 25823
rect 24995 25789 25004 25823
rect 24952 25780 25004 25789
rect 22928 25712 22980 25764
rect 23112 25712 23164 25764
rect 25504 25780 25556 25832
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 28540 25891 28592 25900
rect 28540 25857 28549 25891
rect 28549 25857 28583 25891
rect 28583 25857 28592 25891
rect 28540 25848 28592 25857
rect 30196 25848 30248 25900
rect 34520 25848 34572 25900
rect 30288 25823 30340 25832
rect 11152 25644 11204 25696
rect 12348 25644 12400 25696
rect 13728 25644 13780 25696
rect 16120 25644 16172 25696
rect 21088 25644 21140 25696
rect 21456 25644 21508 25696
rect 24952 25644 25004 25696
rect 25320 25644 25372 25696
rect 25780 25687 25832 25696
rect 25780 25653 25789 25687
rect 25789 25653 25823 25687
rect 25823 25653 25832 25687
rect 25780 25644 25832 25653
rect 29920 25712 29972 25764
rect 30288 25789 30297 25823
rect 30297 25789 30331 25823
rect 30331 25789 30340 25823
rect 30288 25780 30340 25789
rect 34428 25712 34480 25764
rect 28448 25644 28500 25696
rect 28816 25644 28868 25696
rect 28908 25644 28960 25696
rect 31852 25644 31904 25696
rect 33692 25644 33744 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 10876 25483 10928 25492
rect 10876 25449 10885 25483
rect 10885 25449 10919 25483
rect 10919 25449 10928 25483
rect 10876 25440 10928 25449
rect 11888 25440 11940 25492
rect 13728 25483 13780 25492
rect 13728 25449 13737 25483
rect 13737 25449 13771 25483
rect 13771 25449 13780 25483
rect 13728 25440 13780 25449
rect 14096 25440 14148 25492
rect 30196 25440 30248 25492
rect 11980 25304 12032 25356
rect 14188 25372 14240 25424
rect 16856 25372 16908 25424
rect 9496 25279 9548 25288
rect 9496 25245 9505 25279
rect 9505 25245 9539 25279
rect 9539 25245 9548 25279
rect 9496 25236 9548 25245
rect 10692 25236 10744 25288
rect 10968 25236 11020 25288
rect 13268 25279 13320 25288
rect 1768 25143 1820 25152
rect 1768 25109 1777 25143
rect 1777 25109 1811 25143
rect 1811 25109 1820 25143
rect 1768 25100 1820 25109
rect 6000 25100 6052 25152
rect 9864 25100 9916 25152
rect 11980 25100 12032 25152
rect 12992 25100 13044 25152
rect 13268 25245 13277 25279
rect 13277 25245 13311 25279
rect 13311 25245 13320 25279
rect 13268 25236 13320 25245
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 14188 25168 14240 25220
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 14464 25168 14516 25177
rect 16580 25168 16632 25220
rect 16856 25211 16908 25220
rect 16856 25177 16865 25211
rect 16865 25177 16899 25211
rect 16899 25177 16908 25211
rect 16856 25168 16908 25177
rect 15752 25100 15804 25152
rect 16028 25100 16080 25152
rect 17040 25168 17092 25220
rect 25688 25372 25740 25424
rect 37648 25372 37700 25424
rect 20260 25236 20312 25288
rect 20628 25279 20680 25288
rect 20628 25245 20637 25279
rect 20637 25245 20671 25279
rect 20671 25245 20680 25279
rect 20628 25236 20680 25245
rect 24216 25236 24268 25288
rect 24768 25236 24820 25288
rect 20536 25168 20588 25220
rect 21456 25211 21508 25220
rect 21456 25177 21465 25211
rect 21465 25177 21499 25211
rect 21499 25177 21508 25211
rect 22008 25211 22060 25220
rect 21456 25168 21508 25177
rect 22008 25177 22017 25211
rect 22017 25177 22051 25211
rect 22051 25177 22060 25211
rect 22008 25168 22060 25177
rect 23572 25168 23624 25220
rect 24584 25168 24636 25220
rect 18328 25100 18380 25152
rect 18512 25143 18564 25152
rect 18512 25109 18521 25143
rect 18521 25109 18555 25143
rect 18555 25109 18564 25143
rect 18512 25100 18564 25109
rect 21180 25100 21232 25152
rect 25504 25211 25556 25220
rect 25504 25177 25513 25211
rect 25513 25177 25547 25211
rect 25547 25177 25556 25211
rect 25504 25168 25556 25177
rect 26700 25168 26752 25220
rect 26516 25100 26568 25152
rect 27252 25304 27304 25356
rect 27620 25347 27672 25356
rect 27620 25313 27629 25347
rect 27629 25313 27663 25347
rect 27663 25313 27672 25347
rect 27620 25304 27672 25313
rect 28540 25304 28592 25356
rect 30104 25304 30156 25356
rect 31760 25347 31812 25356
rect 31760 25313 31769 25347
rect 31769 25313 31803 25347
rect 31803 25313 31812 25347
rect 31760 25304 31812 25313
rect 33692 25347 33744 25356
rect 33692 25313 33701 25347
rect 33701 25313 33735 25347
rect 33735 25313 33744 25347
rect 33692 25304 33744 25313
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 27804 25168 27856 25220
rect 28816 25168 28868 25220
rect 29828 25211 29880 25220
rect 29828 25177 29837 25211
rect 29837 25177 29871 25211
rect 29871 25177 29880 25211
rect 29828 25168 29880 25177
rect 29920 25211 29972 25220
rect 29920 25177 29929 25211
rect 29929 25177 29963 25211
rect 29963 25177 29972 25211
rect 29920 25168 29972 25177
rect 31484 25211 31536 25220
rect 28080 25100 28132 25152
rect 28448 25100 28500 25152
rect 31484 25177 31493 25211
rect 31493 25177 31527 25211
rect 31527 25177 31536 25211
rect 31484 25168 31536 25177
rect 31576 25211 31628 25220
rect 31576 25177 31585 25211
rect 31585 25177 31619 25211
rect 31619 25177 31628 25211
rect 33784 25211 33836 25220
rect 31576 25168 31628 25177
rect 33784 25177 33793 25211
rect 33793 25177 33827 25211
rect 33827 25177 33836 25211
rect 33784 25168 33836 25177
rect 30932 25100 30984 25152
rect 33416 25100 33468 25152
rect 33968 25100 34020 25152
rect 34428 25168 34480 25220
rect 38660 25168 38712 25220
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7288 24896 7340 24948
rect 10692 24896 10744 24948
rect 9680 24828 9732 24880
rect 12164 24871 12216 24880
rect 1768 24803 1820 24812
rect 1768 24769 1777 24803
rect 1777 24769 1811 24803
rect 1811 24769 1820 24803
rect 1768 24760 1820 24769
rect 9404 24735 9456 24744
rect 9404 24701 9413 24735
rect 9413 24701 9447 24735
rect 9447 24701 9456 24735
rect 9404 24692 9456 24701
rect 9588 24692 9640 24744
rect 8208 24624 8260 24676
rect 12164 24837 12173 24871
rect 12173 24837 12207 24871
rect 12207 24837 12216 24871
rect 12164 24828 12216 24837
rect 12716 24803 12768 24812
rect 10600 24692 10652 24744
rect 12716 24769 12725 24803
rect 12725 24769 12759 24803
rect 12759 24769 12768 24803
rect 12716 24760 12768 24769
rect 16488 24896 16540 24948
rect 13452 24760 13504 24812
rect 14004 24760 14056 24812
rect 13268 24692 13320 24744
rect 15108 24624 15160 24676
rect 15384 24760 15436 24812
rect 16672 24760 16724 24812
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 19156 24803 19208 24812
rect 16764 24692 16816 24744
rect 17132 24692 17184 24744
rect 17316 24735 17368 24744
rect 17316 24701 17325 24735
rect 17325 24701 17359 24735
rect 17359 24701 17368 24735
rect 17316 24692 17368 24701
rect 17592 24692 17644 24744
rect 18328 24692 18380 24744
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 20904 24871 20956 24880
rect 20904 24837 20913 24871
rect 20913 24837 20947 24871
rect 20947 24837 20956 24871
rect 26700 24896 26752 24948
rect 27896 24896 27948 24948
rect 20904 24828 20956 24837
rect 24216 24871 24268 24880
rect 24216 24837 24225 24871
rect 24225 24837 24259 24871
rect 24259 24837 24268 24871
rect 24216 24828 24268 24837
rect 23940 24760 23992 24812
rect 19708 24624 19760 24676
rect 20720 24692 20772 24744
rect 22836 24735 22888 24744
rect 22836 24701 22845 24735
rect 22845 24701 22879 24735
rect 22879 24701 22888 24735
rect 22836 24692 22888 24701
rect 23020 24692 23072 24744
rect 24492 24692 24544 24744
rect 25412 24760 25464 24812
rect 25688 24760 25740 24812
rect 25964 24692 26016 24744
rect 26332 24803 26384 24812
rect 26332 24769 26341 24803
rect 26341 24769 26375 24803
rect 26375 24769 26384 24803
rect 27436 24828 27488 24880
rect 29920 24828 29972 24880
rect 30288 24871 30340 24880
rect 30288 24837 30297 24871
rect 30297 24837 30331 24871
rect 30331 24837 30340 24871
rect 30288 24828 30340 24837
rect 26332 24760 26384 24769
rect 26700 24692 26752 24744
rect 1860 24556 1912 24608
rect 9588 24556 9640 24608
rect 13268 24556 13320 24608
rect 13360 24556 13412 24608
rect 14648 24599 14700 24608
rect 14648 24565 14657 24599
rect 14657 24565 14691 24599
rect 14691 24565 14700 24599
rect 14648 24556 14700 24565
rect 15292 24599 15344 24608
rect 15292 24565 15301 24599
rect 15301 24565 15335 24599
rect 15335 24565 15344 24599
rect 15292 24556 15344 24565
rect 15936 24556 15988 24608
rect 23848 24624 23900 24676
rect 24308 24624 24360 24676
rect 27988 24692 28040 24744
rect 29828 24760 29880 24812
rect 32864 24760 32916 24812
rect 33784 24760 33836 24812
rect 35348 24760 35400 24812
rect 29000 24735 29052 24744
rect 29000 24701 29009 24735
rect 29009 24701 29043 24735
rect 29043 24701 29052 24735
rect 29000 24692 29052 24701
rect 30012 24692 30064 24744
rect 30196 24735 30248 24744
rect 30196 24701 30205 24735
rect 30205 24701 30239 24735
rect 30239 24701 30248 24735
rect 30196 24692 30248 24701
rect 32036 24692 32088 24744
rect 29184 24624 29236 24676
rect 23480 24556 23532 24608
rect 26056 24556 26108 24608
rect 27620 24556 27672 24608
rect 29092 24556 29144 24608
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9864 24352 9916 24404
rect 10600 24352 10652 24404
rect 11428 24352 11480 24404
rect 11980 24352 12032 24404
rect 13268 24352 13320 24404
rect 15016 24352 15068 24404
rect 9404 24259 9456 24268
rect 9404 24225 9413 24259
rect 9413 24225 9447 24259
rect 9447 24225 9456 24259
rect 9404 24216 9456 24225
rect 12164 24284 12216 24336
rect 14556 24284 14608 24336
rect 11244 24216 11296 24268
rect 12348 24216 12400 24268
rect 12532 24259 12584 24268
rect 12532 24225 12541 24259
rect 12541 24225 12575 24259
rect 12575 24225 12584 24259
rect 12532 24216 12584 24225
rect 13268 24216 13320 24268
rect 20260 24352 20312 24404
rect 24216 24352 24268 24404
rect 24768 24352 24820 24404
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 1860 24148 1912 24200
rect 13728 24148 13780 24200
rect 19892 24284 19944 24336
rect 15936 24259 15988 24268
rect 15936 24225 15945 24259
rect 15945 24225 15979 24259
rect 15979 24225 15988 24259
rect 15936 24216 15988 24225
rect 16856 24216 16908 24268
rect 17776 24216 17828 24268
rect 18236 24216 18288 24268
rect 24124 24284 24176 24336
rect 24860 24284 24912 24336
rect 20536 24216 20588 24268
rect 21272 24216 21324 24268
rect 25504 24352 25556 24404
rect 26516 24352 26568 24404
rect 37464 24352 37516 24404
rect 25688 24284 25740 24336
rect 26424 24284 26476 24336
rect 19708 24148 19760 24200
rect 20444 24148 20496 24200
rect 25504 24216 25556 24268
rect 25320 24148 25372 24200
rect 26424 24148 26476 24200
rect 26608 24327 26660 24336
rect 26608 24293 26617 24327
rect 26617 24293 26651 24327
rect 26651 24293 26660 24327
rect 26608 24284 26660 24293
rect 27988 24284 28040 24336
rect 30564 24284 30616 24336
rect 31760 24284 31812 24336
rect 28448 24259 28500 24268
rect 28448 24225 28457 24259
rect 28457 24225 28491 24259
rect 28491 24225 28500 24259
rect 28448 24216 28500 24225
rect 30012 24259 30064 24268
rect 30012 24225 30021 24259
rect 30021 24225 30055 24259
rect 30055 24225 30064 24259
rect 30012 24216 30064 24225
rect 31024 24259 31076 24268
rect 31024 24225 31033 24259
rect 31033 24225 31067 24259
rect 31067 24225 31076 24259
rect 31024 24216 31076 24225
rect 31300 24216 31352 24268
rect 32312 24216 32364 24268
rect 34612 24216 34664 24268
rect 37740 24216 37792 24268
rect 38292 24191 38344 24200
rect 11060 24080 11112 24132
rect 11244 24080 11296 24132
rect 12072 24123 12124 24132
rect 12072 24089 12081 24123
rect 12081 24089 12115 24123
rect 12115 24089 12124 24123
rect 12072 24080 12124 24089
rect 15108 24080 15160 24132
rect 5540 24012 5592 24064
rect 10600 24012 10652 24064
rect 13820 24012 13872 24064
rect 15844 24012 15896 24064
rect 16028 24123 16080 24132
rect 16028 24089 16037 24123
rect 16037 24089 16071 24123
rect 16071 24089 16080 24123
rect 16028 24080 16080 24089
rect 17040 24080 17092 24132
rect 18236 24080 18288 24132
rect 18420 24080 18472 24132
rect 19616 24080 19668 24132
rect 18512 24012 18564 24064
rect 18880 24012 18932 24064
rect 20720 24080 20772 24132
rect 21180 24123 21232 24132
rect 21180 24089 21189 24123
rect 21189 24089 21223 24123
rect 21223 24089 21232 24123
rect 23020 24123 23072 24132
rect 21180 24080 21232 24089
rect 23020 24089 23029 24123
rect 23029 24089 23063 24123
rect 23063 24089 23072 24123
rect 23020 24080 23072 24089
rect 23848 24080 23900 24132
rect 24124 24080 24176 24132
rect 27988 24080 28040 24132
rect 25412 24012 25464 24064
rect 27436 24012 27488 24064
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 32220 24123 32272 24132
rect 32220 24089 32229 24123
rect 32229 24089 32263 24123
rect 32263 24089 32272 24123
rect 32220 24080 32272 24089
rect 34060 24012 34112 24064
rect 38108 24055 38160 24064
rect 38108 24021 38117 24055
rect 38117 24021 38151 24055
rect 38151 24021 38160 24055
rect 38108 24012 38160 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1676 23808 1728 23860
rect 2412 23851 2464 23860
rect 2412 23817 2421 23851
rect 2421 23817 2455 23851
rect 2455 23817 2464 23851
rect 2412 23808 2464 23817
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 2596 23715 2648 23724
rect 2596 23681 2605 23715
rect 2605 23681 2639 23715
rect 2639 23681 2648 23715
rect 2596 23672 2648 23681
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 14464 23808 14516 23860
rect 18236 23851 18288 23860
rect 11060 23783 11112 23792
rect 11060 23749 11069 23783
rect 11069 23749 11103 23783
rect 11103 23749 11112 23783
rect 13820 23783 13872 23792
rect 11060 23740 11112 23749
rect 6460 23604 6512 23656
rect 9956 23604 10008 23656
rect 11612 23672 11664 23724
rect 10784 23536 10836 23588
rect 13820 23749 13829 23783
rect 13829 23749 13863 23783
rect 13863 23749 13872 23783
rect 13820 23740 13872 23749
rect 14648 23740 14700 23792
rect 17776 23740 17828 23792
rect 18236 23817 18245 23851
rect 18245 23817 18279 23851
rect 18279 23817 18288 23851
rect 18236 23808 18288 23817
rect 19892 23808 19944 23860
rect 23296 23808 23348 23860
rect 28448 23808 28500 23860
rect 30288 23808 30340 23860
rect 32220 23808 32272 23860
rect 34796 23808 34848 23860
rect 38016 23808 38068 23860
rect 18880 23783 18932 23792
rect 18880 23749 18889 23783
rect 18889 23749 18923 23783
rect 18923 23749 18932 23783
rect 18880 23740 18932 23749
rect 19524 23740 19576 23792
rect 20720 23740 20772 23792
rect 21916 23740 21968 23792
rect 22376 23740 22428 23792
rect 24308 23783 24360 23792
rect 24308 23749 24317 23783
rect 24317 23749 24351 23783
rect 24351 23749 24360 23783
rect 24308 23740 24360 23749
rect 28908 23783 28960 23792
rect 28908 23749 28917 23783
rect 28917 23749 28951 23783
rect 28951 23749 28960 23783
rect 28908 23740 28960 23749
rect 30564 23740 30616 23792
rect 31484 23740 31536 23792
rect 15936 23604 15988 23656
rect 16488 23536 16540 23588
rect 12072 23468 12124 23520
rect 12900 23468 12952 23520
rect 12992 23468 13044 23520
rect 17040 23672 17092 23724
rect 17408 23672 17460 23724
rect 18420 23672 18472 23724
rect 24216 23715 24268 23724
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 20536 23604 20588 23656
rect 20720 23647 20772 23656
rect 20720 23613 20729 23647
rect 20729 23613 20763 23647
rect 20763 23613 20772 23647
rect 20720 23604 20772 23613
rect 21732 23604 21784 23656
rect 23204 23604 23256 23656
rect 25228 23672 25280 23724
rect 25688 23672 25740 23724
rect 24952 23604 25004 23656
rect 25596 23604 25648 23656
rect 22008 23536 22060 23588
rect 29828 23672 29880 23724
rect 30288 23715 30340 23724
rect 30288 23681 30297 23715
rect 30297 23681 30331 23715
rect 30331 23681 30340 23715
rect 30288 23672 30340 23681
rect 26884 23604 26936 23656
rect 27528 23647 27580 23656
rect 27528 23613 27537 23647
rect 27537 23613 27571 23647
rect 27571 23613 27580 23647
rect 27528 23604 27580 23613
rect 28172 23604 28224 23656
rect 28816 23647 28868 23656
rect 28816 23613 28825 23647
rect 28825 23613 28859 23647
rect 28859 23613 28868 23647
rect 28816 23604 28868 23613
rect 29092 23647 29144 23656
rect 29092 23613 29101 23647
rect 29101 23613 29135 23647
rect 29135 23613 29144 23647
rect 29092 23604 29144 23613
rect 30748 23536 30800 23588
rect 31852 23672 31904 23724
rect 33876 23715 33928 23724
rect 33876 23681 33885 23715
rect 33885 23681 33919 23715
rect 33919 23681 33928 23715
rect 33876 23672 33928 23681
rect 37924 23672 37976 23724
rect 34520 23604 34572 23656
rect 32864 23536 32916 23588
rect 16856 23468 16908 23520
rect 17500 23468 17552 23520
rect 23664 23511 23716 23520
rect 23664 23477 23673 23511
rect 23673 23477 23707 23511
rect 23707 23477 23716 23511
rect 23664 23468 23716 23477
rect 24952 23511 25004 23520
rect 24952 23477 24961 23511
rect 24961 23477 24995 23511
rect 24995 23477 25004 23511
rect 24952 23468 25004 23477
rect 25228 23468 25280 23520
rect 27436 23468 27488 23520
rect 30472 23468 30524 23520
rect 31024 23511 31076 23520
rect 31024 23477 31033 23511
rect 31033 23477 31067 23511
rect 31067 23477 31076 23511
rect 31024 23468 31076 23477
rect 31852 23468 31904 23520
rect 32680 23468 32732 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4068 23264 4120 23316
rect 10140 23264 10192 23316
rect 11244 23264 11296 23316
rect 13912 23264 13964 23316
rect 15200 23264 15252 23316
rect 15660 23264 15712 23316
rect 22468 23264 22520 23316
rect 23296 23264 23348 23316
rect 23940 23307 23992 23316
rect 23940 23273 23949 23307
rect 23949 23273 23983 23307
rect 23983 23273 23992 23307
rect 23940 23264 23992 23273
rect 25504 23264 25556 23316
rect 27804 23307 27856 23316
rect 10784 23196 10836 23248
rect 14096 23196 14148 23248
rect 24032 23196 24084 23248
rect 14648 23171 14700 23180
rect 14648 23137 14657 23171
rect 14657 23137 14691 23171
rect 14691 23137 14700 23171
rect 14648 23128 14700 23137
rect 15936 23128 15988 23180
rect 17132 23128 17184 23180
rect 22928 23171 22980 23180
rect 22928 23137 22937 23171
rect 22937 23137 22971 23171
rect 22971 23137 22980 23171
rect 22928 23128 22980 23137
rect 25780 23196 25832 23248
rect 27804 23273 27813 23307
rect 27813 23273 27847 23307
rect 27847 23273 27856 23307
rect 27804 23264 27856 23273
rect 28908 23264 28960 23316
rect 31576 23264 31628 23316
rect 31668 23264 31720 23316
rect 33048 23264 33100 23316
rect 26240 23128 26292 23180
rect 33232 23196 33284 23248
rect 5540 23060 5592 23112
rect 7840 23103 7892 23112
rect 7840 23069 7849 23103
rect 7849 23069 7883 23103
rect 7883 23069 7892 23103
rect 7840 23060 7892 23069
rect 8852 23060 8904 23112
rect 940 22992 992 23044
rect 10784 23060 10836 23112
rect 11796 23060 11848 23112
rect 14096 23060 14148 23112
rect 20260 23060 20312 23112
rect 20444 23060 20496 23112
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 11704 22992 11756 23044
rect 7748 22924 7800 22976
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 15936 23035 15988 23044
rect 15936 23001 15945 23035
rect 15945 23001 15979 23035
rect 15979 23001 15988 23035
rect 15936 22992 15988 23001
rect 17408 23035 17460 23044
rect 16580 22924 16632 22976
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 17500 23035 17552 23044
rect 17500 23001 17509 23035
rect 17509 23001 17543 23035
rect 17543 23001 17552 23035
rect 19524 23035 19576 23044
rect 17500 22992 17552 23001
rect 19524 23001 19533 23035
rect 19533 23001 19567 23035
rect 19567 23001 19576 23035
rect 19524 22992 19576 23001
rect 22376 23035 22428 23044
rect 22376 23001 22385 23035
rect 22385 23001 22419 23035
rect 22419 23001 22428 23035
rect 22376 22992 22428 23001
rect 23664 23060 23716 23112
rect 24492 23060 24544 23112
rect 26148 23103 26200 23112
rect 26148 23069 26157 23103
rect 26157 23069 26191 23103
rect 26191 23069 26200 23103
rect 26148 23060 26200 23069
rect 27068 23103 27120 23112
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 33784 23128 33836 23180
rect 29092 23060 29144 23112
rect 29368 23060 29420 23112
rect 31208 23060 31260 23112
rect 35348 23060 35400 23112
rect 24768 23035 24820 23044
rect 24768 23001 24777 23035
rect 24777 23001 24811 23035
rect 24811 23001 24820 23035
rect 24768 22992 24820 23001
rect 21916 22924 21968 22976
rect 25412 22924 25464 22976
rect 26056 22992 26108 23044
rect 26700 22992 26752 23044
rect 26240 22967 26292 22976
rect 26240 22933 26249 22967
rect 26249 22933 26283 22967
rect 26283 22933 26292 22967
rect 26240 22924 26292 22933
rect 27344 22924 27396 22976
rect 29828 22992 29880 23044
rect 28540 22924 28592 22976
rect 30932 22992 30984 23044
rect 32036 23035 32088 23044
rect 32036 23001 32045 23035
rect 32045 23001 32079 23035
rect 32079 23001 32088 23035
rect 32036 22992 32088 23001
rect 33048 23035 33100 23044
rect 33048 23001 33057 23035
rect 33057 23001 33091 23035
rect 33091 23001 33100 23035
rect 33048 22992 33100 23001
rect 33968 22924 34020 22976
rect 38016 22924 38068 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 7748 22695 7800 22704
rect 7748 22661 7757 22695
rect 7757 22661 7791 22695
rect 7791 22661 7800 22695
rect 7748 22652 7800 22661
rect 10232 22695 10284 22704
rect 10232 22661 10241 22695
rect 10241 22661 10275 22695
rect 10275 22661 10284 22695
rect 10232 22652 10284 22661
rect 10600 22652 10652 22704
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 8392 22516 8444 22568
rect 9404 22559 9456 22568
rect 9404 22525 9413 22559
rect 9413 22525 9447 22559
rect 9447 22525 9456 22559
rect 9404 22516 9456 22525
rect 10140 22559 10192 22568
rect 10140 22525 10149 22559
rect 10149 22525 10183 22559
rect 10183 22525 10192 22559
rect 10140 22516 10192 22525
rect 11244 22652 11296 22704
rect 13728 22720 13780 22772
rect 13360 22695 13412 22704
rect 13360 22661 13369 22695
rect 13369 22661 13403 22695
rect 13403 22661 13412 22695
rect 13360 22652 13412 22661
rect 12992 22584 13044 22636
rect 15108 22695 15160 22704
rect 15108 22661 15117 22695
rect 15117 22661 15151 22695
rect 15151 22661 15160 22695
rect 15108 22652 15160 22661
rect 15660 22652 15712 22704
rect 19432 22720 19484 22772
rect 19984 22720 20036 22772
rect 24492 22720 24544 22772
rect 29276 22720 29328 22772
rect 29644 22720 29696 22772
rect 29920 22720 29972 22772
rect 31668 22720 31720 22772
rect 20628 22652 20680 22704
rect 23480 22652 23532 22704
rect 24952 22652 25004 22704
rect 25136 22652 25188 22704
rect 27344 22695 27396 22704
rect 17224 22627 17276 22636
rect 17224 22593 17233 22627
rect 17233 22593 17267 22627
rect 17267 22593 17276 22627
rect 17224 22584 17276 22593
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 19524 22627 19576 22636
rect 19524 22593 19533 22627
rect 19533 22593 19567 22627
rect 19567 22593 19576 22627
rect 19524 22584 19576 22593
rect 21364 22584 21416 22636
rect 25504 22584 25556 22636
rect 27344 22661 27353 22695
rect 27353 22661 27387 22695
rect 27387 22661 27396 22695
rect 27344 22652 27396 22661
rect 28540 22695 28592 22704
rect 28540 22661 28549 22695
rect 28549 22661 28583 22695
rect 28583 22661 28592 22695
rect 28540 22652 28592 22661
rect 29552 22652 29604 22704
rect 29828 22652 29880 22704
rect 31024 22652 31076 22704
rect 32220 22652 32272 22704
rect 37924 22720 37976 22772
rect 38108 22652 38160 22704
rect 15200 22516 15252 22568
rect 21272 22516 21324 22568
rect 22376 22559 22428 22568
rect 22376 22525 22385 22559
rect 22385 22525 22419 22559
rect 22419 22525 22428 22559
rect 22376 22516 22428 22525
rect 22560 22516 22612 22568
rect 25044 22516 25096 22568
rect 27252 22559 27304 22568
rect 7840 22448 7892 22500
rect 21180 22448 21232 22500
rect 5540 22380 5592 22432
rect 10324 22380 10376 22432
rect 12164 22380 12216 22432
rect 17868 22380 17920 22432
rect 18144 22380 18196 22432
rect 19064 22380 19116 22432
rect 22100 22448 22152 22500
rect 27252 22525 27261 22559
rect 27261 22525 27295 22559
rect 27295 22525 27304 22559
rect 27252 22516 27304 22525
rect 27436 22516 27488 22568
rect 25136 22380 25188 22432
rect 26332 22423 26384 22432
rect 26332 22389 26341 22423
rect 26341 22389 26375 22423
rect 26375 22389 26384 22423
rect 26332 22380 26384 22389
rect 29920 22448 29972 22500
rect 30748 22516 30800 22568
rect 31484 22516 31536 22568
rect 35348 22584 35400 22636
rect 38016 22627 38068 22636
rect 38016 22593 38025 22627
rect 38025 22593 38059 22627
rect 38059 22593 38068 22627
rect 38016 22584 38068 22593
rect 31668 22516 31720 22568
rect 34612 22516 34664 22568
rect 30380 22448 30432 22500
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 30748 22380 30800 22432
rect 30932 22380 30984 22432
rect 32312 22380 32364 22432
rect 33140 22380 33192 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8392 22219 8444 22228
rect 8392 22185 8401 22219
rect 8401 22185 8435 22219
rect 8435 22185 8444 22219
rect 8392 22176 8444 22185
rect 17408 22176 17460 22228
rect 18236 22176 18288 22228
rect 18328 22176 18380 22228
rect 20260 22176 20312 22228
rect 1952 22108 2004 22160
rect 8208 22108 8260 22160
rect 11704 22108 11756 22160
rect 12348 22108 12400 22160
rect 1768 21879 1820 21888
rect 1768 21845 1777 21879
rect 1777 21845 1811 21879
rect 1811 21845 1820 21879
rect 1768 21836 1820 21845
rect 9956 22040 10008 22092
rect 10140 22083 10192 22092
rect 10140 22049 10149 22083
rect 10149 22049 10183 22083
rect 10183 22049 10192 22083
rect 12900 22108 12952 22160
rect 16948 22108 17000 22160
rect 10140 22040 10192 22049
rect 13820 22040 13872 22092
rect 14464 22040 14516 22092
rect 15200 22040 15252 22092
rect 5540 21972 5592 22024
rect 8484 21972 8536 22024
rect 12992 21972 13044 22024
rect 13452 21972 13504 22024
rect 10140 21904 10192 21956
rect 11152 21947 11204 21956
rect 11152 21913 11161 21947
rect 11161 21913 11195 21947
rect 11195 21913 11204 21947
rect 11152 21904 11204 21913
rect 11704 21947 11756 21956
rect 11704 21913 11713 21947
rect 11713 21913 11747 21947
rect 11747 21913 11756 21947
rect 11704 21904 11756 21913
rect 11796 21947 11848 21956
rect 11796 21913 11805 21947
rect 11805 21913 11839 21947
rect 11839 21913 11848 21947
rect 11796 21904 11848 21913
rect 13084 21904 13136 21956
rect 16304 21947 16356 21956
rect 10324 21836 10376 21888
rect 13820 21836 13872 21888
rect 16304 21913 16313 21947
rect 16313 21913 16347 21947
rect 16347 21913 16356 21947
rect 16304 21904 16356 21913
rect 16764 21904 16816 21956
rect 17316 22040 17368 22092
rect 19892 22040 19944 22092
rect 21180 22108 21232 22160
rect 23480 22108 23532 22160
rect 23756 22176 23808 22228
rect 33140 22176 33192 22228
rect 27252 22108 27304 22160
rect 23572 22083 23624 22092
rect 23572 22049 23581 22083
rect 23581 22049 23615 22083
rect 23615 22049 23624 22083
rect 23572 22040 23624 22049
rect 25964 22083 26016 22092
rect 25964 22049 25973 22083
rect 25973 22049 26007 22083
rect 26007 22049 26016 22083
rect 25964 22040 26016 22049
rect 26056 22040 26108 22092
rect 29644 22108 29696 22160
rect 32312 22108 32364 22160
rect 19432 21972 19484 22024
rect 22744 21972 22796 22024
rect 23848 21972 23900 22024
rect 28448 22040 28500 22092
rect 30380 22040 30432 22092
rect 33784 22083 33836 22092
rect 33784 22049 33793 22083
rect 33793 22049 33827 22083
rect 33827 22049 33836 22083
rect 33784 22040 33836 22049
rect 34520 22040 34572 22092
rect 17408 21904 17460 21956
rect 17868 21947 17920 21956
rect 17868 21913 17877 21947
rect 17877 21913 17911 21947
rect 17911 21913 17920 21947
rect 17868 21904 17920 21913
rect 21272 21904 21324 21956
rect 25136 21947 25188 21956
rect 25136 21913 25145 21947
rect 25145 21913 25179 21947
rect 25179 21913 25188 21947
rect 25136 21904 25188 21913
rect 25228 21947 25280 21956
rect 25228 21913 25237 21947
rect 25237 21913 25271 21947
rect 25271 21913 25280 21947
rect 25228 21904 25280 21913
rect 25504 21904 25556 21956
rect 26332 21904 26384 21956
rect 26884 21947 26936 21956
rect 26884 21913 26893 21947
rect 26893 21913 26927 21947
rect 26927 21913 26936 21947
rect 26884 21904 26936 21913
rect 27528 21904 27580 21956
rect 31760 21972 31812 22024
rect 32220 21972 32272 22024
rect 32772 21972 32824 22024
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 28908 21904 28960 21956
rect 29644 21904 29696 21956
rect 30932 21947 30984 21956
rect 30932 21913 30941 21947
rect 30941 21913 30975 21947
rect 30975 21913 30984 21947
rect 30932 21904 30984 21913
rect 22284 21836 22336 21888
rect 22928 21836 22980 21888
rect 27988 21836 28040 21888
rect 30012 21836 30064 21888
rect 32496 21904 32548 21956
rect 32404 21879 32456 21888
rect 32404 21845 32413 21879
rect 32413 21845 32447 21879
rect 32447 21845 32456 21879
rect 32404 21836 32456 21845
rect 36360 21972 36412 22024
rect 38292 22015 38344 22024
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 38016 21904 38068 21956
rect 33876 21836 33928 21888
rect 36544 21836 36596 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 10232 21632 10284 21684
rect 11704 21632 11756 21684
rect 11796 21632 11848 21684
rect 16304 21632 16356 21684
rect 16396 21632 16448 21684
rect 19800 21632 19852 21684
rect 19984 21632 20036 21684
rect 22192 21632 22244 21684
rect 22744 21632 22796 21684
rect 27068 21632 27120 21684
rect 27804 21675 27856 21684
rect 27804 21641 27813 21675
rect 27813 21641 27847 21675
rect 27847 21641 27856 21675
rect 27804 21632 27856 21641
rect 10692 21564 10744 21616
rect 11152 21564 11204 21616
rect 12716 21564 12768 21616
rect 14648 21564 14700 21616
rect 16672 21564 16724 21616
rect 17224 21607 17276 21616
rect 17224 21573 17233 21607
rect 17233 21573 17267 21607
rect 17267 21573 17276 21607
rect 17224 21564 17276 21573
rect 19340 21564 19392 21616
rect 10324 21539 10376 21548
rect 10324 21505 10333 21539
rect 10333 21505 10367 21539
rect 10367 21505 10376 21539
rect 10324 21496 10376 21505
rect 10508 21496 10560 21548
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 12532 21496 12584 21548
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 18604 21496 18656 21548
rect 19248 21496 19300 21548
rect 19616 21539 19668 21548
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 21272 21564 21324 21616
rect 13084 21428 13136 21480
rect 10784 21360 10836 21412
rect 11244 21360 11296 21412
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 12072 21360 12124 21412
rect 14464 21428 14516 21480
rect 15200 21428 15252 21480
rect 15844 21428 15896 21480
rect 17408 21428 17460 21480
rect 20536 21496 20588 21548
rect 20904 21539 20956 21548
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 21180 21496 21232 21548
rect 21824 21496 21876 21548
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 23572 21564 23624 21616
rect 23940 21564 23992 21616
rect 25504 21564 25556 21616
rect 28908 21564 28960 21616
rect 30104 21564 30156 21616
rect 32404 21564 32456 21616
rect 27620 21539 27672 21548
rect 27620 21505 27629 21539
rect 27629 21505 27663 21539
rect 27663 21505 27672 21539
rect 27620 21496 27672 21505
rect 29552 21539 29604 21548
rect 29552 21505 29561 21539
rect 29561 21505 29595 21539
rect 29595 21505 29604 21539
rect 29552 21496 29604 21505
rect 19892 21428 19944 21480
rect 23756 21428 23808 21480
rect 24124 21471 24176 21480
rect 24124 21437 24133 21471
rect 24133 21437 24167 21471
rect 24167 21437 24176 21471
rect 25136 21471 25188 21480
rect 24124 21428 24176 21437
rect 25136 21437 25145 21471
rect 25145 21437 25179 21471
rect 25179 21437 25188 21471
rect 25136 21428 25188 21437
rect 25964 21471 26016 21480
rect 25964 21437 25973 21471
rect 25973 21437 26007 21471
rect 26007 21437 26016 21471
rect 25964 21428 26016 21437
rect 28264 21428 28316 21480
rect 28632 21428 28684 21480
rect 30564 21496 30616 21548
rect 17132 21292 17184 21344
rect 18880 21292 18932 21344
rect 19432 21292 19484 21344
rect 19800 21292 19852 21344
rect 20904 21292 20956 21344
rect 22192 21292 22244 21344
rect 22284 21292 22336 21344
rect 24860 21360 24912 21412
rect 27436 21292 27488 21344
rect 28632 21292 28684 21344
rect 29644 21360 29696 21412
rect 31852 21496 31904 21548
rect 32220 21496 32272 21548
rect 32588 21496 32640 21548
rect 32956 21539 33008 21548
rect 32956 21505 32965 21539
rect 32965 21505 32999 21539
rect 32999 21505 33008 21539
rect 32956 21496 33008 21505
rect 33600 21539 33652 21548
rect 33600 21505 33609 21539
rect 33609 21505 33643 21539
rect 33643 21505 33652 21539
rect 33600 21496 33652 21505
rect 36360 21496 36412 21548
rect 29920 21360 29972 21412
rect 30380 21292 30432 21344
rect 32496 21292 32548 21344
rect 33416 21292 33468 21344
rect 34336 21335 34388 21344
rect 34336 21301 34345 21335
rect 34345 21301 34379 21335
rect 34379 21301 34388 21335
rect 34336 21292 34388 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 10140 21088 10192 21140
rect 15384 21088 15436 21140
rect 12532 21020 12584 21072
rect 12900 21020 12952 21072
rect 13452 21020 13504 21072
rect 17040 21088 17092 21140
rect 17132 21088 17184 21140
rect 23940 21131 23992 21140
rect 23940 21097 23949 21131
rect 23949 21097 23983 21131
rect 23983 21097 23992 21131
rect 23940 21088 23992 21097
rect 24768 21088 24820 21140
rect 24952 21088 25004 21140
rect 26148 21088 26200 21140
rect 27620 21088 27672 21140
rect 37280 21088 37332 21140
rect 37924 21088 37976 21140
rect 6828 20884 6880 20936
rect 13636 20952 13688 21004
rect 13452 20884 13504 20936
rect 10692 20816 10744 20868
rect 1768 20791 1820 20800
rect 1768 20757 1777 20791
rect 1777 20757 1811 20791
rect 1811 20757 1820 20791
rect 1768 20748 1820 20757
rect 4068 20748 4120 20800
rect 10508 20748 10560 20800
rect 11152 20748 11204 20800
rect 18052 20952 18104 21004
rect 14096 20748 14148 20800
rect 14740 20884 14792 20936
rect 15936 20859 15988 20868
rect 15936 20825 15945 20859
rect 15945 20825 15979 20859
rect 15979 20825 15988 20859
rect 15936 20816 15988 20825
rect 17040 20748 17092 20800
rect 17500 20859 17552 20868
rect 17500 20825 17509 20859
rect 17509 20825 17543 20859
rect 17543 20825 17552 20859
rect 17500 20816 17552 20825
rect 17684 20816 17736 20868
rect 21824 20952 21876 21004
rect 24124 21020 24176 21072
rect 27528 21020 27580 21072
rect 24308 20952 24360 21004
rect 25136 20952 25188 21004
rect 26240 20952 26292 21004
rect 27988 20995 28040 21004
rect 27988 20961 27997 20995
rect 27997 20961 28031 20995
rect 28031 20961 28040 20995
rect 27988 20952 28040 20961
rect 28264 20995 28316 21004
rect 28264 20961 28273 20995
rect 28273 20961 28307 20995
rect 28307 20961 28316 20995
rect 28264 20952 28316 20961
rect 30196 20952 30248 21004
rect 21548 20884 21600 20936
rect 23940 20884 23992 20936
rect 24952 20884 25004 20936
rect 29184 20884 29236 20936
rect 19892 20859 19944 20868
rect 17592 20748 17644 20800
rect 19892 20825 19901 20859
rect 19901 20825 19935 20859
rect 19935 20825 19944 20859
rect 19892 20816 19944 20825
rect 19984 20859 20036 20868
rect 19984 20825 19993 20859
rect 19993 20825 20027 20859
rect 20027 20825 20036 20859
rect 19984 20816 20036 20825
rect 20812 20816 20864 20868
rect 21088 20816 21140 20868
rect 21916 20816 21968 20868
rect 22284 20859 22336 20868
rect 22284 20825 22293 20859
rect 22293 20825 22327 20859
rect 22327 20825 22336 20859
rect 22284 20816 22336 20825
rect 23296 20816 23348 20868
rect 18604 20748 18656 20800
rect 19156 20748 19208 20800
rect 19616 20748 19668 20800
rect 20536 20748 20588 20800
rect 21548 20791 21600 20800
rect 21548 20757 21557 20791
rect 21557 20757 21591 20791
rect 21591 20757 21600 20791
rect 21548 20748 21600 20757
rect 21640 20748 21692 20800
rect 25504 20748 25556 20800
rect 25688 20748 25740 20800
rect 26332 20748 26384 20800
rect 28080 20859 28132 20868
rect 28080 20825 28089 20859
rect 28089 20825 28123 20859
rect 28123 20825 28132 20859
rect 28080 20816 28132 20825
rect 28632 20816 28684 20868
rect 30012 20816 30064 20868
rect 30840 21020 30892 21072
rect 31116 21020 31168 21072
rect 31944 21020 31996 21072
rect 35440 21020 35492 21072
rect 30932 20952 30984 21004
rect 34336 20952 34388 21004
rect 32772 20884 32824 20936
rect 33232 20884 33284 20936
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 31944 20859 31996 20868
rect 31944 20825 31953 20859
rect 31953 20825 31987 20859
rect 31987 20825 31996 20859
rect 31944 20816 31996 20825
rect 32220 20816 32272 20868
rect 32496 20859 32548 20868
rect 32496 20825 32505 20859
rect 32505 20825 32539 20859
rect 32539 20825 32548 20859
rect 32496 20816 32548 20825
rect 33876 20816 33928 20868
rect 35900 20816 35952 20868
rect 33048 20791 33100 20800
rect 33048 20757 33057 20791
rect 33057 20757 33091 20791
rect 33091 20757 33100 20791
rect 33048 20748 33100 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6828 20587 6880 20596
rect 6828 20553 6837 20587
rect 6837 20553 6871 20587
rect 6871 20553 6880 20587
rect 6828 20544 6880 20553
rect 12808 20544 12860 20596
rect 1860 20408 1912 20460
rect 7564 20408 7616 20460
rect 13084 20476 13136 20528
rect 13268 20476 13320 20528
rect 15292 20476 15344 20528
rect 17224 20544 17276 20596
rect 19984 20544 20036 20596
rect 21548 20544 21600 20596
rect 16764 20476 16816 20528
rect 17040 20519 17092 20528
rect 17040 20485 17049 20519
rect 17049 20485 17083 20519
rect 17083 20485 17092 20519
rect 17040 20476 17092 20485
rect 18880 20519 18932 20528
rect 18880 20485 18889 20519
rect 18889 20485 18923 20519
rect 18923 20485 18932 20519
rect 18880 20476 18932 20485
rect 22192 20519 22244 20528
rect 22192 20485 22201 20519
rect 22201 20485 22235 20519
rect 22235 20485 22244 20519
rect 22192 20476 22244 20485
rect 22284 20476 22336 20528
rect 22560 20476 22612 20528
rect 23756 20476 23808 20528
rect 24216 20544 24268 20596
rect 25412 20544 25464 20596
rect 25504 20544 25556 20596
rect 29460 20544 29512 20596
rect 29736 20544 29788 20596
rect 30012 20544 30064 20596
rect 30932 20544 30984 20596
rect 31300 20544 31352 20596
rect 31576 20544 31628 20596
rect 24400 20476 24452 20528
rect 25228 20476 25280 20528
rect 27344 20519 27396 20528
rect 27344 20485 27353 20519
rect 27353 20485 27387 20519
rect 27387 20485 27396 20519
rect 27344 20476 27396 20485
rect 30380 20476 30432 20528
rect 32404 20519 32456 20528
rect 12900 20408 12952 20460
rect 13360 20408 13412 20460
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 14556 20340 14608 20392
rect 14832 20340 14884 20392
rect 15200 20383 15252 20392
rect 15200 20349 15209 20383
rect 15209 20349 15243 20383
rect 15243 20349 15252 20383
rect 15200 20340 15252 20349
rect 17868 20383 17920 20392
rect 6644 20272 6696 20324
rect 17868 20349 17877 20383
rect 17877 20349 17911 20383
rect 17911 20349 17920 20383
rect 17868 20340 17920 20349
rect 18236 20340 18288 20392
rect 1768 20247 1820 20256
rect 1768 20213 1777 20247
rect 1777 20213 1811 20247
rect 1811 20213 1820 20247
rect 1768 20204 1820 20213
rect 11704 20204 11756 20256
rect 12348 20204 12400 20256
rect 14464 20204 14516 20256
rect 16396 20204 16448 20256
rect 16764 20204 16816 20256
rect 17776 20204 17828 20256
rect 18236 20204 18288 20256
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 20076 20340 20128 20392
rect 22376 20340 22428 20392
rect 22560 20340 22612 20392
rect 24216 20340 24268 20392
rect 24308 20383 24360 20392
rect 24308 20349 24317 20383
rect 24317 20349 24351 20383
rect 24351 20349 24360 20383
rect 24308 20340 24360 20349
rect 22284 20272 22336 20324
rect 22836 20272 22888 20324
rect 25780 20408 25832 20460
rect 26884 20408 26936 20460
rect 27068 20408 27120 20460
rect 27620 20383 27672 20392
rect 21456 20204 21508 20256
rect 23020 20204 23072 20256
rect 26240 20247 26292 20256
rect 26240 20213 26249 20247
rect 26249 20213 26283 20247
rect 26283 20213 26292 20247
rect 26240 20204 26292 20213
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 27896 20340 27948 20392
rect 28816 20383 28868 20392
rect 28816 20349 28825 20383
rect 28825 20349 28859 20383
rect 28859 20349 28868 20383
rect 28816 20340 28868 20349
rect 29000 20340 29052 20392
rect 29460 20340 29512 20392
rect 30380 20340 30432 20392
rect 32404 20485 32413 20519
rect 32413 20485 32447 20519
rect 32447 20485 32456 20519
rect 32404 20476 32456 20485
rect 33416 20476 33468 20528
rect 34060 20476 34112 20528
rect 33692 20408 33744 20460
rect 34152 20451 34204 20460
rect 34152 20417 34161 20451
rect 34161 20417 34195 20451
rect 34195 20417 34204 20451
rect 34152 20408 34204 20417
rect 27436 20272 27488 20324
rect 30564 20272 30616 20324
rect 31024 20272 31076 20324
rect 29920 20204 29972 20256
rect 30196 20204 30248 20256
rect 32956 20315 33008 20324
rect 32956 20281 32965 20315
rect 32965 20281 32999 20315
rect 32999 20281 33008 20315
rect 32956 20272 33008 20281
rect 32128 20204 32180 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7932 20000 7984 20052
rect 15568 20000 15620 20052
rect 15936 20000 15988 20052
rect 17500 20000 17552 20052
rect 17776 20000 17828 20052
rect 23664 20000 23716 20052
rect 6184 19932 6236 19984
rect 13176 19932 13228 19984
rect 15844 19932 15896 19984
rect 20168 19932 20220 19984
rect 20628 19932 20680 19984
rect 22100 19932 22152 19984
rect 11612 19864 11664 19916
rect 12348 19864 12400 19916
rect 21916 19864 21968 19916
rect 24032 19932 24084 19984
rect 23756 19864 23808 19916
rect 25136 20000 25188 20052
rect 25872 20000 25924 20052
rect 26148 20000 26200 20052
rect 28356 20000 28408 20052
rect 25320 19932 25372 19984
rect 28264 19932 28316 19984
rect 25044 19864 25096 19916
rect 27436 19907 27488 19916
rect 27436 19873 27445 19907
rect 27445 19873 27479 19907
rect 27479 19873 27488 19907
rect 27436 19864 27488 19873
rect 28724 19907 28776 19916
rect 28724 19873 28733 19907
rect 28733 19873 28767 19907
rect 28767 19873 28776 19907
rect 28724 19864 28776 19873
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 13636 19796 13688 19848
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 15568 19796 15620 19848
rect 16672 19839 16724 19848
rect 16672 19805 16681 19839
rect 16681 19805 16715 19839
rect 16715 19805 16724 19839
rect 16672 19796 16724 19805
rect 17500 19796 17552 19848
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 26148 19839 26200 19848
rect 26148 19805 26157 19839
rect 26157 19805 26191 19839
rect 26191 19805 26200 19839
rect 26148 19796 26200 19805
rect 27988 19796 28040 19848
rect 29552 19932 29604 19984
rect 10968 19728 11020 19780
rect 11704 19771 11756 19780
rect 11704 19737 11713 19771
rect 11713 19737 11747 19771
rect 11747 19737 11756 19771
rect 11704 19728 11756 19737
rect 8576 19660 8628 19712
rect 15108 19728 15160 19780
rect 15476 19771 15528 19780
rect 15476 19737 15485 19771
rect 15485 19737 15519 19771
rect 15519 19737 15528 19771
rect 15476 19728 15528 19737
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 14004 19660 14056 19712
rect 14740 19660 14792 19712
rect 15016 19660 15068 19712
rect 18144 19771 18196 19780
rect 18144 19737 18153 19771
rect 18153 19737 18187 19771
rect 18187 19737 18196 19771
rect 18144 19728 18196 19737
rect 18880 19728 18932 19780
rect 21456 19771 21508 19780
rect 19340 19660 19392 19712
rect 21456 19737 21465 19771
rect 21465 19737 21499 19771
rect 21499 19737 21508 19771
rect 21456 19728 21508 19737
rect 22376 19771 22428 19780
rect 22376 19737 22385 19771
rect 22385 19737 22419 19771
rect 22419 19737 22428 19771
rect 22376 19728 22428 19737
rect 23020 19771 23072 19780
rect 23020 19737 23029 19771
rect 23029 19737 23063 19771
rect 23063 19737 23072 19771
rect 23020 19728 23072 19737
rect 24216 19728 24268 19780
rect 20904 19660 20956 19712
rect 22560 19660 22612 19712
rect 23664 19660 23716 19712
rect 27896 19728 27948 19780
rect 29368 19728 29420 19780
rect 30196 20000 30248 20052
rect 30380 20000 30432 20052
rect 31024 19932 31076 19984
rect 31944 20000 31996 20052
rect 33416 20000 33468 20052
rect 29920 19864 29972 19916
rect 34612 19864 34664 19916
rect 38752 19864 38804 19916
rect 30564 19796 30616 19848
rect 31944 19796 31996 19848
rect 32220 19796 32272 19848
rect 32312 19839 32364 19848
rect 32312 19805 32321 19839
rect 32321 19805 32355 19839
rect 32355 19805 32364 19839
rect 32956 19839 33008 19848
rect 32312 19796 32364 19805
rect 32956 19805 32965 19839
rect 32965 19805 32999 19839
rect 32999 19805 33008 19839
rect 32956 19796 33008 19805
rect 34152 19796 34204 19848
rect 34796 19796 34848 19848
rect 31208 19771 31260 19780
rect 28816 19660 28868 19712
rect 29736 19660 29788 19712
rect 31208 19737 31217 19771
rect 31217 19737 31251 19771
rect 31251 19737 31260 19771
rect 31208 19728 31260 19737
rect 31300 19771 31352 19780
rect 31300 19737 31309 19771
rect 31309 19737 31343 19771
rect 31343 19737 31352 19771
rect 31300 19728 31352 19737
rect 30196 19660 30248 19712
rect 31392 19660 31444 19712
rect 34428 19728 34480 19780
rect 38108 19771 38160 19780
rect 38108 19737 38117 19771
rect 38117 19737 38151 19771
rect 38151 19737 38160 19771
rect 38108 19728 38160 19737
rect 32404 19703 32456 19712
rect 32404 19669 32413 19703
rect 32413 19669 32447 19703
rect 32447 19669 32456 19703
rect 32404 19660 32456 19669
rect 33324 19660 33376 19712
rect 34704 19660 34756 19712
rect 35348 19660 35400 19712
rect 37648 19660 37700 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 7564 19499 7616 19508
rect 7564 19465 7573 19499
rect 7573 19465 7607 19499
rect 7607 19465 7616 19499
rect 7564 19456 7616 19465
rect 8484 19456 8536 19508
rect 10968 19456 11020 19508
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 13268 19456 13320 19508
rect 14280 19456 14332 19508
rect 1768 19320 1820 19372
rect 5448 19320 5500 19372
rect 9772 19388 9824 19440
rect 10140 19431 10192 19440
rect 10140 19397 10149 19431
rect 10149 19397 10183 19431
rect 10183 19397 10192 19431
rect 10140 19388 10192 19397
rect 11796 19388 11848 19440
rect 11980 19388 12032 19440
rect 15016 19388 15068 19440
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 12900 19320 12952 19372
rect 12532 19252 12584 19304
rect 14740 19320 14792 19372
rect 17408 19431 17460 19440
rect 17408 19397 17417 19431
rect 17417 19397 17451 19431
rect 17451 19397 17460 19431
rect 17408 19388 17460 19397
rect 18604 19431 18656 19440
rect 18604 19397 18613 19431
rect 18613 19397 18647 19431
rect 18647 19397 18656 19431
rect 18604 19388 18656 19397
rect 19340 19388 19392 19440
rect 20352 19388 20404 19440
rect 20904 19388 20956 19440
rect 21088 19431 21140 19440
rect 21088 19397 21097 19431
rect 21097 19397 21131 19431
rect 21131 19397 21140 19431
rect 21088 19388 21140 19397
rect 22100 19431 22152 19440
rect 22100 19397 22109 19431
rect 22109 19397 22143 19431
rect 22143 19397 22152 19431
rect 22100 19388 22152 19397
rect 23020 19388 23072 19440
rect 23664 19431 23716 19440
rect 23664 19397 23666 19431
rect 23666 19397 23700 19431
rect 23700 19397 23716 19431
rect 23664 19388 23716 19397
rect 23940 19388 23992 19440
rect 26240 19388 26292 19440
rect 27344 19431 27396 19440
rect 27344 19397 27353 19431
rect 27353 19397 27387 19431
rect 27387 19397 27396 19431
rect 27344 19388 27396 19397
rect 28080 19456 28132 19508
rect 31576 19456 31628 19508
rect 29736 19431 29788 19440
rect 29736 19397 29745 19431
rect 29745 19397 29779 19431
rect 29779 19397 29788 19431
rect 29736 19388 29788 19397
rect 30012 19388 30064 19440
rect 15200 19363 15252 19372
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 15384 19320 15436 19372
rect 16304 19320 16356 19372
rect 16396 19320 16448 19372
rect 21824 19320 21876 19372
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 22836 19363 22888 19372
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 20076 19295 20128 19304
rect 6552 19184 6604 19236
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 18880 19184 18932 19236
rect 20076 19261 20085 19295
rect 20085 19261 20119 19295
rect 20119 19261 20128 19295
rect 20076 19252 20128 19261
rect 22836 19329 22845 19363
rect 22845 19329 22879 19363
rect 22879 19329 22888 19363
rect 22836 19320 22888 19329
rect 23388 19320 23440 19372
rect 24124 19295 24176 19304
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 27068 19320 27120 19372
rect 27252 19295 27304 19304
rect 27252 19261 27261 19295
rect 27261 19261 27295 19295
rect 27295 19261 27304 19295
rect 27252 19252 27304 19261
rect 27344 19252 27396 19304
rect 28448 19320 28500 19372
rect 28540 19320 28592 19372
rect 28908 19320 28960 19372
rect 29460 19320 29512 19372
rect 33324 19456 33376 19508
rect 32404 19388 32456 19440
rect 36268 19499 36320 19508
rect 36268 19465 36277 19499
rect 36277 19465 36311 19499
rect 36311 19465 36320 19499
rect 36268 19456 36320 19465
rect 38016 19456 38068 19508
rect 33508 19431 33560 19440
rect 33508 19397 33517 19431
rect 33517 19397 33551 19431
rect 33551 19397 33560 19431
rect 33508 19388 33560 19397
rect 34060 19388 34112 19440
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 34520 19363 34572 19372
rect 34520 19329 34529 19363
rect 34529 19329 34563 19363
rect 34563 19329 34572 19363
rect 34520 19320 34572 19329
rect 38292 19363 38344 19372
rect 28356 19252 28408 19304
rect 29644 19295 29696 19304
rect 20720 19184 20772 19236
rect 29644 19261 29653 19295
rect 29653 19261 29687 19295
rect 29687 19261 29696 19295
rect 29644 19252 29696 19261
rect 30012 19295 30064 19304
rect 30012 19261 30021 19295
rect 30021 19261 30055 19295
rect 30055 19261 30064 19295
rect 30012 19252 30064 19261
rect 30932 19252 30984 19304
rect 24492 19116 24544 19168
rect 26976 19116 27028 19168
rect 27068 19116 27120 19168
rect 28540 19116 28592 19168
rect 28724 19116 28776 19168
rect 30012 19116 30064 19168
rect 30656 19116 30708 19168
rect 33140 19252 33192 19304
rect 33232 19252 33284 19304
rect 38292 19329 38301 19363
rect 38301 19329 38335 19363
rect 38335 19329 38344 19363
rect 38292 19320 38344 19329
rect 37464 19252 37516 19304
rect 31576 19184 31628 19236
rect 33508 19184 33560 19236
rect 32404 19159 32456 19168
rect 32404 19125 32413 19159
rect 32413 19125 32447 19159
rect 32447 19125 32456 19159
rect 32404 19116 32456 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 10140 18912 10192 18964
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 17408 18912 17460 18964
rect 18604 18955 18656 18964
rect 18604 18921 18613 18955
rect 18613 18921 18647 18955
rect 18647 18921 18656 18955
rect 18604 18912 18656 18921
rect 14648 18844 14700 18896
rect 19524 18912 19576 18964
rect 19892 18912 19944 18964
rect 24216 18912 24268 18964
rect 25964 18912 26016 18964
rect 18880 18844 18932 18896
rect 27252 18844 27304 18896
rect 28080 18912 28132 18964
rect 29828 18912 29880 18964
rect 31024 18912 31076 18964
rect 27436 18844 27488 18896
rect 27528 18844 27580 18896
rect 29000 18844 29052 18896
rect 34428 18912 34480 18964
rect 16580 18776 16632 18828
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 11152 18683 11204 18692
rect 11152 18649 11161 18683
rect 11161 18649 11195 18683
rect 11195 18649 11204 18683
rect 11152 18640 11204 18649
rect 11244 18640 11296 18692
rect 15568 18708 15620 18760
rect 16120 18708 16172 18760
rect 18604 18776 18656 18828
rect 19340 18776 19392 18828
rect 23204 18776 23256 18828
rect 31116 18776 31168 18828
rect 34888 18844 34940 18896
rect 31668 18776 31720 18828
rect 33140 18819 33192 18828
rect 33140 18785 33149 18819
rect 33149 18785 33183 18819
rect 33183 18785 33192 18819
rect 33140 18776 33192 18785
rect 35900 18776 35952 18828
rect 38568 18776 38620 18828
rect 18052 18708 18104 18760
rect 19064 18708 19116 18760
rect 19892 18640 19944 18692
rect 21640 18708 21692 18760
rect 22284 18708 22336 18760
rect 24492 18708 24544 18760
rect 28264 18708 28316 18760
rect 34704 18708 34756 18760
rect 38844 18708 38896 18760
rect 8576 18572 8628 18624
rect 9680 18572 9732 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 16120 18572 16172 18624
rect 23020 18683 23072 18692
rect 23020 18649 23029 18683
rect 23029 18649 23063 18683
rect 23063 18649 23072 18683
rect 25780 18683 25832 18692
rect 23020 18640 23072 18649
rect 25780 18649 25789 18683
rect 25789 18649 25823 18683
rect 25823 18649 25832 18683
rect 25780 18640 25832 18649
rect 20720 18615 20772 18624
rect 20720 18581 20729 18615
rect 20729 18581 20763 18615
rect 20763 18581 20772 18615
rect 20720 18572 20772 18581
rect 21916 18572 21968 18624
rect 22836 18572 22888 18624
rect 23664 18572 23716 18624
rect 25688 18572 25740 18624
rect 26700 18640 26752 18692
rect 27344 18683 27396 18692
rect 27344 18649 27353 18683
rect 27353 18649 27387 18683
rect 27387 18649 27396 18683
rect 27344 18640 27396 18649
rect 27436 18683 27488 18692
rect 27436 18649 27445 18683
rect 27445 18649 27479 18683
rect 27479 18649 27488 18683
rect 27436 18640 27488 18649
rect 27620 18640 27672 18692
rect 27988 18640 28040 18692
rect 28540 18640 28592 18692
rect 27896 18572 27948 18624
rect 28724 18572 28776 18624
rect 29920 18683 29972 18692
rect 29920 18649 29929 18683
rect 29929 18649 29963 18683
rect 29963 18649 29972 18683
rect 29920 18640 29972 18649
rect 30656 18640 30708 18692
rect 31024 18683 31076 18692
rect 31024 18649 31033 18683
rect 31033 18649 31067 18683
rect 31067 18649 31076 18683
rect 31024 18640 31076 18649
rect 30932 18572 30984 18624
rect 32036 18640 32088 18692
rect 34060 18640 34112 18692
rect 32312 18572 32364 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 8300 18368 8352 18420
rect 11520 18368 11572 18420
rect 15660 18411 15712 18420
rect 15660 18377 15669 18411
rect 15669 18377 15703 18411
rect 15703 18377 15712 18411
rect 15660 18368 15712 18377
rect 6736 18343 6788 18352
rect 6736 18309 6745 18343
rect 6745 18309 6779 18343
rect 6779 18309 6788 18343
rect 6736 18300 6788 18309
rect 12164 18343 12216 18352
rect 12164 18309 12173 18343
rect 12173 18309 12207 18343
rect 12207 18309 12216 18343
rect 12164 18300 12216 18309
rect 12716 18343 12768 18352
rect 12716 18309 12725 18343
rect 12725 18309 12759 18343
rect 12759 18309 12768 18343
rect 12716 18300 12768 18309
rect 12900 18300 12952 18352
rect 13912 18300 13964 18352
rect 15108 18300 15160 18352
rect 23664 18368 23716 18420
rect 18052 18343 18104 18352
rect 18052 18309 18061 18343
rect 18061 18309 18095 18343
rect 18095 18309 18104 18343
rect 18052 18300 18104 18309
rect 18144 18300 18196 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 8024 18232 8076 18284
rect 6092 18164 6144 18216
rect 7656 18207 7708 18216
rect 7656 18173 7665 18207
rect 7665 18173 7699 18207
rect 7699 18173 7708 18207
rect 7656 18164 7708 18173
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 8944 18164 8996 18216
rect 11152 18096 11204 18148
rect 17592 18232 17644 18284
rect 18328 18207 18380 18216
rect 18328 18173 18337 18207
rect 18337 18173 18371 18207
rect 18371 18173 18380 18207
rect 18328 18164 18380 18173
rect 19892 18300 19944 18352
rect 21088 18300 21140 18352
rect 25964 18368 26016 18420
rect 28632 18368 28684 18420
rect 25320 18300 25372 18352
rect 26332 18300 26384 18352
rect 27252 18300 27304 18352
rect 28908 18368 28960 18420
rect 30288 18368 30340 18420
rect 30932 18368 30984 18420
rect 28816 18300 28868 18352
rect 29644 18300 29696 18352
rect 33968 18368 34020 18420
rect 34888 18411 34940 18420
rect 34888 18377 34897 18411
rect 34897 18377 34931 18411
rect 34931 18377 34940 18411
rect 34888 18368 34940 18377
rect 20076 18232 20128 18284
rect 23664 18232 23716 18284
rect 28540 18275 28592 18284
rect 9312 18028 9364 18080
rect 9404 18028 9456 18080
rect 10140 18028 10192 18080
rect 10600 18028 10652 18080
rect 20352 18096 20404 18148
rect 23204 18164 23256 18216
rect 24768 18207 24820 18216
rect 24768 18173 24777 18207
rect 24777 18173 24811 18207
rect 24811 18173 24820 18207
rect 24768 18164 24820 18173
rect 28080 18164 28132 18216
rect 28540 18241 28549 18275
rect 28549 18241 28583 18275
rect 28583 18241 28592 18275
rect 28540 18232 28592 18241
rect 18328 18028 18380 18080
rect 18604 18028 18656 18080
rect 19432 18028 19484 18080
rect 20076 18028 20128 18080
rect 20720 18028 20772 18080
rect 22192 18028 22244 18080
rect 23020 18071 23072 18080
rect 23020 18037 23029 18071
rect 23029 18037 23063 18071
rect 23063 18037 23072 18071
rect 23020 18028 23072 18037
rect 28908 18164 28960 18216
rect 33048 18232 33100 18284
rect 33508 18275 33560 18284
rect 30196 18207 30248 18216
rect 30196 18173 30205 18207
rect 30205 18173 30239 18207
rect 30239 18173 30248 18207
rect 30196 18164 30248 18173
rect 31116 18164 31168 18216
rect 31576 18164 31628 18216
rect 32036 18164 32088 18216
rect 33508 18241 33517 18275
rect 33517 18241 33551 18275
rect 33551 18241 33560 18275
rect 33508 18232 33560 18241
rect 37464 18300 37516 18352
rect 35624 18275 35676 18284
rect 35624 18241 35633 18275
rect 35633 18241 35667 18275
rect 35667 18241 35676 18275
rect 35624 18232 35676 18241
rect 38108 18275 38160 18284
rect 38108 18241 38117 18275
rect 38117 18241 38151 18275
rect 38151 18241 38160 18275
rect 38108 18232 38160 18241
rect 33232 18096 33284 18148
rect 37280 18096 37332 18148
rect 27528 18028 27580 18080
rect 27896 18028 27948 18080
rect 28264 18028 28316 18080
rect 28632 18028 28684 18080
rect 32772 18028 32824 18080
rect 37924 18028 37976 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 6736 17824 6788 17876
rect 15016 17824 15068 17876
rect 16488 17824 16540 17876
rect 16580 17824 16632 17876
rect 20812 17824 20864 17876
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 21456 17824 21508 17876
rect 9404 17756 9456 17808
rect 11704 17756 11756 17808
rect 8576 17688 8628 17740
rect 15108 17756 15160 17808
rect 15384 17756 15436 17808
rect 25688 17756 25740 17808
rect 25780 17756 25832 17808
rect 26608 17756 26660 17808
rect 27344 17799 27396 17808
rect 14924 17688 14976 17740
rect 16580 17688 16632 17740
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 8760 17620 8812 17672
rect 10600 17620 10652 17672
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 9036 17552 9088 17604
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 9680 17552 9732 17604
rect 7012 17484 7064 17536
rect 8208 17484 8260 17536
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 11796 17552 11848 17604
rect 12992 17552 13044 17604
rect 15476 17620 15528 17672
rect 16120 17620 16172 17672
rect 24492 17688 24544 17740
rect 26056 17688 26108 17740
rect 27344 17765 27353 17799
rect 27353 17765 27387 17799
rect 27387 17765 27396 17799
rect 27344 17756 27396 17765
rect 27160 17688 27212 17740
rect 27712 17688 27764 17740
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 16488 17552 16540 17604
rect 13728 17484 13780 17536
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 15292 17484 15344 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 16028 17484 16080 17536
rect 16856 17552 16908 17604
rect 19524 17620 19576 17672
rect 21548 17620 21600 17672
rect 23572 17620 23624 17672
rect 19340 17552 19392 17604
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 18144 17484 18196 17493
rect 20720 17552 20772 17604
rect 20812 17552 20864 17604
rect 21916 17595 21968 17604
rect 21916 17561 21925 17595
rect 21925 17561 21959 17595
rect 21959 17561 21968 17595
rect 21916 17552 21968 17561
rect 24676 17552 24728 17604
rect 25596 17552 25648 17604
rect 25688 17595 25740 17604
rect 25688 17561 25697 17595
rect 25697 17561 25731 17595
rect 25731 17561 25740 17595
rect 25688 17552 25740 17561
rect 32404 17756 32456 17808
rect 28264 17688 28316 17740
rect 29736 17688 29788 17740
rect 28448 17620 28500 17672
rect 19892 17484 19944 17536
rect 21456 17484 21508 17536
rect 21732 17484 21784 17536
rect 22560 17484 22612 17536
rect 23940 17484 23992 17536
rect 30932 17620 30984 17672
rect 30012 17595 30064 17604
rect 30012 17561 30021 17595
rect 30021 17561 30055 17595
rect 30055 17561 30064 17595
rect 30012 17552 30064 17561
rect 30104 17595 30156 17604
rect 30104 17561 30113 17595
rect 30113 17561 30147 17595
rect 30147 17561 30156 17595
rect 30104 17552 30156 17561
rect 30472 17552 30524 17604
rect 31300 17552 31352 17604
rect 31576 17595 31628 17604
rect 31576 17561 31585 17595
rect 31585 17561 31619 17595
rect 31619 17561 31628 17595
rect 31576 17552 31628 17561
rect 31116 17484 31168 17536
rect 31852 17552 31904 17604
rect 32220 17595 32272 17604
rect 32220 17561 32229 17595
rect 32229 17561 32263 17595
rect 32263 17561 32272 17595
rect 32220 17552 32272 17561
rect 32772 17867 32824 17876
rect 32772 17833 32781 17867
rect 32781 17833 32815 17867
rect 32815 17833 32824 17867
rect 32772 17824 32824 17833
rect 32864 17756 32916 17808
rect 34520 17756 34572 17808
rect 33232 17688 33284 17740
rect 33324 17663 33376 17672
rect 33324 17629 33333 17663
rect 33333 17629 33367 17663
rect 33367 17629 33376 17663
rect 33324 17620 33376 17629
rect 33968 17663 34020 17672
rect 33968 17629 33977 17663
rect 33977 17629 34011 17663
rect 34011 17629 34020 17663
rect 33968 17620 34020 17629
rect 33048 17484 33100 17536
rect 33140 17484 33192 17536
rect 37188 17484 37240 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7012 17255 7064 17264
rect 7012 17221 7021 17255
rect 7021 17221 7055 17255
rect 7055 17221 7064 17255
rect 7012 17212 7064 17221
rect 9680 17280 9732 17332
rect 11704 17280 11756 17332
rect 8116 17255 8168 17264
rect 8116 17221 8125 17255
rect 8125 17221 8159 17255
rect 8159 17221 8168 17255
rect 8116 17212 8168 17221
rect 8208 17255 8260 17264
rect 8208 17221 8217 17255
rect 8217 17221 8251 17255
rect 8251 17221 8260 17255
rect 8208 17212 8260 17221
rect 9772 17212 9824 17264
rect 10508 17212 10560 17264
rect 10876 17212 10928 17264
rect 5080 17144 5132 17196
rect 5448 17144 5500 17196
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 10968 17187 11020 17196
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 6736 17076 6788 17128
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 14464 17187 14516 17196
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 11428 17076 11480 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 12716 17076 12768 17128
rect 16856 17280 16908 17332
rect 18052 17280 18104 17332
rect 15200 17212 15252 17264
rect 18328 17255 18380 17264
rect 14832 17076 14884 17128
rect 15660 17119 15712 17128
rect 15660 17085 15669 17119
rect 15669 17085 15703 17119
rect 15703 17085 15712 17119
rect 18328 17221 18337 17255
rect 18337 17221 18371 17255
rect 18371 17221 18380 17255
rect 18328 17212 18380 17221
rect 20076 17212 20128 17264
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 17040 17144 17092 17196
rect 20812 17212 20864 17264
rect 21732 17212 21784 17264
rect 23296 17212 23348 17264
rect 15660 17076 15712 17085
rect 18420 17076 18472 17128
rect 8208 17008 8260 17060
rect 12256 17008 12308 17060
rect 17960 17008 18012 17060
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 13544 16983 13596 16992
rect 13544 16949 13553 16983
rect 13553 16949 13587 16983
rect 13587 16949 13596 16983
rect 13544 16940 13596 16949
rect 15108 16940 15160 16992
rect 17868 16940 17920 16992
rect 20444 17144 20496 17196
rect 20076 17076 20128 17128
rect 21272 17076 21324 17128
rect 23296 17119 23348 17128
rect 23296 17085 23305 17119
rect 23305 17085 23339 17119
rect 23339 17085 23348 17119
rect 23296 17076 23348 17085
rect 23940 17255 23992 17264
rect 23940 17221 23949 17255
rect 23949 17221 23983 17255
rect 23983 17221 23992 17255
rect 23940 17212 23992 17221
rect 27620 17280 27672 17332
rect 30288 17280 30340 17332
rect 32312 17280 32364 17332
rect 33048 17323 33100 17332
rect 33048 17289 33057 17323
rect 33057 17289 33091 17323
rect 33091 17289 33100 17323
rect 33048 17280 33100 17289
rect 35624 17280 35676 17332
rect 25504 17255 25556 17264
rect 25504 17221 25513 17255
rect 25513 17221 25547 17255
rect 25547 17221 25556 17255
rect 25504 17212 25556 17221
rect 24032 17076 24084 17128
rect 25504 17076 25556 17128
rect 28264 17212 28316 17264
rect 30104 17212 30156 17264
rect 31300 17212 31352 17264
rect 34796 17212 34848 17264
rect 27804 17144 27856 17196
rect 26424 17119 26476 17128
rect 26424 17085 26433 17119
rect 26433 17085 26467 17119
rect 26467 17085 26476 17119
rect 26424 17076 26476 17085
rect 27344 17119 27396 17128
rect 27344 17085 27353 17119
rect 27353 17085 27387 17119
rect 27387 17085 27396 17119
rect 27344 17076 27396 17085
rect 27988 17076 28040 17128
rect 29368 17119 29420 17128
rect 29368 17085 29377 17119
rect 29377 17085 29411 17119
rect 29411 17085 29420 17119
rect 29368 17076 29420 17085
rect 30656 17076 30708 17128
rect 30748 17076 30800 17128
rect 32312 17187 32364 17196
rect 32312 17153 32321 17187
rect 32321 17153 32355 17187
rect 32355 17153 32364 17187
rect 32312 17144 32364 17153
rect 32956 17187 33008 17196
rect 32956 17153 32965 17187
rect 32965 17153 32999 17187
rect 32999 17153 33008 17187
rect 32956 17144 33008 17153
rect 38292 17187 38344 17196
rect 31024 17119 31076 17128
rect 31024 17085 31033 17119
rect 31033 17085 31067 17119
rect 31067 17085 31076 17119
rect 31024 17076 31076 17085
rect 20720 17008 20772 17060
rect 38292 17153 38301 17187
rect 38301 17153 38335 17187
rect 38335 17153 38344 17187
rect 38292 17144 38344 17153
rect 20812 16940 20864 16992
rect 24768 16940 24820 16992
rect 26424 16940 26476 16992
rect 29368 16940 29420 16992
rect 30656 16940 30708 16992
rect 38108 16983 38160 16992
rect 38108 16949 38117 16983
rect 38117 16949 38151 16983
rect 38151 16949 38160 16983
rect 38108 16940 38160 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 12256 16736 12308 16788
rect 12716 16736 12768 16788
rect 9404 16668 9456 16720
rect 10968 16668 11020 16720
rect 16212 16736 16264 16788
rect 16948 16736 17000 16788
rect 5264 16600 5316 16652
rect 7380 16643 7432 16652
rect 7380 16609 7389 16643
rect 7389 16609 7423 16643
rect 7423 16609 7432 16643
rect 7380 16600 7432 16609
rect 8300 16600 8352 16652
rect 11428 16532 11480 16584
rect 12164 16532 12216 16584
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 13452 16668 13504 16720
rect 13820 16668 13872 16720
rect 16396 16668 16448 16720
rect 19892 16736 19944 16788
rect 20536 16736 20588 16788
rect 20812 16736 20864 16788
rect 13728 16600 13780 16652
rect 16120 16600 16172 16652
rect 13452 16532 13504 16584
rect 15200 16532 15252 16584
rect 18604 16600 18656 16652
rect 21732 16668 21784 16720
rect 25504 16736 25556 16788
rect 25596 16736 25648 16788
rect 26424 16736 26476 16788
rect 30196 16736 30248 16788
rect 24492 16668 24544 16720
rect 24860 16600 24912 16652
rect 29460 16668 29512 16720
rect 18512 16532 18564 16584
rect 19340 16532 19392 16584
rect 24584 16575 24636 16584
rect 2228 16464 2280 16516
rect 5816 16464 5868 16516
rect 9220 16507 9272 16516
rect 9220 16473 9229 16507
rect 9229 16473 9263 16507
rect 9263 16473 9272 16507
rect 9220 16464 9272 16473
rect 10232 16507 10284 16516
rect 1492 16396 1544 16448
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 6920 16396 6972 16448
rect 9036 16396 9088 16448
rect 10232 16473 10241 16507
rect 10241 16473 10275 16507
rect 10275 16473 10284 16507
rect 10232 16464 10284 16473
rect 10600 16464 10652 16516
rect 15660 16507 15712 16516
rect 15660 16473 15669 16507
rect 15669 16473 15703 16507
rect 15703 16473 15712 16507
rect 15660 16464 15712 16473
rect 10968 16396 11020 16448
rect 11796 16396 11848 16448
rect 12624 16396 12676 16448
rect 12716 16396 12768 16448
rect 13084 16396 13136 16448
rect 13360 16396 13412 16448
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 14924 16396 14976 16448
rect 15108 16396 15160 16448
rect 17960 16464 18012 16516
rect 19892 16464 19944 16516
rect 20536 16464 20588 16516
rect 21456 16464 21508 16516
rect 22192 16464 22244 16516
rect 23020 16464 23072 16516
rect 17316 16396 17368 16448
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 19432 16396 19484 16448
rect 20260 16396 20312 16448
rect 20904 16396 20956 16448
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 27804 16600 27856 16652
rect 28724 16600 28776 16652
rect 31668 16736 31720 16788
rect 34704 16736 34756 16788
rect 31024 16668 31076 16720
rect 32680 16668 32732 16720
rect 25320 16532 25372 16541
rect 28632 16532 28684 16584
rect 31760 16600 31812 16652
rect 37556 16668 37608 16720
rect 38108 16600 38160 16652
rect 25688 16464 25740 16516
rect 23296 16396 23348 16448
rect 23388 16396 23440 16448
rect 25504 16396 25556 16448
rect 27804 16464 27856 16516
rect 28264 16464 28316 16516
rect 28816 16464 28868 16516
rect 29644 16464 29696 16516
rect 30012 16464 30064 16516
rect 30932 16464 30984 16516
rect 31392 16464 31444 16516
rect 31852 16464 31904 16516
rect 32588 16507 32640 16516
rect 32588 16473 32597 16507
rect 32597 16473 32631 16507
rect 32631 16473 32640 16507
rect 33508 16507 33560 16516
rect 32588 16464 32640 16473
rect 33508 16473 33517 16507
rect 33517 16473 33551 16507
rect 33551 16473 33560 16507
rect 33508 16464 33560 16473
rect 27160 16396 27212 16448
rect 27252 16396 27304 16448
rect 34060 16439 34112 16448
rect 34060 16405 34069 16439
rect 34069 16405 34103 16439
rect 34103 16405 34112 16439
rect 34060 16396 34112 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 8484 16192 8536 16244
rect 10324 16192 10376 16244
rect 13636 16192 13688 16244
rect 14280 16192 14332 16244
rect 15660 16192 15712 16244
rect 24124 16235 24176 16244
rect 6828 16167 6880 16176
rect 6828 16133 6837 16167
rect 6837 16133 6871 16167
rect 6871 16133 6880 16167
rect 6828 16124 6880 16133
rect 8392 16167 8444 16176
rect 8392 16133 8401 16167
rect 8401 16133 8435 16167
rect 8435 16133 8444 16167
rect 8392 16124 8444 16133
rect 10232 16167 10284 16176
rect 10232 16133 10241 16167
rect 10241 16133 10275 16167
rect 10275 16133 10284 16167
rect 10232 16124 10284 16133
rect 10784 16124 10836 16176
rect 12072 16124 12124 16176
rect 12808 16167 12860 16176
rect 12808 16133 12817 16167
rect 12817 16133 12851 16167
rect 12851 16133 12860 16167
rect 12808 16124 12860 16133
rect 13544 16124 13596 16176
rect 8576 15988 8628 16040
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 10140 16031 10192 16040
rect 8668 15988 8720 15997
rect 10140 15997 10149 16031
rect 10149 15997 10183 16031
rect 10183 15997 10192 16031
rect 10140 15988 10192 15997
rect 10508 15988 10560 16040
rect 12992 16056 13044 16108
rect 13636 16056 13688 16108
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 16028 15988 16080 16040
rect 16212 15988 16264 16040
rect 16764 16124 16816 16176
rect 17316 16124 17368 16176
rect 18144 16124 18196 16176
rect 19340 16124 19392 16176
rect 20168 16124 20220 16176
rect 22008 16124 22060 16176
rect 22468 16167 22520 16176
rect 20536 16056 20588 16108
rect 22192 16056 22244 16108
rect 17960 16031 18012 16040
rect 17960 15997 17969 16031
rect 17969 15997 18003 16031
rect 18003 15997 18012 16031
rect 17960 15988 18012 15997
rect 18788 16031 18840 16040
rect 18788 15997 18797 16031
rect 18797 15997 18831 16031
rect 18831 15997 18840 16031
rect 18788 15988 18840 15997
rect 22468 16133 22477 16167
rect 22477 16133 22511 16167
rect 22511 16133 22520 16167
rect 22468 16124 22520 16133
rect 22560 16167 22612 16176
rect 22560 16133 22569 16167
rect 22569 16133 22603 16167
rect 22603 16133 22612 16167
rect 22560 16124 22612 16133
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 5172 15852 5224 15904
rect 7012 15852 7064 15904
rect 12808 15852 12860 15904
rect 13636 15852 13688 15904
rect 23112 15920 23164 15972
rect 16764 15852 16816 15904
rect 16856 15852 16908 15904
rect 19616 15852 19668 15904
rect 20260 15852 20312 15904
rect 21824 15852 21876 15904
rect 24124 16201 24133 16235
rect 24133 16201 24167 16235
rect 24167 16201 24176 16235
rect 24124 16192 24176 16201
rect 23480 16124 23532 16176
rect 24032 16099 24084 16108
rect 24032 16065 24041 16099
rect 24041 16065 24075 16099
rect 24075 16065 24084 16099
rect 24032 16056 24084 16065
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 24952 16056 25004 16108
rect 27712 16192 27764 16244
rect 27896 16124 27948 16176
rect 23480 16031 23532 16040
rect 23480 15997 23489 16031
rect 23489 15997 23523 16031
rect 23523 15997 23532 16031
rect 23480 15988 23532 15997
rect 26148 15988 26200 16040
rect 27252 16031 27304 16040
rect 27252 15997 27261 16031
rect 27261 15997 27295 16031
rect 27295 15997 27304 16031
rect 27252 15988 27304 15997
rect 29552 16124 29604 16176
rect 30104 16192 30156 16244
rect 31300 16192 31352 16244
rect 31760 16192 31812 16244
rect 34060 16192 34112 16244
rect 28632 16056 28684 16108
rect 29644 16099 29696 16108
rect 29644 16065 29653 16099
rect 29653 16065 29687 16099
rect 29687 16065 29696 16099
rect 29644 16056 29696 16065
rect 30840 16124 30892 16176
rect 30564 16056 30616 16108
rect 31116 16056 31168 16108
rect 31668 16056 31720 16108
rect 37188 16056 37240 16108
rect 24860 15852 24912 15904
rect 25228 15852 25280 15904
rect 25504 15852 25556 15904
rect 28356 15988 28408 16040
rect 31944 15988 31996 16040
rect 33508 15988 33560 16040
rect 34520 15988 34572 16040
rect 27896 15920 27948 15972
rect 30564 15920 30616 15972
rect 31392 15920 31444 15972
rect 33140 15920 33192 15972
rect 27988 15852 28040 15904
rect 30656 15852 30708 15904
rect 31760 15852 31812 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8300 15648 8352 15700
rect 9036 15648 9088 15700
rect 14556 15648 14608 15700
rect 14924 15648 14976 15700
rect 17684 15648 17736 15700
rect 17776 15648 17828 15700
rect 20076 15648 20128 15700
rect 7012 15580 7064 15632
rect 17960 15580 18012 15632
rect 6736 15512 6788 15564
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 9220 15512 9272 15564
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 12164 15512 12216 15564
rect 4988 15444 5040 15496
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 12440 15444 12492 15496
rect 14280 15512 14332 15564
rect 1676 15419 1728 15428
rect 1676 15385 1685 15419
rect 1685 15385 1719 15419
rect 1719 15385 1728 15419
rect 1676 15376 1728 15385
rect 1860 15419 1912 15428
rect 1860 15385 1869 15419
rect 1869 15385 1903 15419
rect 1903 15385 1912 15419
rect 1860 15376 1912 15385
rect 5908 15419 5960 15428
rect 5908 15385 5917 15419
rect 5917 15385 5951 15419
rect 5951 15385 5960 15419
rect 5908 15376 5960 15385
rect 5448 15308 5500 15360
rect 7012 15376 7064 15428
rect 7380 15419 7432 15428
rect 7380 15385 7389 15419
rect 7389 15385 7423 15419
rect 7423 15385 7432 15419
rect 7380 15376 7432 15385
rect 9772 15419 9824 15428
rect 9772 15385 9781 15419
rect 9781 15385 9815 15419
rect 9815 15385 9824 15419
rect 13452 15444 13504 15496
rect 15200 15512 15252 15564
rect 17776 15512 17828 15564
rect 9772 15376 9824 15385
rect 14372 15376 14424 15428
rect 15844 15444 15896 15496
rect 16396 15444 16448 15496
rect 16856 15444 16908 15496
rect 15384 15376 15436 15428
rect 18420 15444 18472 15496
rect 20720 15580 20772 15632
rect 18972 15512 19024 15564
rect 23112 15648 23164 15700
rect 25136 15648 25188 15700
rect 25320 15648 25372 15700
rect 26332 15648 26384 15700
rect 27436 15648 27488 15700
rect 28080 15648 28132 15700
rect 30472 15691 30524 15700
rect 30472 15657 30481 15691
rect 30481 15657 30515 15691
rect 30515 15657 30524 15691
rect 30472 15648 30524 15657
rect 32588 15648 32640 15700
rect 22560 15580 22612 15632
rect 23020 15580 23072 15632
rect 25412 15580 25464 15632
rect 26148 15580 26200 15632
rect 32772 15580 32824 15632
rect 18880 15444 18932 15496
rect 22284 15512 22336 15564
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 20076 15444 20128 15496
rect 12072 15308 12124 15360
rect 12256 15308 12308 15360
rect 13820 15308 13872 15360
rect 15016 15308 15068 15360
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 16212 15351 16264 15360
rect 16212 15317 16221 15351
rect 16221 15317 16255 15351
rect 16255 15317 16264 15351
rect 16212 15308 16264 15317
rect 17316 15308 17368 15360
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 19340 15376 19392 15428
rect 20168 15376 20220 15428
rect 20076 15308 20128 15360
rect 20352 15351 20404 15360
rect 20352 15317 20361 15351
rect 20361 15317 20395 15351
rect 20395 15317 20404 15351
rect 20352 15308 20404 15317
rect 20812 15444 20864 15496
rect 20720 15376 20772 15428
rect 23296 15512 23348 15564
rect 24860 15555 24912 15564
rect 23664 15487 23716 15496
rect 23664 15453 23673 15487
rect 23673 15453 23707 15487
rect 23707 15453 23716 15487
rect 23664 15444 23716 15453
rect 24400 15444 24452 15496
rect 24860 15521 24869 15555
rect 24869 15521 24903 15555
rect 24903 15521 24912 15555
rect 24860 15512 24912 15521
rect 27620 15512 27672 15564
rect 25136 15444 25188 15496
rect 26516 15444 26568 15496
rect 26608 15444 26660 15496
rect 27436 15444 27488 15496
rect 24492 15376 24544 15428
rect 29000 15444 29052 15496
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 33140 15512 33192 15564
rect 31024 15487 31076 15496
rect 31024 15453 31033 15487
rect 31033 15453 31067 15487
rect 31067 15453 31076 15487
rect 31024 15444 31076 15453
rect 31576 15444 31628 15496
rect 38016 15487 38068 15496
rect 38016 15453 38025 15487
rect 38025 15453 38059 15487
rect 38059 15453 38068 15487
rect 38016 15444 38068 15453
rect 28080 15419 28132 15428
rect 28080 15385 28089 15419
rect 28089 15385 28123 15419
rect 28123 15385 28132 15419
rect 28080 15376 28132 15385
rect 28264 15376 28316 15428
rect 23480 15308 23532 15360
rect 23664 15308 23716 15360
rect 24032 15308 24084 15360
rect 25780 15308 25832 15360
rect 26332 15308 26384 15360
rect 32312 15376 32364 15428
rect 30656 15308 30708 15360
rect 32588 15308 32640 15360
rect 34520 15376 34572 15428
rect 35716 15376 35768 15428
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 8484 15104 8536 15156
rect 6920 15079 6972 15088
rect 6920 15045 6929 15079
rect 6929 15045 6963 15079
rect 6963 15045 6972 15079
rect 6920 15036 6972 15045
rect 8300 15079 8352 15088
rect 8300 15045 8309 15079
rect 8309 15045 8343 15079
rect 8343 15045 8352 15079
rect 8300 15036 8352 15045
rect 10140 15079 10192 15088
rect 10140 15045 10149 15079
rect 10149 15045 10183 15079
rect 10183 15045 10192 15079
rect 10140 15036 10192 15045
rect 15384 15036 15436 15088
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 14464 14968 14516 15020
rect 15476 15011 15528 15020
rect 7012 14900 7064 14952
rect 7840 14900 7892 14952
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 6736 14832 6788 14884
rect 1124 14764 1176 14816
rect 6092 14764 6144 14816
rect 7656 14764 7708 14816
rect 9772 14900 9824 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 13084 14900 13136 14952
rect 14004 14900 14056 14952
rect 15108 14900 15160 14952
rect 12900 14764 12952 14816
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 15844 15104 15896 15156
rect 16488 15104 16540 15156
rect 18328 15036 18380 15088
rect 18696 15079 18748 15088
rect 18696 15045 18705 15079
rect 18705 15045 18739 15079
rect 18739 15045 18748 15079
rect 18696 15036 18748 15045
rect 24400 15104 24452 15156
rect 27344 15104 27396 15156
rect 28172 15104 28224 15156
rect 30104 15104 30156 15156
rect 33416 15104 33468 15156
rect 17776 14968 17828 15020
rect 26148 15036 26200 15088
rect 27252 15036 27304 15088
rect 27896 15036 27948 15088
rect 28080 15036 28132 15088
rect 30656 15079 30708 15088
rect 30656 15045 30665 15079
rect 30665 15045 30699 15079
rect 30699 15045 30708 15079
rect 30656 15036 30708 15045
rect 32220 15036 32272 15088
rect 20812 14968 20864 15020
rect 21732 14968 21784 15020
rect 23756 14968 23808 15020
rect 25136 14968 25188 15020
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 18972 14900 19024 14952
rect 21456 14900 21508 14952
rect 22928 14900 22980 14952
rect 23480 14900 23532 14952
rect 24952 14900 25004 14952
rect 26516 14968 26568 15020
rect 27528 14968 27580 15020
rect 26148 14900 26200 14952
rect 17224 14832 17276 14884
rect 22560 14832 22612 14884
rect 24308 14832 24360 14884
rect 28356 14900 28408 14952
rect 29000 14968 29052 15020
rect 29736 15011 29788 15020
rect 29736 14977 29745 15011
rect 29745 14977 29779 15011
rect 29779 14977 29788 15011
rect 29736 14968 29788 14977
rect 29644 14900 29696 14952
rect 29828 14900 29880 14952
rect 27436 14832 27488 14884
rect 29368 14832 29420 14884
rect 29920 14832 29972 14884
rect 16396 14764 16448 14816
rect 16948 14764 17000 14816
rect 19064 14764 19116 14816
rect 19340 14764 19392 14816
rect 20536 14764 20588 14816
rect 24124 14764 24176 14816
rect 24952 14764 25004 14816
rect 26056 14764 26108 14816
rect 27712 14764 27764 14816
rect 28448 14764 28500 14816
rect 29000 14764 29052 14816
rect 38108 14968 38160 15020
rect 37832 14807 37884 14816
rect 37832 14773 37841 14807
rect 37841 14773 37875 14807
rect 37875 14773 37884 14807
rect 37832 14764 37884 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14560 2372 14612
rect 6552 14560 6604 14612
rect 9036 14560 9088 14612
rect 10048 14560 10100 14612
rect 8576 14492 8628 14544
rect 11980 14492 12032 14544
rect 5908 14424 5960 14476
rect 8208 14424 8260 14476
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 13912 14424 13964 14476
rect 5908 14288 5960 14340
rect 6552 14331 6604 14340
rect 6552 14297 6561 14331
rect 6561 14297 6595 14331
rect 6595 14297 6604 14331
rect 6552 14288 6604 14297
rect 7564 14288 7616 14340
rect 9312 14331 9364 14340
rect 9312 14297 9321 14331
rect 9321 14297 9355 14331
rect 9355 14297 9364 14331
rect 9312 14288 9364 14297
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 7472 14220 7524 14272
rect 12164 14220 12216 14272
rect 12440 14356 12492 14408
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 13268 14356 13320 14408
rect 15936 14424 15988 14476
rect 14004 14288 14056 14340
rect 15200 14399 15252 14408
rect 15200 14365 15209 14399
rect 15209 14365 15243 14399
rect 15243 14365 15252 14399
rect 15200 14356 15252 14365
rect 15476 14356 15528 14408
rect 18696 14560 18748 14612
rect 19340 14560 19392 14612
rect 20168 14560 20220 14612
rect 21272 14560 21324 14612
rect 22560 14560 22612 14612
rect 25136 14560 25188 14612
rect 26792 14560 26844 14612
rect 28908 14603 28960 14612
rect 28908 14569 28917 14603
rect 28917 14569 28951 14603
rect 28951 14569 28960 14603
rect 28908 14560 28960 14569
rect 38016 14560 38068 14612
rect 22376 14492 22428 14544
rect 23756 14492 23808 14544
rect 27344 14492 27396 14544
rect 29736 14492 29788 14544
rect 16856 14424 16908 14476
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 17132 14399 17184 14408
rect 16580 14356 16632 14365
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 17960 14331 18012 14340
rect 17960 14297 17969 14331
rect 17969 14297 18003 14331
rect 18003 14297 18012 14331
rect 19340 14356 19392 14408
rect 22192 14424 22244 14476
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 24860 14424 24912 14476
rect 26240 14424 26292 14476
rect 27252 14424 27304 14476
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 23756 14356 23808 14365
rect 24492 14356 24544 14408
rect 27160 14356 27212 14408
rect 18880 14331 18932 14340
rect 17960 14288 18012 14297
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 15844 14220 15896 14272
rect 16028 14220 16080 14272
rect 16304 14220 16356 14272
rect 18880 14297 18889 14331
rect 18889 14297 18923 14331
rect 18923 14297 18932 14331
rect 18880 14288 18932 14297
rect 19248 14288 19300 14340
rect 18696 14220 18748 14272
rect 19524 14220 19576 14272
rect 22468 14288 22520 14340
rect 19984 14220 20036 14272
rect 21732 14220 21784 14272
rect 27344 14288 27396 14340
rect 27620 14356 27672 14408
rect 33048 14356 33100 14408
rect 37556 14399 37608 14408
rect 37556 14365 37565 14399
rect 37565 14365 37599 14399
rect 37599 14365 37608 14399
rect 37556 14356 37608 14365
rect 37924 14356 37976 14408
rect 29368 14288 29420 14340
rect 29828 14288 29880 14340
rect 30196 14331 30248 14340
rect 30196 14297 30205 14331
rect 30205 14297 30239 14331
rect 30239 14297 30248 14331
rect 30196 14288 30248 14297
rect 31484 14288 31536 14340
rect 27620 14220 27672 14272
rect 30656 14220 30708 14272
rect 37464 14220 37516 14272
rect 37924 14220 37976 14272
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 7380 14016 7432 14068
rect 8300 14016 8352 14068
rect 8392 14016 8444 14068
rect 5448 13880 5500 13932
rect 7012 13880 7064 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 10048 14016 10100 14068
rect 11888 14016 11940 14068
rect 9496 13991 9548 14000
rect 9496 13957 9505 13991
rect 9505 13957 9539 13991
rect 9539 13957 9548 13991
rect 9496 13948 9548 13957
rect 10416 13948 10468 14000
rect 15292 14016 15344 14068
rect 18696 14016 18748 14068
rect 18880 14016 18932 14068
rect 19156 14016 19208 14068
rect 21364 14016 21416 14068
rect 21548 14016 21600 14068
rect 22284 14016 22336 14068
rect 23756 14016 23808 14068
rect 23940 14016 23992 14068
rect 13360 13991 13412 14000
rect 13360 13957 13369 13991
rect 13369 13957 13403 13991
rect 13403 13957 13412 13991
rect 13360 13948 13412 13957
rect 13820 13948 13872 14000
rect 15108 13948 15160 14000
rect 8668 13744 8720 13796
rect 9220 13812 9272 13864
rect 9588 13812 9640 13864
rect 12992 13880 13044 13932
rect 12348 13855 12400 13864
rect 12348 13821 12357 13855
rect 12357 13821 12391 13855
rect 12391 13821 12400 13855
rect 12348 13812 12400 13821
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 12532 13744 12584 13796
rect 14832 13812 14884 13864
rect 17408 13948 17460 14000
rect 17684 13948 17736 14000
rect 18788 13948 18840 14000
rect 19340 13948 19392 14000
rect 20720 13948 20772 14000
rect 27712 14016 27764 14068
rect 28448 14016 28500 14068
rect 30196 14016 30248 14068
rect 27988 13948 28040 14000
rect 16488 13880 16540 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 19616 13880 19668 13932
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 29092 13880 29144 13932
rect 30564 13923 30616 13932
rect 30564 13889 30573 13923
rect 30573 13889 30607 13923
rect 30607 13889 30616 13923
rect 30564 13880 30616 13889
rect 30932 13880 30984 13932
rect 18420 13812 18472 13864
rect 19340 13812 19392 13864
rect 19432 13812 19484 13864
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 22100 13855 22152 13864
rect 22100 13821 22109 13855
rect 22109 13821 22143 13855
rect 22143 13821 22152 13855
rect 22100 13812 22152 13821
rect 7288 13676 7340 13728
rect 11612 13676 11664 13728
rect 14464 13676 14516 13728
rect 15200 13676 15252 13728
rect 15936 13676 15988 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 18236 13744 18288 13796
rect 18696 13744 18748 13796
rect 21180 13744 21232 13796
rect 22008 13744 22060 13796
rect 26700 13812 26752 13864
rect 27160 13855 27212 13864
rect 26240 13744 26292 13796
rect 27160 13821 27169 13855
rect 27169 13821 27203 13855
rect 27203 13821 27212 13855
rect 27160 13812 27212 13821
rect 26976 13744 27028 13796
rect 27528 13812 27580 13864
rect 28448 13812 28500 13864
rect 28908 13744 28960 13796
rect 29092 13744 29144 13796
rect 25136 13719 25188 13728
rect 25136 13685 25166 13719
rect 25166 13685 25188 13719
rect 25136 13676 25188 13685
rect 25504 13676 25556 13728
rect 30564 13744 30616 13796
rect 30840 13744 30892 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2044 13404 2096 13456
rect 5540 13404 5592 13456
rect 8392 13336 8444 13388
rect 9312 13472 9364 13524
rect 9496 13472 9548 13524
rect 10140 13472 10192 13524
rect 12532 13472 12584 13524
rect 15384 13472 15436 13524
rect 13360 13404 13412 13456
rect 12992 13336 13044 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 5172 13268 5224 13320
rect 7196 13268 7248 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 10048 13268 10100 13320
rect 10876 13268 10928 13320
rect 16212 13336 16264 13388
rect 16856 13336 16908 13388
rect 17776 13336 17828 13388
rect 18052 13472 18104 13524
rect 18512 13472 18564 13524
rect 20720 13472 20772 13524
rect 13636 13268 13688 13320
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15476 13268 15528 13320
rect 19616 13268 19668 13320
rect 20260 13268 20312 13320
rect 20536 13268 20588 13320
rect 21272 13472 21324 13524
rect 22376 13472 22428 13524
rect 23204 13472 23256 13524
rect 22928 13404 22980 13456
rect 24492 13404 24544 13456
rect 20904 13336 20956 13388
rect 8576 13243 8628 13252
rect 3976 13132 4028 13184
rect 8576 13209 8585 13243
rect 8585 13209 8619 13243
rect 8619 13209 8628 13243
rect 8576 13200 8628 13209
rect 14280 13200 14332 13252
rect 16488 13200 16540 13252
rect 17224 13200 17276 13252
rect 21180 13268 21232 13320
rect 22192 13336 22244 13388
rect 22652 13336 22704 13388
rect 23388 13379 23440 13388
rect 23388 13345 23397 13379
rect 23397 13345 23431 13379
rect 23431 13345 23440 13379
rect 23388 13336 23440 13345
rect 24768 13379 24820 13388
rect 24768 13345 24777 13379
rect 24777 13345 24811 13379
rect 24811 13345 24820 13379
rect 24768 13336 24820 13345
rect 37556 13472 37608 13524
rect 26332 13404 26384 13456
rect 26884 13404 26936 13456
rect 27712 13404 27764 13456
rect 27896 13404 27948 13456
rect 27160 13336 27212 13388
rect 23480 13268 23532 13320
rect 28080 13268 28132 13320
rect 33876 13268 33928 13320
rect 38292 13311 38344 13320
rect 38292 13277 38301 13311
rect 38301 13277 38335 13311
rect 38335 13277 38344 13311
rect 38292 13268 38344 13277
rect 16212 13132 16264 13184
rect 17776 13132 17828 13184
rect 19984 13132 20036 13184
rect 20536 13132 20588 13184
rect 20812 13175 20864 13184
rect 20812 13141 20821 13175
rect 20821 13141 20855 13175
rect 20855 13141 20864 13175
rect 20812 13132 20864 13141
rect 24952 13200 25004 13252
rect 25044 13243 25096 13252
rect 25044 13209 25053 13243
rect 25053 13209 25087 13243
rect 25087 13209 25096 13243
rect 25044 13200 25096 13209
rect 26516 13200 26568 13252
rect 26976 13200 27028 13252
rect 27896 13200 27948 13252
rect 28816 13200 28868 13252
rect 30012 13200 30064 13252
rect 23204 13132 23256 13184
rect 23940 13175 23992 13184
rect 23940 13141 23949 13175
rect 23949 13141 23983 13175
rect 23983 13141 23992 13175
rect 23940 13132 23992 13141
rect 24492 13132 24544 13184
rect 29552 13132 29604 13184
rect 30288 13132 30340 13184
rect 35992 13132 36044 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 9220 12928 9272 12980
rect 1952 12860 2004 12912
rect 7288 12860 7340 12912
rect 8852 12860 8904 12912
rect 9036 12860 9088 12912
rect 10140 12860 10192 12912
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 3884 12724 3936 12776
rect 7104 12656 7156 12708
rect 9128 12792 9180 12844
rect 11704 12835 11756 12844
rect 8392 12724 8444 12776
rect 7380 12656 7432 12708
rect 8024 12656 8076 12708
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12532 12928 12584 12980
rect 13084 12928 13136 12980
rect 14004 12860 14056 12912
rect 14464 12903 14516 12912
rect 14464 12869 14473 12903
rect 14473 12869 14507 12903
rect 14507 12869 14516 12903
rect 14464 12860 14516 12869
rect 15936 12928 15988 12980
rect 17776 12903 17828 12912
rect 17776 12869 17785 12903
rect 17785 12869 17819 12903
rect 17819 12869 17828 12903
rect 17776 12860 17828 12869
rect 18328 12860 18380 12912
rect 13084 12724 13136 12776
rect 14464 12724 14516 12776
rect 16856 12792 16908 12844
rect 20260 12928 20312 12980
rect 21088 12860 21140 12912
rect 23940 12860 23992 12912
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 24400 12792 24452 12844
rect 27988 12928 28040 12980
rect 28264 12928 28316 12980
rect 34520 12928 34572 12980
rect 28816 12792 28868 12844
rect 30288 12792 30340 12844
rect 33140 12792 33192 12844
rect 34796 12792 34848 12844
rect 38108 12835 38160 12844
rect 38108 12801 38117 12835
rect 38117 12801 38151 12835
rect 38151 12801 38160 12835
rect 38108 12792 38160 12801
rect 19708 12724 19760 12776
rect 21180 12724 21232 12776
rect 22376 12724 22428 12776
rect 3792 12631 3844 12640
rect 3792 12597 3801 12631
rect 3801 12597 3835 12631
rect 3835 12597 3844 12631
rect 3792 12588 3844 12597
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 6736 12588 6788 12640
rect 9404 12588 9456 12640
rect 9588 12588 9640 12640
rect 9956 12588 10008 12640
rect 17408 12656 17460 12708
rect 19156 12656 19208 12708
rect 21548 12656 21600 12708
rect 24216 12724 24268 12776
rect 34152 12724 34204 12776
rect 32404 12656 32456 12708
rect 15936 12588 15988 12640
rect 19340 12588 19392 12640
rect 19708 12588 19760 12640
rect 21916 12588 21968 12640
rect 24952 12588 25004 12640
rect 25596 12588 25648 12640
rect 27344 12588 27396 12640
rect 29092 12588 29144 12640
rect 38016 12588 38068 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5080 12427 5132 12436
rect 5080 12393 5089 12427
rect 5089 12393 5123 12427
rect 5123 12393 5132 12427
rect 5080 12384 5132 12393
rect 6000 12384 6052 12436
rect 7012 12316 7064 12368
rect 10232 12384 10284 12436
rect 11336 12384 11388 12436
rect 11980 12384 12032 12436
rect 17960 12384 18012 12436
rect 19432 12384 19484 12436
rect 19616 12384 19668 12436
rect 6000 12248 6052 12300
rect 5448 12180 5500 12232
rect 7196 12180 7248 12232
rect 9588 12248 9640 12300
rect 9680 12248 9732 12300
rect 19984 12316 20036 12368
rect 10048 12248 10100 12300
rect 10508 12248 10560 12300
rect 12532 12248 12584 12300
rect 12716 12248 12768 12300
rect 12992 12248 13044 12300
rect 13636 12248 13688 12300
rect 15200 12248 15252 12300
rect 17868 12248 17920 12300
rect 19432 12248 19484 12300
rect 21180 12384 21232 12436
rect 22560 12384 22612 12436
rect 23112 12316 23164 12368
rect 26424 12384 26476 12436
rect 26976 12384 27028 12436
rect 28632 12427 28684 12436
rect 28632 12393 28641 12427
rect 28641 12393 28675 12427
rect 28675 12393 28684 12427
rect 28632 12384 28684 12393
rect 31024 12384 31076 12436
rect 34796 12384 34848 12436
rect 8484 12180 8536 12232
rect 11520 12180 11572 12232
rect 17408 12180 17460 12232
rect 22652 12180 22704 12232
rect 25596 12316 25648 12368
rect 30564 12316 30616 12368
rect 31576 12316 31628 12368
rect 24492 12248 24544 12300
rect 25504 12248 25556 12300
rect 27160 12248 27212 12300
rect 27344 12248 27396 12300
rect 28356 12180 28408 12232
rect 5724 12112 5776 12164
rect 11704 12112 11756 12164
rect 11980 12155 12032 12164
rect 11980 12121 11989 12155
rect 11989 12121 12023 12155
rect 12023 12121 12032 12155
rect 11980 12112 12032 12121
rect 12440 12112 12492 12164
rect 7564 12044 7616 12096
rect 8300 12044 8352 12096
rect 8392 12044 8444 12096
rect 9772 12044 9824 12096
rect 15660 12112 15712 12164
rect 16212 12112 16264 12164
rect 17132 12112 17184 12164
rect 20444 12155 20496 12164
rect 20444 12121 20453 12155
rect 20453 12121 20487 12155
rect 20487 12121 20496 12155
rect 20444 12112 20496 12121
rect 18328 12044 18380 12096
rect 18880 12044 18932 12096
rect 22468 12112 22520 12164
rect 23112 12112 23164 12164
rect 25504 12112 25556 12164
rect 25964 12155 26016 12164
rect 25964 12121 25973 12155
rect 25973 12121 26007 12155
rect 26007 12121 26016 12155
rect 25964 12112 26016 12121
rect 26332 12044 26384 12096
rect 28908 12112 28960 12164
rect 29736 12044 29788 12096
rect 30472 12044 30524 12096
rect 33508 12112 33560 12164
rect 31760 12044 31812 12096
rect 32128 12044 32180 12096
rect 32680 12044 32732 12096
rect 37372 12180 37424 12232
rect 37004 12112 37056 12164
rect 36176 12044 36228 12096
rect 39028 12044 39080 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 9772 11840 9824 11892
rect 6276 11772 6328 11824
rect 7380 11772 7432 11824
rect 8392 11815 8444 11824
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 7196 11704 7248 11756
rect 8392 11781 8401 11815
rect 8401 11781 8435 11815
rect 8435 11781 8444 11815
rect 8392 11772 8444 11781
rect 7748 11704 7800 11756
rect 4620 11636 4672 11688
rect 5816 11636 5868 11688
rect 6552 11636 6604 11688
rect 6828 11568 6880 11620
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 2320 11500 2372 11509
rect 3240 11500 3292 11552
rect 7196 11500 7248 11552
rect 8392 11636 8444 11688
rect 8484 11636 8536 11688
rect 9680 11772 9732 11824
rect 10140 11840 10192 11892
rect 10232 11840 10284 11892
rect 15660 11840 15712 11892
rect 18236 11840 18288 11892
rect 10784 11772 10836 11824
rect 12072 11772 12124 11824
rect 14740 11772 14792 11824
rect 14832 11772 14884 11824
rect 19432 11840 19484 11892
rect 20444 11840 20496 11892
rect 26976 11840 27028 11892
rect 18512 11772 18564 11824
rect 19064 11772 19116 11824
rect 20260 11772 20312 11824
rect 23756 11815 23808 11824
rect 23756 11781 23765 11815
rect 23765 11781 23799 11815
rect 23799 11781 23808 11815
rect 23756 11772 23808 11781
rect 26056 11772 26108 11824
rect 9312 11568 9364 11620
rect 9680 11568 9732 11620
rect 10048 11636 10100 11688
rect 22100 11704 22152 11756
rect 25504 11704 25556 11756
rect 31208 11840 31260 11892
rect 31668 11840 31720 11892
rect 32588 11883 32640 11892
rect 32588 11849 32597 11883
rect 32597 11849 32631 11883
rect 32631 11849 32640 11883
rect 32588 11840 32640 11849
rect 27344 11772 27396 11824
rect 27712 11772 27764 11824
rect 30656 11772 30708 11824
rect 30012 11704 30064 11756
rect 32680 11772 32732 11824
rect 31392 11704 31444 11756
rect 12348 11679 12400 11688
rect 12348 11645 12357 11679
rect 12357 11645 12391 11679
rect 12391 11645 12400 11679
rect 12348 11636 12400 11645
rect 12624 11679 12676 11688
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 13268 11636 13320 11688
rect 10140 11568 10192 11620
rect 10692 11568 10744 11620
rect 11060 11568 11112 11620
rect 12072 11500 12124 11552
rect 13912 11500 13964 11552
rect 14004 11500 14056 11552
rect 14280 11500 14332 11552
rect 17960 11636 18012 11688
rect 21272 11636 21324 11688
rect 21364 11636 21416 11688
rect 27160 11679 27212 11688
rect 15200 11500 15252 11552
rect 15844 11500 15896 11552
rect 16672 11500 16724 11552
rect 18696 11500 18748 11552
rect 19708 11500 19760 11552
rect 24308 11500 24360 11552
rect 27160 11645 27169 11679
rect 27169 11645 27203 11679
rect 27203 11645 27212 11679
rect 27160 11636 27212 11645
rect 26424 11568 26476 11620
rect 27068 11568 27120 11620
rect 29184 11679 29236 11688
rect 29184 11645 29193 11679
rect 29193 11645 29227 11679
rect 29227 11645 29236 11679
rect 29184 11636 29236 11645
rect 30656 11636 30708 11688
rect 32312 11636 32364 11688
rect 35348 11772 35400 11824
rect 36084 11747 36136 11756
rect 36084 11713 36093 11747
rect 36093 11713 36127 11747
rect 36127 11713 36136 11747
rect 36084 11704 36136 11713
rect 29736 11568 29788 11620
rect 30012 11568 30064 11620
rect 37280 11704 37332 11756
rect 38936 11568 38988 11620
rect 30104 11500 30156 11552
rect 30840 11500 30892 11552
rect 38108 11500 38160 11552
rect 38292 11500 38344 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3148 11296 3200 11348
rect 7288 11296 7340 11348
rect 7656 11296 7708 11348
rect 1032 11228 1084 11280
rect 4988 11160 5040 11212
rect 5172 11160 5224 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 4068 11092 4120 11144
rect 4896 11024 4948 11076
rect 1768 10999 1820 11008
rect 1768 10965 1777 10999
rect 1777 10965 1811 10999
rect 1811 10965 1820 10999
rect 1768 10956 1820 10965
rect 4620 10956 4672 11008
rect 5080 11024 5132 11076
rect 6092 11092 6144 11144
rect 6460 11092 6512 11144
rect 7380 11228 7432 11280
rect 7748 11228 7800 11280
rect 10048 11296 10100 11348
rect 10140 11296 10192 11348
rect 11244 11296 11296 11348
rect 11704 11296 11756 11348
rect 7656 11160 7708 11212
rect 7840 11203 7892 11212
rect 7840 11169 7849 11203
rect 7849 11169 7883 11203
rect 7883 11169 7892 11203
rect 7840 11160 7892 11169
rect 12440 11296 12492 11348
rect 14096 11296 14148 11348
rect 15476 11296 15528 11348
rect 18144 11296 18196 11348
rect 17132 11228 17184 11280
rect 23112 11296 23164 11348
rect 25136 11296 25188 11348
rect 23756 11228 23808 11280
rect 37464 11271 37516 11280
rect 37464 11237 37473 11271
rect 37473 11237 37507 11271
rect 37507 11237 37516 11271
rect 37464 11228 37516 11237
rect 38660 11228 38712 11280
rect 14004 11160 14056 11212
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15476 11203 15528 11212
rect 15200 11160 15252 11169
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 20260 11160 20312 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 14280 11135 14332 11144
rect 14280 11101 14281 11135
rect 14281 11101 14315 11135
rect 14315 11101 14332 11135
rect 14280 11092 14332 11101
rect 15108 11092 15160 11144
rect 5908 11024 5960 11076
rect 7564 11067 7616 11076
rect 7564 11033 7573 11067
rect 7573 11033 7607 11067
rect 7607 11033 7616 11067
rect 7564 11024 7616 11033
rect 10140 11024 10192 11076
rect 11336 11024 11388 11076
rect 12256 11024 12308 11076
rect 14924 11024 14976 11076
rect 6000 10956 6052 11008
rect 8484 10956 8536 11008
rect 9864 10956 9916 11008
rect 13636 10956 13688 11008
rect 20720 11024 20772 11076
rect 22008 11160 22060 11212
rect 22100 11160 22152 11212
rect 22652 11160 22704 11212
rect 26240 11203 26292 11212
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 29368 11160 29420 11212
rect 29552 11160 29604 11212
rect 30288 11160 30340 11212
rect 24584 11092 24636 11144
rect 24676 11092 24728 11144
rect 18696 10956 18748 11008
rect 18880 10956 18932 11008
rect 24768 11024 24820 11076
rect 29092 11092 29144 11144
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30564 11160 30616 11212
rect 30932 11160 30984 11212
rect 30472 11092 30524 11144
rect 31576 11160 31628 11212
rect 36268 11160 36320 11212
rect 38108 11160 38160 11212
rect 31944 11092 31996 11144
rect 35900 11092 35952 11144
rect 37372 11135 37424 11144
rect 37372 11101 37381 11135
rect 37381 11101 37415 11135
rect 37415 11101 37424 11135
rect 37372 11092 37424 11101
rect 38660 11092 38712 11144
rect 31760 11067 31812 11076
rect 31760 11033 31769 11067
rect 31769 11033 31803 11067
rect 31803 11033 31812 11067
rect 32588 11067 32640 11076
rect 31760 11024 31812 11033
rect 32588 11033 32597 11067
rect 32597 11033 32631 11067
rect 32631 11033 32640 11067
rect 32588 11024 32640 11033
rect 34060 11024 34112 11076
rect 36544 11024 36596 11076
rect 38108 11067 38160 11076
rect 38108 11033 38117 11067
rect 38117 11033 38151 11067
rect 38151 11033 38160 11067
rect 38108 11024 38160 11033
rect 24400 10956 24452 11008
rect 26332 10956 26384 11008
rect 26792 10956 26844 11008
rect 29092 10956 29144 11008
rect 29736 10999 29788 11008
rect 29736 10965 29745 10999
rect 29745 10965 29779 10999
rect 29779 10965 29788 10999
rect 29736 10956 29788 10965
rect 31116 10999 31168 11008
rect 31116 10965 31125 10999
rect 31125 10965 31159 10999
rect 31159 10965 31168 10999
rect 31116 10956 31168 10965
rect 32772 10956 32824 11008
rect 36084 10956 36136 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 2780 10616 2832 10668
rect 3332 10684 3384 10736
rect 5816 10752 5868 10804
rect 7656 10752 7708 10804
rect 5632 10684 5684 10736
rect 7196 10727 7248 10736
rect 7196 10693 7205 10727
rect 7205 10693 7239 10727
rect 7239 10693 7248 10727
rect 7196 10684 7248 10693
rect 7288 10684 7340 10736
rect 8300 10684 8352 10736
rect 9404 10752 9456 10804
rect 10784 10752 10836 10804
rect 11980 10752 12032 10804
rect 14280 10752 14332 10804
rect 17132 10752 17184 10804
rect 17868 10752 17920 10804
rect 21088 10752 21140 10804
rect 24400 10752 24452 10804
rect 9956 10727 10008 10736
rect 9956 10693 9965 10727
rect 9965 10693 9999 10727
rect 9999 10693 10008 10727
rect 9956 10684 10008 10693
rect 2964 10616 3016 10668
rect 4620 10616 4672 10668
rect 5540 10616 5592 10668
rect 12624 10684 12676 10736
rect 14464 10727 14516 10736
rect 14464 10693 14473 10727
rect 14473 10693 14507 10727
rect 14507 10693 14516 10727
rect 14464 10684 14516 10693
rect 12440 10625 12449 10652
rect 12449 10625 12483 10652
rect 12483 10625 12492 10652
rect 12440 10600 12492 10625
rect 13820 10616 13872 10668
rect 14372 10616 14424 10668
rect 16488 10616 16540 10668
rect 20812 10684 20864 10736
rect 29184 10752 29236 10804
rect 24952 10684 25004 10736
rect 25964 10684 26016 10736
rect 26792 10684 26844 10736
rect 29460 10727 29512 10736
rect 29460 10693 29469 10727
rect 29469 10693 29503 10727
rect 29503 10693 29512 10727
rect 29460 10684 29512 10693
rect 32404 10752 32456 10804
rect 32588 10795 32640 10804
rect 32588 10761 32597 10795
rect 32597 10761 32631 10795
rect 32631 10761 32640 10795
rect 32588 10752 32640 10761
rect 29920 10684 29972 10736
rect 30104 10684 30156 10736
rect 30288 10684 30340 10736
rect 6920 10548 6972 10600
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 8392 10548 8444 10600
rect 9680 10548 9732 10600
rect 9956 10548 10008 10600
rect 10232 10548 10284 10600
rect 13176 10548 13228 10600
rect 13452 10548 13504 10600
rect 3332 10480 3384 10532
rect 2504 10412 2556 10464
rect 3424 10412 3476 10464
rect 3608 10455 3660 10464
rect 3608 10421 3617 10455
rect 3617 10421 3651 10455
rect 3651 10421 3660 10455
rect 3608 10412 3660 10421
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 5816 10412 5868 10464
rect 7380 10412 7432 10464
rect 9588 10412 9640 10464
rect 15660 10455 15712 10464
rect 15660 10421 15669 10455
rect 15669 10421 15703 10455
rect 15703 10421 15712 10455
rect 15660 10412 15712 10421
rect 18328 10548 18380 10600
rect 18420 10548 18472 10600
rect 18788 10480 18840 10532
rect 22560 10480 22612 10532
rect 17868 10412 17920 10464
rect 18052 10412 18104 10464
rect 18328 10412 18380 10464
rect 19892 10412 19944 10464
rect 21916 10412 21968 10464
rect 25044 10548 25096 10600
rect 27160 10591 27212 10600
rect 27160 10557 27169 10591
rect 27169 10557 27203 10591
rect 27203 10557 27212 10591
rect 27160 10548 27212 10557
rect 28080 10548 28132 10600
rect 30380 10548 30432 10600
rect 30748 10684 30800 10736
rect 30748 10548 30800 10600
rect 26056 10480 26108 10532
rect 26332 10412 26384 10464
rect 29000 10412 29052 10464
rect 30288 10480 30340 10532
rect 32036 10616 32088 10668
rect 33140 10616 33192 10668
rect 38752 10684 38804 10736
rect 35624 10616 35676 10668
rect 36728 10659 36780 10668
rect 36728 10625 36737 10659
rect 36737 10625 36771 10659
rect 36771 10625 36780 10659
rect 36728 10616 36780 10625
rect 38108 10659 38160 10668
rect 38108 10625 38117 10659
rect 38117 10625 38151 10659
rect 38151 10625 38160 10659
rect 38108 10616 38160 10625
rect 31668 10548 31720 10600
rect 31208 10412 31260 10464
rect 33416 10412 33468 10464
rect 35532 10412 35584 10464
rect 35900 10412 35952 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2964 10208 3016 10260
rect 6276 10251 6328 10260
rect 6276 10217 6285 10251
rect 6285 10217 6319 10251
rect 6319 10217 6328 10251
rect 6276 10208 6328 10217
rect 7472 10208 7524 10260
rect 1492 10140 1544 10192
rect 7104 10140 7156 10192
rect 11980 10208 12032 10260
rect 12348 10208 12400 10260
rect 15660 10208 15712 10260
rect 2596 10072 2648 10124
rect 7564 10115 7616 10124
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 2136 10004 2188 10056
rect 2504 10004 2556 10056
rect 2872 10004 2924 10056
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 9864 10072 9916 10124
rect 4988 10004 5040 10056
rect 5356 10004 5408 10056
rect 5816 10004 5868 10056
rect 6276 10004 6328 10056
rect 7196 10004 7248 10056
rect 9404 10004 9456 10056
rect 11520 10004 11572 10056
rect 14556 10072 14608 10124
rect 16396 10072 16448 10124
rect 18420 10072 18472 10124
rect 13084 10004 13136 10056
rect 13268 10004 13320 10056
rect 16856 10004 16908 10056
rect 24124 10208 24176 10260
rect 25044 10208 25096 10260
rect 31208 10208 31260 10260
rect 32220 10208 32272 10260
rect 32496 10208 32548 10260
rect 33600 10208 33652 10260
rect 37556 10208 37608 10260
rect 37924 10208 37976 10260
rect 18880 10183 18932 10192
rect 18880 10149 18889 10183
rect 18889 10149 18923 10183
rect 18923 10149 18932 10183
rect 18880 10140 18932 10149
rect 26976 10140 27028 10192
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 22744 10072 22796 10124
rect 26332 10072 26384 10124
rect 27620 10140 27672 10192
rect 31484 10140 31536 10192
rect 31944 10140 31996 10192
rect 29828 10072 29880 10124
rect 31116 10072 31168 10124
rect 20444 10004 20496 10056
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 27160 10004 27212 10056
rect 34520 10140 34572 10192
rect 36268 10072 36320 10124
rect 6644 9936 6696 9988
rect 7656 9979 7708 9988
rect 7656 9945 7665 9979
rect 7665 9945 7699 9979
rect 7699 9945 7708 9979
rect 11980 9979 12032 9988
rect 7656 9936 7708 9945
rect 2412 9868 2464 9920
rect 4804 9868 4856 9920
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 11244 9911 11296 9920
rect 11244 9877 11253 9911
rect 11253 9877 11287 9911
rect 11287 9877 11296 9911
rect 11244 9868 11296 9877
rect 11980 9945 11989 9979
rect 11989 9945 12023 9979
rect 12023 9945 12032 9979
rect 11980 9936 12032 9945
rect 12256 9936 12308 9988
rect 14648 9868 14700 9920
rect 15292 9936 15344 9988
rect 25688 9936 25740 9988
rect 26056 9936 26108 9988
rect 27436 9936 27488 9988
rect 27896 9936 27948 9988
rect 32036 10004 32088 10056
rect 33324 10004 33376 10056
rect 33692 10004 33744 10056
rect 34152 10047 34204 10056
rect 34152 10013 34161 10047
rect 34161 10013 34195 10047
rect 34195 10013 34204 10047
rect 34152 10004 34204 10013
rect 19892 9868 19944 9920
rect 20260 9868 20312 9920
rect 26700 9868 26752 9920
rect 31576 9936 31628 9988
rect 32588 9936 32640 9988
rect 29828 9868 29880 9920
rect 33784 9868 33836 9920
rect 34612 9868 34664 9920
rect 35440 10004 35492 10056
rect 36912 10047 36964 10056
rect 36912 10013 36921 10047
rect 36921 10013 36955 10047
rect 36955 10013 36964 10047
rect 36912 10004 36964 10013
rect 37372 10047 37424 10056
rect 37372 10013 37381 10047
rect 37381 10013 37415 10047
rect 37415 10013 37424 10047
rect 37372 10004 37424 10013
rect 38384 10004 38436 10056
rect 35808 9936 35860 9988
rect 36636 9868 36688 9920
rect 38108 9868 38160 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 1308 9664 1360 9716
rect 5540 9664 5592 9716
rect 6920 9664 6972 9716
rect 1400 9528 1452 9580
rect 5908 9596 5960 9648
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 7748 9596 7800 9648
rect 8024 9639 8076 9648
rect 8024 9605 8033 9639
rect 8033 9605 8067 9639
rect 8067 9605 8076 9639
rect 8024 9596 8076 9605
rect 8760 9596 8812 9648
rect 9128 9596 9180 9648
rect 10968 9596 11020 9648
rect 11612 9596 11664 9648
rect 12532 9596 12584 9648
rect 13636 9596 13688 9648
rect 14832 9639 14884 9648
rect 14832 9605 14841 9639
rect 14841 9605 14875 9639
rect 14875 9605 14884 9639
rect 14832 9596 14884 9605
rect 16120 9596 16172 9648
rect 20996 9639 21048 9648
rect 20996 9605 21005 9639
rect 21005 9605 21039 9639
rect 21039 9605 21048 9639
rect 20996 9596 21048 9605
rect 22376 9596 22428 9648
rect 22836 9596 22888 9648
rect 24768 9596 24820 9648
rect 27712 9596 27764 9648
rect 28448 9664 28500 9716
rect 29092 9664 29144 9716
rect 34152 9664 34204 9716
rect 36636 9664 36688 9716
rect 37096 9664 37148 9716
rect 30288 9639 30340 9648
rect 30288 9605 30297 9639
rect 30297 9605 30331 9639
rect 30331 9605 30340 9639
rect 30288 9596 30340 9605
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 2228 9460 2280 9512
rect 4620 9528 4672 9580
rect 4712 9528 4764 9580
rect 5448 9528 5500 9580
rect 5540 9528 5592 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 16580 9528 16632 9580
rect 17132 9528 17184 9580
rect 4896 9460 4948 9512
rect 5908 9460 5960 9512
rect 6828 9460 6880 9512
rect 7932 9503 7984 9512
rect 3884 9392 3936 9444
rect 4068 9392 4120 9444
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 5448 9324 5500 9376
rect 6736 9324 6788 9376
rect 6920 9392 6972 9444
rect 7288 9392 7340 9444
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 11704 9503 11756 9512
rect 8760 9392 8812 9444
rect 11704 9469 11713 9503
rect 11713 9469 11747 9503
rect 11747 9469 11756 9503
rect 11704 9460 11756 9469
rect 12440 9460 12492 9512
rect 14280 9460 14332 9512
rect 15844 9460 15896 9512
rect 16212 9460 16264 9512
rect 16488 9460 16540 9512
rect 17592 9460 17644 9512
rect 16764 9392 16816 9444
rect 10968 9324 11020 9376
rect 13176 9324 13228 9376
rect 14924 9324 14976 9376
rect 17316 9324 17368 9376
rect 18420 9528 18472 9580
rect 18880 9528 18932 9580
rect 20352 9528 20404 9580
rect 20812 9528 20864 9580
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 26976 9528 27028 9580
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 18236 9460 18288 9512
rect 18512 9460 18564 9512
rect 19248 9460 19300 9512
rect 21456 9460 21508 9512
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 18880 9324 18932 9376
rect 19340 9324 19392 9376
rect 19616 9324 19668 9376
rect 22652 9460 22704 9512
rect 24676 9460 24728 9512
rect 25136 9503 25188 9512
rect 22284 9324 22336 9376
rect 24768 9324 24820 9376
rect 25136 9469 25145 9503
rect 25145 9469 25179 9503
rect 25179 9469 25188 9503
rect 25136 9460 25188 9469
rect 26148 9460 26200 9512
rect 29552 9528 29604 9580
rect 34520 9596 34572 9648
rect 33048 9528 33100 9580
rect 33140 9528 33192 9580
rect 34152 9528 34204 9580
rect 34244 9571 34296 9580
rect 34244 9537 34253 9571
rect 34253 9537 34287 9571
rect 34287 9537 34296 9571
rect 34244 9528 34296 9537
rect 34428 9528 34480 9580
rect 35808 9571 35860 9580
rect 35808 9537 35817 9571
rect 35817 9537 35851 9571
rect 35851 9537 35860 9571
rect 35808 9528 35860 9537
rect 36452 9571 36504 9580
rect 36452 9537 36461 9571
rect 36461 9537 36495 9571
rect 36495 9537 36504 9571
rect 36452 9528 36504 9537
rect 36820 9528 36872 9580
rect 28632 9460 28684 9512
rect 26332 9324 26384 9376
rect 26976 9324 27028 9376
rect 29920 9392 29972 9444
rect 28908 9367 28960 9376
rect 28908 9333 28917 9367
rect 28917 9333 28951 9367
rect 28951 9333 28960 9367
rect 29460 9367 29512 9376
rect 28908 9324 28960 9333
rect 29460 9333 29469 9367
rect 29469 9333 29503 9367
rect 29503 9333 29512 9367
rect 29460 9324 29512 9333
rect 30288 9460 30340 9512
rect 31852 9460 31904 9512
rect 33324 9460 33376 9512
rect 30380 9392 30432 9444
rect 33692 9435 33744 9444
rect 33692 9401 33701 9435
rect 33701 9401 33735 9435
rect 33735 9401 33744 9435
rect 33692 9392 33744 9401
rect 37372 9392 37424 9444
rect 31760 9324 31812 9376
rect 32220 9324 32272 9376
rect 33140 9324 33192 9376
rect 33876 9324 33928 9376
rect 34336 9367 34388 9376
rect 34336 9333 34345 9367
rect 34345 9333 34379 9367
rect 34379 9333 34388 9367
rect 34336 9324 34388 9333
rect 34796 9324 34848 9376
rect 37464 9324 37516 9376
rect 38016 9324 38068 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3240 9120 3292 9172
rect 8208 9120 8260 9172
rect 4068 9052 4120 9104
rect 2228 8984 2280 9036
rect 7932 9052 7984 9104
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 6184 8984 6236 9036
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 6460 8984 6512 9036
rect 8116 8984 8168 9036
rect 8944 8984 8996 9036
rect 5540 8916 5592 8968
rect 6000 8916 6052 8968
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 9404 9052 9456 9104
rect 12256 9052 12308 9104
rect 14188 9052 14240 9104
rect 11796 8984 11848 9036
rect 17316 9120 17368 9172
rect 18236 9120 18288 9172
rect 19616 9120 19668 9172
rect 22100 9120 22152 9172
rect 22192 9120 22244 9172
rect 23388 9120 23440 9172
rect 26056 9120 26108 9172
rect 7012 8916 7064 8925
rect 3056 8848 3108 8900
rect 3516 8780 3568 8832
rect 3976 8848 4028 8900
rect 6368 8848 6420 8900
rect 5540 8780 5592 8832
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 7840 8848 7892 8900
rect 9036 8848 9088 8900
rect 9588 8891 9640 8900
rect 9588 8857 9597 8891
rect 9597 8857 9631 8891
rect 9631 8857 9640 8891
rect 9588 8848 9640 8857
rect 9772 8848 9824 8900
rect 9956 8848 10008 8900
rect 10876 8848 10928 8900
rect 11520 8848 11572 8900
rect 12256 8848 12308 8900
rect 8760 8780 8812 8832
rect 14556 8984 14608 9036
rect 16580 8984 16632 9036
rect 17500 8984 17552 9036
rect 17592 8984 17644 9036
rect 13360 8916 13412 8968
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 19984 8984 20036 9036
rect 20812 9027 20864 9036
rect 20812 8993 20821 9027
rect 20821 8993 20855 9027
rect 20855 8993 20864 9027
rect 20812 8984 20864 8993
rect 22100 8984 22152 9036
rect 18512 8916 18564 8968
rect 19340 8916 19392 8968
rect 24032 9052 24084 9104
rect 27804 9120 27856 9172
rect 29460 9052 29512 9104
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 23296 8984 23348 9036
rect 23020 8916 23072 8968
rect 24400 8984 24452 9036
rect 26332 8984 26384 9036
rect 26884 8984 26936 9036
rect 28172 8984 28224 9036
rect 34336 9120 34388 9172
rect 36452 9120 36504 9172
rect 37004 9163 37056 9172
rect 37004 9129 37013 9163
rect 37013 9129 37047 9163
rect 37047 9129 37056 9163
rect 37004 9120 37056 9129
rect 31116 9052 31168 9104
rect 34980 9052 35032 9104
rect 37280 9052 37332 9104
rect 29644 8984 29696 9036
rect 30288 8984 30340 9036
rect 30748 9027 30800 9036
rect 30748 8993 30757 9027
rect 30757 8993 30791 9027
rect 30791 8993 30800 9027
rect 30748 8984 30800 8993
rect 13084 8848 13136 8900
rect 13728 8848 13780 8900
rect 14556 8848 14608 8900
rect 15016 8848 15068 8900
rect 17132 8891 17184 8900
rect 17132 8857 17141 8891
rect 17141 8857 17175 8891
rect 17175 8857 17184 8891
rect 17132 8848 17184 8857
rect 19432 8891 19484 8900
rect 19432 8857 19441 8891
rect 19441 8857 19475 8891
rect 19475 8857 19484 8891
rect 19432 8848 19484 8857
rect 27344 8916 27396 8968
rect 28448 8959 28500 8968
rect 28448 8925 28457 8959
rect 28457 8925 28491 8959
rect 28491 8925 28500 8959
rect 28448 8916 28500 8925
rect 29000 8916 29052 8968
rect 24860 8848 24912 8900
rect 13176 8780 13228 8832
rect 21180 8780 21232 8832
rect 22008 8780 22060 8832
rect 23848 8780 23900 8832
rect 24952 8780 25004 8832
rect 25596 8780 25648 8832
rect 27712 8848 27764 8900
rect 31760 8984 31812 9036
rect 31852 9027 31904 9036
rect 31852 8993 31861 9027
rect 31861 8993 31895 9027
rect 31895 8993 31904 9027
rect 31852 8984 31904 8993
rect 34244 8984 34296 9036
rect 32772 8916 32824 8968
rect 33232 8959 33284 8968
rect 33232 8925 33241 8959
rect 33241 8925 33275 8959
rect 33275 8925 33284 8959
rect 33232 8916 33284 8925
rect 33508 8916 33560 8968
rect 33876 8959 33928 8968
rect 33876 8925 33885 8959
rect 33885 8925 33919 8959
rect 33919 8925 33928 8959
rect 33876 8916 33928 8925
rect 34520 8916 34572 8968
rect 35716 8959 35768 8968
rect 26884 8780 26936 8832
rect 27068 8780 27120 8832
rect 29000 8780 29052 8832
rect 30472 8780 30524 8832
rect 31668 8780 31720 8832
rect 33140 8848 33192 8900
rect 35256 8848 35308 8900
rect 34796 8780 34848 8832
rect 35716 8925 35725 8959
rect 35725 8925 35759 8959
rect 35759 8925 35768 8959
rect 35716 8916 35768 8925
rect 36544 8959 36596 8968
rect 36544 8925 36553 8959
rect 36553 8925 36587 8959
rect 36587 8925 36596 8959
rect 36544 8916 36596 8925
rect 35808 8848 35860 8900
rect 37832 8916 37884 8968
rect 37188 8780 37240 8832
rect 37832 8780 37884 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4712 8576 4764 8628
rect 5448 8551 5500 8560
rect 5448 8517 5450 8551
rect 5450 8517 5484 8551
rect 5484 8517 5500 8551
rect 5448 8508 5500 8517
rect 6828 8551 6880 8560
rect 6828 8517 6830 8551
rect 6830 8517 6864 8551
rect 6864 8517 6880 8551
rect 8116 8576 8168 8628
rect 9772 8576 9824 8628
rect 6828 8508 6880 8517
rect 8576 8508 8628 8560
rect 11244 8576 11296 8628
rect 12440 8576 12492 8628
rect 11888 8508 11940 8560
rect 12532 8508 12584 8560
rect 14280 8576 14332 8628
rect 12900 8508 12952 8560
rect 16580 8576 16632 8628
rect 16856 8576 16908 8628
rect 16304 8508 16356 8560
rect 16396 8508 16448 8560
rect 18972 8508 19024 8560
rect 19432 8576 19484 8628
rect 2596 8440 2648 8492
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 4252 8440 4304 8492
rect 2872 8372 2924 8424
rect 6368 8440 6420 8492
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 11612 8440 11664 8492
rect 11796 8440 11848 8492
rect 19340 8508 19392 8560
rect 21732 8508 21784 8560
rect 24768 8576 24820 8628
rect 32404 8619 32456 8628
rect 21916 8440 21968 8492
rect 23848 8440 23900 8492
rect 27068 8508 27120 8560
rect 27344 8508 27396 8560
rect 6828 8372 6880 8424
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 8852 8372 8904 8424
rect 1952 8304 2004 8356
rect 3240 8304 3292 8356
rect 6920 8304 6972 8356
rect 7380 8304 7432 8356
rect 7656 8304 7708 8356
rect 8208 8304 8260 8356
rect 9772 8372 9824 8424
rect 10140 8372 10192 8424
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 17132 8372 17184 8424
rect 18420 8372 18472 8424
rect 21088 8415 21140 8424
rect 14096 8347 14148 8356
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 16120 8304 16172 8356
rect 21088 8381 21097 8415
rect 21097 8381 21131 8415
rect 21131 8381 21140 8415
rect 21088 8372 21140 8381
rect 21180 8372 21232 8424
rect 22836 8372 22888 8424
rect 24952 8372 25004 8424
rect 25136 8372 25188 8424
rect 27160 8415 27212 8424
rect 25504 8304 25556 8356
rect 25780 8304 25832 8356
rect 26332 8304 26384 8356
rect 27160 8381 27169 8415
rect 27169 8381 27203 8415
rect 27203 8381 27212 8415
rect 27160 8372 27212 8381
rect 27988 8372 28040 8424
rect 29184 8440 29236 8492
rect 29368 8440 29420 8492
rect 32404 8585 32413 8619
rect 32413 8585 32447 8619
rect 32447 8585 32456 8619
rect 32404 8576 32456 8585
rect 32956 8576 33008 8628
rect 34980 8619 35032 8628
rect 32036 8508 32088 8560
rect 34980 8585 34989 8619
rect 34989 8585 35023 8619
rect 35023 8585 35032 8619
rect 34980 8576 35032 8585
rect 30380 8415 30432 8424
rect 30380 8381 30389 8415
rect 30389 8381 30423 8415
rect 30423 8381 30432 8415
rect 30380 8372 30432 8381
rect 30564 8372 30616 8424
rect 31024 8372 31076 8424
rect 31668 8372 31720 8424
rect 32680 8440 32732 8492
rect 33232 8440 33284 8492
rect 34520 8440 34572 8492
rect 35440 8440 35492 8492
rect 36268 8508 36320 8560
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 38016 8483 38068 8492
rect 38016 8449 38025 8483
rect 38025 8449 38059 8483
rect 38059 8449 38068 8483
rect 38016 8440 38068 8449
rect 35624 8372 35676 8424
rect 30932 8304 30984 8356
rect 3700 8236 3752 8288
rect 4068 8236 4120 8288
rect 6368 8236 6420 8288
rect 9680 8236 9732 8288
rect 11888 8236 11940 8288
rect 12256 8236 12308 8288
rect 14556 8236 14608 8288
rect 16764 8236 16816 8288
rect 19064 8236 19116 8288
rect 19156 8236 19208 8288
rect 19432 8236 19484 8288
rect 21088 8236 21140 8288
rect 24952 8236 25004 8288
rect 25872 8236 25924 8288
rect 26148 8236 26200 8288
rect 28724 8236 28776 8288
rect 30288 8236 30340 8288
rect 33876 8304 33928 8356
rect 34520 8304 34572 8356
rect 34888 8304 34940 8356
rect 35256 8304 35308 8356
rect 35440 8304 35492 8356
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 38200 8347 38252 8356
rect 38200 8313 38209 8347
rect 38209 8313 38243 8347
rect 38243 8313 38252 8347
rect 38200 8304 38252 8313
rect 31668 8236 31720 8288
rect 34244 8236 34296 8288
rect 34428 8236 34480 8288
rect 37004 8236 37056 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1400 8032 1452 8084
rect 1584 8032 1636 8084
rect 4712 8075 4764 8084
rect 4712 8041 4721 8075
rect 4721 8041 4755 8075
rect 4755 8041 4764 8075
rect 4712 8032 4764 8041
rect 5356 8075 5408 8084
rect 5356 8041 5365 8075
rect 5365 8041 5399 8075
rect 5399 8041 5408 8075
rect 5356 8032 5408 8041
rect 6184 8032 6236 8084
rect 15752 8032 15804 8084
rect 16948 8032 17000 8084
rect 20812 8032 20864 8084
rect 20996 8032 21048 8084
rect 24768 8032 24820 8084
rect 24860 8032 24912 8084
rect 27896 8032 27948 8084
rect 31944 8032 31996 8084
rect 32036 8032 32088 8084
rect 33140 8032 33192 8084
rect 33968 8032 34020 8084
rect 34428 8032 34480 8084
rect 34704 8032 34756 8084
rect 35624 8075 35676 8084
rect 35624 8041 35633 8075
rect 35633 8041 35667 8075
rect 35667 8041 35676 8075
rect 35624 8032 35676 8041
rect 3792 7964 3844 8016
rect 8024 7964 8076 8016
rect 11060 7964 11112 8016
rect 13084 7964 13136 8016
rect 16212 7964 16264 8016
rect 3056 7828 3108 7880
rect 4896 7828 4948 7880
rect 5448 7896 5500 7948
rect 7012 7896 7064 7948
rect 7380 7896 7432 7948
rect 7840 7896 7892 7948
rect 9220 7896 9272 7948
rect 12348 7896 12400 7948
rect 12440 7896 12492 7948
rect 13544 7896 13596 7948
rect 15292 7896 15344 7948
rect 15568 7896 15620 7948
rect 5356 7828 5408 7880
rect 9404 7828 9456 7880
rect 11336 7828 11388 7880
rect 11520 7828 11572 7880
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 13912 7828 13964 7880
rect 14648 7828 14700 7880
rect 16304 7828 16356 7880
rect 16856 7896 16908 7948
rect 18512 7964 18564 8016
rect 19340 7896 19392 7948
rect 26148 7964 26200 8016
rect 28080 7964 28132 8016
rect 28908 7964 28960 8016
rect 30932 7964 30984 8016
rect 32496 7964 32548 8016
rect 34244 7964 34296 8016
rect 20168 7896 20220 7948
rect 21180 7896 21232 7948
rect 22008 7939 22060 7948
rect 22008 7905 22017 7939
rect 22017 7905 22051 7939
rect 22051 7905 22060 7939
rect 22008 7896 22060 7905
rect 23020 7896 23072 7948
rect 17040 7828 17092 7880
rect 18512 7828 18564 7880
rect 24400 7828 24452 7880
rect 25964 7828 26016 7880
rect 26976 7896 27028 7948
rect 27160 7896 27212 7948
rect 27620 7828 27672 7880
rect 5724 7760 5776 7812
rect 5816 7760 5868 7812
rect 6092 7803 6144 7812
rect 6092 7769 6101 7803
rect 6101 7769 6135 7803
rect 6135 7769 6144 7803
rect 6092 7760 6144 7769
rect 6828 7760 6880 7812
rect 7380 7760 7432 7812
rect 8576 7803 8628 7812
rect 1768 7735 1820 7744
rect 1768 7701 1777 7735
rect 1777 7701 1811 7735
rect 1811 7701 1820 7735
rect 1768 7692 1820 7701
rect 2504 7692 2556 7744
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 4068 7692 4120 7744
rect 7196 7692 7248 7744
rect 8576 7769 8585 7803
rect 8585 7769 8619 7803
rect 8619 7769 8628 7803
rect 8576 7760 8628 7769
rect 10508 7760 10560 7812
rect 12072 7760 12124 7812
rect 12992 7760 13044 7812
rect 7840 7692 7892 7744
rect 9128 7692 9180 7744
rect 11244 7692 11296 7744
rect 11336 7692 11388 7744
rect 15476 7760 15528 7812
rect 16488 7760 16540 7812
rect 16580 7692 16632 7744
rect 17132 7692 17184 7744
rect 18972 7760 19024 7812
rect 19432 7760 19484 7812
rect 18328 7692 18380 7744
rect 22192 7760 22244 7812
rect 26148 7760 26200 7812
rect 26240 7760 26292 7812
rect 26516 7803 26568 7812
rect 26516 7769 26525 7803
rect 26525 7769 26559 7803
rect 26559 7769 26568 7803
rect 26516 7760 26568 7769
rect 21272 7692 21324 7744
rect 21824 7692 21876 7744
rect 22560 7692 22612 7744
rect 31668 7896 31720 7948
rect 35716 7896 35768 7948
rect 36084 7896 36136 7948
rect 27896 7828 27948 7880
rect 28264 7803 28316 7812
rect 28264 7769 28273 7803
rect 28273 7769 28307 7803
rect 28307 7769 28316 7803
rect 28264 7760 28316 7769
rect 28540 7828 28592 7880
rect 29368 7828 29420 7880
rect 33232 7828 33284 7880
rect 33508 7871 33560 7880
rect 33508 7837 33517 7871
rect 33517 7837 33551 7871
rect 33551 7837 33560 7871
rect 33508 7828 33560 7837
rect 34244 7828 34296 7880
rect 36820 7871 36872 7880
rect 27896 7692 27948 7744
rect 30012 7692 30064 7744
rect 33600 7803 33652 7812
rect 31576 7692 31628 7744
rect 31668 7692 31720 7744
rect 33600 7769 33609 7803
rect 33609 7769 33643 7803
rect 33643 7769 33652 7803
rect 33600 7760 33652 7769
rect 36820 7837 36829 7871
rect 36829 7837 36863 7871
rect 36863 7837 36872 7871
rect 36820 7828 36872 7837
rect 37924 7828 37976 7880
rect 34060 7692 34112 7744
rect 38108 7760 38160 7812
rect 35256 7692 35308 7744
rect 35716 7692 35768 7744
rect 38200 7735 38252 7744
rect 38200 7701 38209 7735
rect 38209 7701 38243 7735
rect 38243 7701 38252 7735
rect 38200 7692 38252 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3976 7531 4028 7540
rect 3976 7497 3985 7531
rect 3985 7497 4019 7531
rect 4019 7497 4028 7531
rect 3976 7488 4028 7497
rect 6092 7488 6144 7540
rect 2136 7463 2188 7472
rect 2136 7429 2145 7463
rect 2145 7429 2179 7463
rect 2179 7429 2188 7463
rect 2136 7420 2188 7429
rect 4804 7420 4856 7472
rect 7564 7420 7616 7472
rect 8392 7420 8444 7472
rect 11336 7488 11388 7540
rect 2964 7352 3016 7404
rect 3792 7352 3844 7404
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4160 7352 4212 7404
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5080 7352 5132 7404
rect 5632 7352 5684 7404
rect 4620 7284 4672 7336
rect 6368 7284 6420 7336
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 7564 7284 7616 7336
rect 9956 7420 10008 7472
rect 10416 7420 10468 7472
rect 11244 7420 11296 7472
rect 14464 7420 14516 7472
rect 14648 7420 14700 7472
rect 15752 7488 15804 7540
rect 16948 7488 17000 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 17776 7488 17828 7540
rect 18328 7420 18380 7472
rect 18696 7420 18748 7472
rect 20812 7488 20864 7540
rect 23572 7488 23624 7540
rect 27160 7488 27212 7540
rect 27344 7488 27396 7540
rect 28080 7488 28132 7540
rect 28264 7488 28316 7540
rect 11796 7352 11848 7404
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 11060 7284 11112 7336
rect 12348 7327 12400 7336
rect 12348 7293 12357 7327
rect 12357 7293 12391 7327
rect 12391 7293 12400 7327
rect 12348 7284 12400 7293
rect 14280 7352 14332 7404
rect 16028 7352 16080 7404
rect 20168 7352 20220 7404
rect 20720 7420 20772 7472
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 22560 7420 22612 7472
rect 25228 7420 25280 7472
rect 27436 7463 27488 7472
rect 27436 7429 27445 7463
rect 27445 7429 27479 7463
rect 27479 7429 27488 7463
rect 27436 7420 27488 7429
rect 28908 7420 28960 7472
rect 30472 7488 30524 7540
rect 31576 7488 31628 7540
rect 32036 7420 32088 7472
rect 32588 7420 32640 7472
rect 34060 7488 34112 7540
rect 35624 7488 35676 7540
rect 36820 7488 36872 7540
rect 37004 7488 37056 7540
rect 34704 7420 34756 7472
rect 35256 7420 35308 7472
rect 20352 7352 20404 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 26240 7352 26292 7404
rect 26976 7352 27028 7404
rect 16764 7284 16816 7336
rect 16856 7284 16908 7336
rect 18512 7284 18564 7336
rect 20996 7284 21048 7336
rect 21548 7284 21600 7336
rect 24032 7284 24084 7336
rect 24216 7327 24268 7336
rect 24216 7293 24225 7327
rect 24225 7293 24259 7327
rect 24259 7293 24268 7327
rect 24216 7284 24268 7293
rect 26700 7284 26752 7336
rect 27528 7284 27580 7336
rect 29092 7352 29144 7404
rect 29368 7395 29420 7404
rect 29368 7361 29377 7395
rect 29377 7361 29411 7395
rect 29411 7361 29420 7395
rect 29368 7352 29420 7361
rect 31852 7352 31904 7404
rect 33140 7352 33192 7404
rect 33508 7395 33560 7404
rect 33508 7361 33517 7395
rect 33517 7361 33551 7395
rect 33551 7361 33560 7395
rect 33508 7352 33560 7361
rect 28908 7284 28960 7336
rect 5448 7216 5500 7268
rect 9036 7216 9088 7268
rect 12256 7216 12308 7268
rect 13728 7216 13780 7268
rect 16396 7216 16448 7268
rect 2688 7148 2740 7200
rect 3516 7148 3568 7200
rect 6552 7148 6604 7200
rect 11796 7148 11848 7200
rect 14740 7148 14792 7200
rect 16212 7148 16264 7200
rect 16948 7148 17000 7200
rect 17132 7148 17184 7200
rect 17500 7148 17552 7200
rect 19432 7216 19484 7268
rect 20628 7216 20680 7268
rect 26608 7216 26660 7268
rect 33692 7284 33744 7336
rect 35716 7284 35768 7336
rect 37004 7352 37056 7404
rect 37924 7352 37976 7404
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 32864 7216 32916 7268
rect 20168 7148 20220 7200
rect 20812 7148 20864 7200
rect 25872 7148 25924 7200
rect 28540 7148 28592 7200
rect 28816 7148 28868 7200
rect 31300 7148 31352 7200
rect 32036 7148 32088 7200
rect 32220 7148 32272 7200
rect 33324 7148 33376 7200
rect 34152 7148 34204 7200
rect 35624 7148 35676 7200
rect 36636 7148 36688 7200
rect 38108 7191 38160 7200
rect 38108 7157 38117 7191
rect 38117 7157 38151 7191
rect 38151 7157 38160 7191
rect 38108 7148 38160 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3608 6944 3660 6996
rect 4160 6944 4212 6996
rect 5080 6944 5132 6996
rect 11888 6944 11940 6996
rect 12072 6944 12124 6996
rect 2964 6876 3016 6928
rect 12440 6944 12492 6996
rect 13728 6944 13780 6996
rect 14464 6944 14516 6996
rect 16948 6944 17000 6996
rect 20352 6944 20404 6996
rect 21548 6944 21600 6996
rect 21640 6944 21692 6996
rect 4804 6808 4856 6860
rect 15384 6876 15436 6928
rect 16120 6876 16172 6928
rect 17500 6876 17552 6928
rect 20628 6876 20680 6928
rect 22284 6944 22336 6996
rect 22836 6944 22888 6996
rect 24032 6944 24084 6996
rect 26332 6944 26384 6996
rect 28264 6944 28316 6996
rect 29828 6944 29880 6996
rect 30012 6987 30064 6996
rect 30012 6953 30042 6987
rect 30042 6953 30064 6987
rect 30012 6944 30064 6953
rect 7564 6808 7616 6860
rect 9312 6808 9364 6860
rect 9404 6808 9456 6860
rect 11704 6808 11756 6860
rect 12348 6808 12400 6860
rect 16856 6808 16908 6860
rect 17040 6808 17092 6860
rect 2136 6740 2188 6792
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 3976 6740 4028 6792
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 5356 6604 5408 6656
rect 5540 6604 5592 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7840 6672 7892 6724
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 9864 6672 9916 6724
rect 10968 6740 11020 6792
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 13360 6740 13412 6792
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 10600 6715 10652 6724
rect 10600 6681 10609 6715
rect 10609 6681 10643 6715
rect 10643 6681 10652 6715
rect 10600 6672 10652 6681
rect 10692 6672 10744 6724
rect 11980 6672 12032 6724
rect 14280 6715 14332 6724
rect 14280 6681 14289 6715
rect 14289 6681 14323 6715
rect 14323 6681 14332 6715
rect 14280 6672 14332 6681
rect 8392 6604 8444 6656
rect 8484 6604 8536 6656
rect 11612 6604 11664 6656
rect 12072 6604 12124 6656
rect 14096 6604 14148 6656
rect 14188 6604 14240 6656
rect 15108 6672 15160 6724
rect 18788 6740 18840 6792
rect 16764 6672 16816 6724
rect 17960 6672 18012 6724
rect 19156 6740 19208 6792
rect 20720 6783 20772 6792
rect 20720 6749 20729 6783
rect 20729 6749 20763 6783
rect 20763 6749 20772 6783
rect 20720 6740 20772 6749
rect 22744 6783 22796 6792
rect 22744 6749 22753 6783
rect 22753 6749 22787 6783
rect 22787 6749 22796 6783
rect 22744 6740 22796 6749
rect 22836 6740 22888 6792
rect 26148 6808 26200 6860
rect 26976 6808 27028 6860
rect 27160 6808 27212 6860
rect 27712 6808 27764 6860
rect 29368 6808 29420 6860
rect 33692 6944 33744 6996
rect 34060 6944 34112 6996
rect 36268 6944 36320 6996
rect 34428 6876 34480 6928
rect 32404 6851 32456 6860
rect 32404 6817 32413 6851
rect 32413 6817 32447 6851
rect 32447 6817 32456 6851
rect 32404 6808 32456 6817
rect 36084 6876 36136 6928
rect 25228 6783 25280 6792
rect 20444 6672 20496 6724
rect 23664 6672 23716 6724
rect 25228 6749 25237 6783
rect 25237 6749 25271 6783
rect 25271 6749 25280 6783
rect 25228 6740 25280 6749
rect 27804 6740 27856 6792
rect 31668 6740 31720 6792
rect 32956 6740 33008 6792
rect 33784 6740 33836 6792
rect 34704 6808 34756 6860
rect 34336 6740 34388 6792
rect 35716 6808 35768 6860
rect 35624 6740 35676 6792
rect 36176 6783 36228 6792
rect 36176 6749 36185 6783
rect 36185 6749 36219 6783
rect 36219 6749 36228 6783
rect 36176 6740 36228 6749
rect 36728 6740 36780 6792
rect 37464 6740 37516 6792
rect 18512 6604 18564 6656
rect 19340 6604 19392 6656
rect 20996 6604 21048 6656
rect 21364 6604 21416 6656
rect 22376 6604 22428 6656
rect 23480 6604 23532 6656
rect 24308 6604 24360 6656
rect 25136 6604 25188 6656
rect 26516 6604 26568 6656
rect 30288 6672 30340 6724
rect 31576 6604 31628 6656
rect 32864 6672 32916 6724
rect 36636 6672 36688 6724
rect 33784 6604 33836 6656
rect 34060 6604 34112 6656
rect 34244 6647 34296 6656
rect 34244 6613 34253 6647
rect 34253 6613 34287 6647
rect 34287 6613 34296 6647
rect 34244 6604 34296 6613
rect 34704 6604 34756 6656
rect 35440 6604 35492 6656
rect 35624 6647 35676 6656
rect 35624 6613 35633 6647
rect 35633 6613 35667 6647
rect 35667 6613 35676 6647
rect 35624 6604 35676 6613
rect 35716 6604 35768 6656
rect 36452 6604 36504 6656
rect 38292 6604 38344 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 6460 6400 6512 6452
rect 3056 6332 3108 6384
rect 3332 6332 3384 6384
rect 5908 6332 5960 6384
rect 1492 6264 1544 6316
rect 2596 6264 2648 6316
rect 3148 6264 3200 6316
rect 4068 6264 4120 6316
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6828 6264 6880 6316
rect 9404 6400 9456 6452
rect 9496 6400 9548 6452
rect 11152 6443 11204 6452
rect 7748 6332 7800 6384
rect 8760 6332 8812 6384
rect 9956 6332 10008 6384
rect 10324 6332 10376 6384
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 11428 6332 11480 6384
rect 10968 6264 11020 6316
rect 12072 6332 12124 6384
rect 13820 6400 13872 6452
rect 14280 6400 14332 6452
rect 14832 6332 14884 6384
rect 19800 6400 19852 6452
rect 20444 6400 20496 6452
rect 22284 6400 22336 6452
rect 11704 6264 11756 6316
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 15016 6264 15068 6316
rect 16488 6332 16540 6384
rect 16580 6332 16632 6384
rect 4804 6196 4856 6248
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 5448 6128 5500 6180
rect 6736 6196 6788 6248
rect 6828 6128 6880 6180
rect 3608 6060 3660 6112
rect 4436 6060 4488 6112
rect 4988 6060 5040 6112
rect 5356 6060 5408 6112
rect 9128 6060 9180 6112
rect 10692 6128 10744 6180
rect 14096 6196 14148 6248
rect 16304 6196 16356 6248
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 17132 6196 17184 6248
rect 17592 6196 17644 6248
rect 18880 6332 18932 6384
rect 20076 6332 20128 6384
rect 22928 6400 22980 6452
rect 23020 6400 23072 6452
rect 25228 6400 25280 6452
rect 26608 6400 26660 6452
rect 28264 6400 28316 6452
rect 28908 6443 28960 6452
rect 28908 6409 28917 6443
rect 28917 6409 28951 6443
rect 28951 6409 28960 6443
rect 28908 6400 28960 6409
rect 29184 6400 29236 6452
rect 29828 6400 29880 6452
rect 20352 6264 20404 6316
rect 24492 6332 24544 6384
rect 25596 6264 25648 6316
rect 26148 6264 26200 6316
rect 18788 6239 18840 6248
rect 11336 6060 11388 6112
rect 14832 6103 14884 6112
rect 14832 6069 14841 6103
rect 14841 6069 14875 6103
rect 14875 6069 14884 6103
rect 14832 6060 14884 6069
rect 15108 6060 15160 6112
rect 17960 6060 18012 6112
rect 18788 6205 18797 6239
rect 18797 6205 18831 6239
rect 18831 6205 18840 6239
rect 18788 6196 18840 6205
rect 18880 6196 18932 6248
rect 20536 6239 20588 6248
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 20628 6196 20680 6248
rect 22008 6239 22060 6248
rect 21732 6128 21784 6180
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22376 6196 22428 6248
rect 23664 6196 23716 6248
rect 24216 6239 24268 6248
rect 24216 6205 24225 6239
rect 24225 6205 24259 6239
rect 24259 6205 24268 6239
rect 24216 6196 24268 6205
rect 25136 6196 25188 6248
rect 27436 6332 27488 6384
rect 36544 6400 36596 6452
rect 32036 6332 32088 6384
rect 32312 6375 32364 6384
rect 32312 6341 32321 6375
rect 32321 6341 32355 6375
rect 32355 6341 32364 6375
rect 32312 6332 32364 6341
rect 34428 6332 34480 6384
rect 27160 6307 27212 6316
rect 27160 6273 27169 6307
rect 27169 6273 27203 6307
rect 27203 6273 27212 6307
rect 27160 6264 27212 6273
rect 29368 6307 29420 6316
rect 29368 6273 29377 6307
rect 29377 6273 29411 6307
rect 29411 6273 29420 6307
rect 29368 6264 29420 6273
rect 31944 6264 31996 6316
rect 33508 6307 33560 6316
rect 33508 6273 33517 6307
rect 33517 6273 33551 6307
rect 33551 6273 33560 6307
rect 33508 6264 33560 6273
rect 33784 6264 33836 6316
rect 36084 6307 36136 6316
rect 36084 6273 36093 6307
rect 36093 6273 36127 6307
rect 36127 6273 36136 6307
rect 36084 6264 36136 6273
rect 20720 6060 20772 6112
rect 22100 6060 22152 6112
rect 22284 6060 22336 6112
rect 26148 6128 26200 6180
rect 27528 6196 27580 6248
rect 29184 6196 29236 6248
rect 31300 6196 31352 6248
rect 32220 6239 32272 6248
rect 32220 6205 32229 6239
rect 32229 6205 32263 6239
rect 32263 6205 32272 6239
rect 32220 6196 32272 6205
rect 32496 6239 32548 6248
rect 32496 6205 32505 6239
rect 32505 6205 32539 6239
rect 32539 6205 32548 6239
rect 32496 6196 32548 6205
rect 34152 6196 34204 6248
rect 35440 6239 35492 6248
rect 30656 6128 30708 6180
rect 35440 6205 35449 6239
rect 35449 6205 35483 6239
rect 35483 6205 35492 6239
rect 35440 6196 35492 6205
rect 35716 6196 35768 6248
rect 23480 6060 23532 6112
rect 30104 6060 30156 6112
rect 31576 6103 31628 6112
rect 31576 6069 31585 6103
rect 31585 6069 31619 6103
rect 31619 6069 31628 6103
rect 31576 6060 31628 6069
rect 31760 6060 31812 6112
rect 35624 6060 35676 6112
rect 38200 6103 38252 6112
rect 38200 6069 38209 6103
rect 38209 6069 38243 6103
rect 38243 6069 38252 6103
rect 38200 6060 38252 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2596 5856 2648 5908
rect 4252 5856 4304 5908
rect 4436 5856 4488 5908
rect 7840 5856 7892 5908
rect 1860 5831 1912 5840
rect 1860 5797 1869 5831
rect 1869 5797 1903 5831
rect 1903 5797 1912 5831
rect 1860 5788 1912 5797
rect 3884 5788 3936 5840
rect 4804 5788 4856 5840
rect 5816 5788 5868 5840
rect 6552 5788 6604 5840
rect 2688 5720 2740 5772
rect 8668 5788 8720 5840
rect 11428 5788 11480 5840
rect 11612 5788 11664 5840
rect 16396 5831 16448 5840
rect 8300 5720 8352 5772
rect 9404 5720 9456 5772
rect 9772 5763 9824 5772
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 11704 5763 11756 5772
rect 9772 5720 9824 5729
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 16396 5797 16405 5831
rect 16405 5797 16439 5831
rect 16439 5797 16448 5831
rect 16396 5788 16448 5797
rect 16304 5720 16356 5772
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 17132 5720 17184 5772
rect 17224 5720 17276 5772
rect 18788 5720 18840 5772
rect 1308 5652 1360 5704
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 6736 5652 6788 5704
rect 8208 5652 8260 5704
rect 1676 5627 1728 5636
rect 1676 5593 1685 5627
rect 1685 5593 1719 5627
rect 1719 5593 1728 5627
rect 1676 5584 1728 5593
rect 4160 5584 4212 5636
rect 5356 5627 5408 5636
rect 5356 5593 5365 5627
rect 5365 5593 5399 5627
rect 5399 5593 5408 5627
rect 5356 5584 5408 5593
rect 5448 5627 5500 5636
rect 5448 5593 5457 5627
rect 5457 5593 5491 5627
rect 5491 5593 5500 5627
rect 6368 5627 6420 5636
rect 5448 5584 5500 5593
rect 6368 5593 6377 5627
rect 6377 5593 6411 5627
rect 6411 5593 6420 5627
rect 6368 5584 6420 5593
rect 6552 5584 6604 5636
rect 7380 5584 7432 5636
rect 16580 5652 16632 5704
rect 20536 5856 20588 5908
rect 22652 5856 22704 5908
rect 22836 5856 22888 5908
rect 21732 5788 21784 5840
rect 20720 5720 20772 5772
rect 22008 5720 22060 5772
rect 24216 5720 24268 5772
rect 32312 5856 32364 5908
rect 27160 5720 27212 5772
rect 27436 5720 27488 5772
rect 1492 5516 1544 5568
rect 7748 5516 7800 5568
rect 7840 5516 7892 5568
rect 9680 5516 9732 5568
rect 10232 5584 10284 5636
rect 12716 5584 12768 5636
rect 14096 5584 14148 5636
rect 15016 5584 15068 5636
rect 17224 5584 17276 5636
rect 17408 5584 17460 5636
rect 18144 5584 18196 5636
rect 18880 5627 18932 5636
rect 18880 5593 18889 5627
rect 18889 5593 18923 5627
rect 18923 5593 18932 5627
rect 18880 5584 18932 5593
rect 11060 5516 11112 5568
rect 14740 5516 14792 5568
rect 20352 5652 20404 5704
rect 22836 5652 22888 5704
rect 20444 5584 20496 5636
rect 20996 5584 21048 5636
rect 22192 5584 22244 5636
rect 19984 5516 20036 5568
rect 24768 5652 24820 5704
rect 27712 5652 27764 5704
rect 29368 5720 29420 5772
rect 31760 5788 31812 5840
rect 33048 5788 33100 5840
rect 33140 5788 33192 5840
rect 33784 5788 33836 5840
rect 34704 5788 34756 5840
rect 35072 5788 35124 5840
rect 35440 5720 35492 5772
rect 29644 5652 29696 5704
rect 31116 5652 31168 5704
rect 34520 5652 34572 5704
rect 26332 5584 26384 5636
rect 26700 5584 26752 5636
rect 28080 5584 28132 5636
rect 28264 5584 28316 5636
rect 30288 5584 30340 5636
rect 23940 5516 23992 5568
rect 26148 5516 26200 5568
rect 26516 5516 26568 5568
rect 31392 5516 31444 5568
rect 31576 5516 31628 5568
rect 32496 5516 32548 5568
rect 35348 5584 35400 5636
rect 35624 5652 35676 5704
rect 37280 5695 37332 5704
rect 37280 5661 37289 5695
rect 37289 5661 37323 5695
rect 37323 5661 37332 5695
rect 37280 5652 37332 5661
rect 37372 5652 37424 5704
rect 34704 5516 34756 5568
rect 35532 5516 35584 5568
rect 37464 5559 37516 5568
rect 37464 5525 37473 5559
rect 37473 5525 37507 5559
rect 37507 5525 37516 5559
rect 37464 5516 37516 5525
rect 38016 5516 38068 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3332 5312 3384 5364
rect 3516 5287 3568 5296
rect 3516 5253 3525 5287
rect 3525 5253 3559 5287
rect 3559 5253 3568 5287
rect 3516 5244 3568 5253
rect 6828 5312 6880 5364
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7380 5312 7432 5364
rect 8300 5312 8352 5364
rect 8392 5312 8444 5364
rect 5172 5244 5224 5296
rect 5632 5244 5684 5296
rect 1124 5176 1176 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 9036 5244 9088 5296
rect 9128 5244 9180 5296
rect 18880 5312 18932 5364
rect 21088 5312 21140 5364
rect 26148 5312 26200 5364
rect 29184 5312 29236 5364
rect 30748 5312 30800 5364
rect 31576 5312 31628 5364
rect 32128 5312 32180 5364
rect 12624 5244 12676 5296
rect 13268 5244 13320 5296
rect 14556 5244 14608 5296
rect 15108 5244 15160 5296
rect 16120 5244 16172 5296
rect 18052 5244 18104 5296
rect 19064 5244 19116 5296
rect 24492 5244 24544 5296
rect 26056 5244 26108 5296
rect 26424 5244 26476 5296
rect 28172 5244 28224 5296
rect 6184 5176 6236 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 4620 5108 4672 5160
rect 5356 5108 5408 5160
rect 7012 5108 7064 5160
rect 7196 5108 7248 5160
rect 8300 5108 8352 5160
rect 9220 5108 9272 5160
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 13636 5108 13688 5160
rect 13820 5108 13872 5160
rect 14280 5108 14332 5160
rect 16764 5151 16816 5160
rect 5632 5040 5684 5092
rect 7840 5040 7892 5092
rect 11520 5040 11572 5092
rect 14096 5040 14148 5092
rect 16304 5083 16356 5092
rect 16304 5049 16313 5083
rect 16313 5049 16347 5083
rect 16347 5049 16356 5083
rect 16304 5040 16356 5049
rect 1308 4972 1360 5024
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 3976 4972 4028 5024
rect 9864 4972 9916 5024
rect 11060 4972 11112 5024
rect 16212 4972 16264 5024
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 17132 5108 17184 5160
rect 21272 5176 21324 5228
rect 23388 5176 23440 5228
rect 20996 5108 21048 5160
rect 22008 5151 22060 5160
rect 22008 5117 22017 5151
rect 22017 5117 22051 5151
rect 22051 5117 22060 5151
rect 22008 5108 22060 5117
rect 24308 5151 24360 5160
rect 23940 5040 23992 5092
rect 19432 4972 19484 5024
rect 21180 4972 21232 5024
rect 22744 4972 22796 5024
rect 24308 5117 24317 5151
rect 24317 5117 24351 5151
rect 24351 5117 24360 5151
rect 24308 5108 24360 5117
rect 25228 5108 25280 5160
rect 27160 5151 27212 5160
rect 27160 5117 27169 5151
rect 27169 5117 27203 5151
rect 27203 5117 27212 5151
rect 27160 5108 27212 5117
rect 30196 5244 30248 5296
rect 31852 5244 31904 5296
rect 31944 5244 31996 5296
rect 33048 5312 33100 5364
rect 35072 5244 35124 5296
rect 29184 5219 29236 5228
rect 29184 5185 29193 5219
rect 29193 5185 29227 5219
rect 29227 5185 29236 5219
rect 29184 5176 29236 5185
rect 29644 5151 29696 5160
rect 26516 5040 26568 5092
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 29644 5108 29696 5117
rect 31392 5108 31444 5160
rect 30932 5040 30984 5092
rect 25780 4972 25832 5024
rect 26700 4972 26752 5024
rect 31760 4972 31812 5024
rect 32220 5151 32272 5160
rect 32220 5117 32229 5151
rect 32229 5117 32263 5151
rect 32263 5117 32272 5151
rect 32496 5151 32548 5160
rect 32220 5108 32272 5117
rect 32496 5117 32505 5151
rect 32505 5117 32539 5151
rect 32539 5117 32548 5151
rect 32496 5108 32548 5117
rect 32588 5108 32640 5160
rect 34888 5151 34940 5160
rect 34888 5117 34897 5151
rect 34897 5117 34931 5151
rect 34931 5117 34940 5151
rect 38108 5176 38160 5228
rect 34888 5108 34940 5117
rect 38568 5108 38620 5160
rect 32312 5040 32364 5092
rect 35624 4972 35676 5024
rect 36820 5015 36872 5024
rect 36820 4981 36829 5015
rect 36829 4981 36863 5015
rect 36863 4981 36872 5015
rect 36820 4972 36872 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 848 4768 900 4820
rect 2228 4768 2280 4820
rect 8208 4768 8260 4820
rect 9772 4768 9824 4820
rect 9864 4768 9916 4820
rect 6644 4700 6696 4752
rect 16212 4768 16264 4820
rect 16580 4700 16632 4752
rect 7748 4632 7800 4684
rect 1952 4564 2004 4616
rect 3056 4607 3108 4616
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 1860 4496 1912 4548
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 4528 4564 4580 4616
rect 6736 4564 6788 4616
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 4804 4496 4856 4548
rect 7564 4496 7616 4548
rect 8944 4632 8996 4684
rect 9680 4632 9732 4684
rect 11060 4564 11112 4616
rect 13820 4632 13872 4684
rect 17224 4768 17276 4820
rect 17316 4768 17368 4820
rect 21180 4768 21232 4820
rect 21272 4768 21324 4820
rect 22192 4768 22244 4820
rect 25964 4768 26016 4820
rect 17132 4632 17184 4684
rect 17224 4632 17276 4684
rect 14096 4564 14148 4616
rect 14280 4564 14332 4616
rect 18328 4632 18380 4684
rect 18880 4632 18932 4684
rect 18696 4564 18748 4616
rect 19248 4564 19300 4616
rect 19984 4564 20036 4616
rect 9220 4539 9272 4548
rect 8668 4428 8720 4480
rect 9220 4505 9229 4539
rect 9229 4505 9263 4539
rect 9263 4505 9272 4539
rect 9220 4496 9272 4505
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 12808 4496 12860 4548
rect 11612 4428 11664 4480
rect 13544 4428 13596 4480
rect 15108 4496 15160 4548
rect 15844 4496 15896 4548
rect 17040 4496 17092 4548
rect 17408 4496 17460 4548
rect 20168 4539 20220 4548
rect 16580 4428 16632 4480
rect 20168 4505 20177 4539
rect 20177 4505 20211 4539
rect 20211 4505 20220 4539
rect 20168 4496 20220 4505
rect 24584 4700 24636 4752
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 23756 4632 23808 4684
rect 24308 4632 24360 4684
rect 25412 4632 25464 4684
rect 23204 4564 23256 4616
rect 24768 4564 24820 4616
rect 27620 4632 27672 4684
rect 33784 4768 33836 4820
rect 21272 4496 21324 4548
rect 24492 4496 24544 4548
rect 21456 4428 21508 4480
rect 21548 4428 21600 4480
rect 24216 4428 24268 4480
rect 25688 4428 25740 4480
rect 25780 4428 25832 4480
rect 26516 4496 26568 4548
rect 28080 4496 28132 4548
rect 29644 4632 29696 4684
rect 32312 4632 32364 4684
rect 32864 4632 32916 4684
rect 33692 4564 33744 4616
rect 34336 4632 34388 4684
rect 39304 4632 39356 4684
rect 34244 4607 34296 4616
rect 34244 4573 34253 4607
rect 34253 4573 34287 4607
rect 34287 4573 34296 4607
rect 34244 4564 34296 4573
rect 36728 4607 36780 4616
rect 27160 4428 27212 4480
rect 31024 4496 31076 4548
rect 31852 4496 31904 4548
rect 32496 4496 32548 4548
rect 32588 4428 32640 4480
rect 33600 4428 33652 4480
rect 33876 4496 33928 4548
rect 36728 4573 36737 4607
rect 36737 4573 36771 4607
rect 36771 4573 36780 4607
rect 36728 4564 36780 4573
rect 38844 4564 38896 4616
rect 38660 4496 38712 4548
rect 35808 4428 35860 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3700 4224 3752 4276
rect 2780 4156 2832 4208
rect 4528 4199 4580 4208
rect 4528 4165 4537 4199
rect 4537 4165 4571 4199
rect 4571 4165 4580 4199
rect 4528 4156 4580 4165
rect 4804 4224 4856 4276
rect 8576 4224 8628 4276
rect 1400 4088 1452 4140
rect 6000 4088 6052 4140
rect 7104 4156 7156 4208
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 14188 4224 14240 4276
rect 16304 4224 16356 4276
rect 13452 4156 13504 4208
rect 14924 4156 14976 4208
rect 15108 4199 15160 4208
rect 15108 4165 15117 4199
rect 15117 4165 15151 4199
rect 15151 4165 15160 4199
rect 15108 4156 15160 4165
rect 18604 4156 18656 4208
rect 18788 4156 18840 4208
rect 20996 4224 21048 4276
rect 24216 4224 24268 4276
rect 24308 4224 24360 4276
rect 24492 4224 24544 4276
rect 30288 4224 30340 4276
rect 30564 4224 30616 4276
rect 31576 4224 31628 4276
rect 31852 4224 31904 4276
rect 32588 4224 32640 4276
rect 32680 4224 32732 4276
rect 21824 4156 21876 4208
rect 22192 4199 22244 4208
rect 22192 4165 22201 4199
rect 22201 4165 22235 4199
rect 22235 4165 22244 4199
rect 22192 4156 22244 4165
rect 17960 4088 18012 4140
rect 20812 4131 20864 4140
rect 20812 4097 20821 4131
rect 20821 4097 20855 4131
rect 20855 4097 20864 4131
rect 20812 4088 20864 4097
rect 25136 4156 25188 4208
rect 25688 4156 25740 4208
rect 27528 4156 27580 4208
rect 31208 4156 31260 4208
rect 2964 4020 3016 4072
rect 3976 4020 4028 4072
rect 4160 4020 4212 4072
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 10784 4063 10836 4072
rect 664 3952 716 4004
rect 3240 3952 3292 4004
rect 6000 3995 6052 4004
rect 6000 3961 6009 3995
rect 6009 3961 6043 3995
rect 6043 3961 6052 3995
rect 6000 3952 6052 3961
rect 8208 3952 8260 4004
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11060 4020 11112 4072
rect 13360 4063 13412 4072
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 1768 3884 1820 3893
rect 2780 3884 2832 3936
rect 7564 3884 7616 3936
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 8760 3884 8812 3936
rect 12992 3884 13044 3936
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 16304 4063 16356 4072
rect 16304 4029 16313 4063
rect 16313 4029 16347 4063
rect 16347 4029 16356 4063
rect 16304 4020 16356 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18328 4063 18380 4072
rect 18328 4029 18337 4063
rect 18337 4029 18371 4063
rect 18371 4029 18380 4063
rect 18328 4020 18380 4029
rect 18420 4020 18472 4072
rect 21824 4020 21876 4072
rect 22376 4020 22428 4072
rect 23480 4020 23532 4072
rect 14096 3884 14148 3936
rect 17500 3927 17552 3936
rect 17500 3893 17509 3927
rect 17509 3893 17543 3927
rect 17543 3893 17552 3927
rect 17500 3884 17552 3893
rect 17684 3884 17736 3936
rect 20904 3952 20956 4004
rect 24216 4020 24268 4072
rect 24860 4020 24912 4072
rect 28540 4088 28592 4140
rect 29644 4131 29696 4140
rect 29644 4097 29653 4131
rect 29653 4097 29687 4131
rect 29687 4097 29696 4131
rect 29644 4088 29696 4097
rect 32312 4156 32364 4208
rect 33416 4156 33468 4208
rect 34152 4131 34204 4140
rect 34152 4097 34161 4131
rect 34161 4097 34195 4131
rect 34195 4097 34204 4131
rect 34152 4088 34204 4097
rect 35900 4088 35952 4140
rect 35992 4088 36044 4140
rect 37096 4088 37148 4140
rect 37556 4088 37608 4140
rect 25596 4020 25648 4072
rect 27160 4063 27212 4072
rect 27160 4029 27169 4063
rect 27169 4029 27203 4063
rect 27203 4029 27212 4063
rect 27160 4020 27212 4029
rect 25504 3952 25556 4004
rect 26240 3952 26292 4004
rect 20260 3884 20312 3936
rect 23020 3884 23072 3936
rect 23112 3884 23164 3936
rect 27252 3884 27304 3936
rect 27620 3884 27672 3936
rect 29184 4063 29236 4072
rect 29184 4029 29193 4063
rect 29193 4029 29227 4063
rect 29227 4029 29236 4063
rect 29184 4020 29236 4029
rect 29460 4020 29512 4072
rect 29920 4063 29972 4072
rect 29920 4029 29929 4063
rect 29929 4029 29963 4063
rect 29963 4029 29972 4063
rect 29920 4020 29972 4029
rect 30472 4020 30524 4072
rect 34428 4020 34480 4072
rect 34704 4020 34756 4072
rect 35440 4020 35492 4072
rect 35624 4063 35676 4072
rect 35624 4029 35633 4063
rect 35633 4029 35667 4063
rect 35667 4029 35676 4063
rect 35624 4020 35676 4029
rect 38660 4020 38712 4072
rect 31300 3884 31352 3936
rect 35348 3952 35400 4004
rect 33508 3884 33560 3936
rect 33784 3884 33836 3936
rect 33968 3884 34020 3936
rect 36268 3952 36320 4004
rect 36084 3884 36136 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3332 3655 3384 3664
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 2044 3408 2096 3460
rect 2596 3340 2648 3392
rect 4712 3680 4764 3732
rect 5908 3680 5960 3732
rect 7564 3680 7616 3732
rect 18788 3680 18840 3732
rect 19432 3680 19484 3732
rect 8116 3612 8168 3664
rect 10876 3612 10928 3664
rect 16580 3612 16632 3664
rect 4252 3544 4304 3596
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 7196 3544 7248 3596
rect 8760 3544 8812 3596
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 10048 3587 10100 3596
rect 10048 3553 10057 3587
rect 10057 3553 10091 3587
rect 10091 3553 10100 3587
rect 10048 3544 10100 3553
rect 6736 3476 6788 3528
rect 4068 3383 4120 3392
rect 4068 3349 4077 3383
rect 4077 3349 4111 3383
rect 4111 3349 4120 3383
rect 4068 3340 4120 3349
rect 4896 3451 4948 3460
rect 4896 3417 4905 3451
rect 4905 3417 4939 3451
rect 4939 3417 4948 3451
rect 4896 3408 4948 3417
rect 6276 3408 6328 3460
rect 7564 3408 7616 3460
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9312 3451 9364 3460
rect 9312 3417 9321 3451
rect 9321 3417 9355 3451
rect 9355 3417 9364 3451
rect 9312 3408 9364 3417
rect 9588 3408 9640 3460
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 18328 3612 18380 3664
rect 18696 3612 18748 3664
rect 22468 3612 22520 3664
rect 14280 3544 14332 3553
rect 20260 3587 20312 3596
rect 20260 3553 20269 3587
rect 20269 3553 20303 3587
rect 20303 3553 20312 3587
rect 20260 3544 20312 3553
rect 21732 3544 21784 3596
rect 28080 3680 28132 3732
rect 38200 3723 38252 3732
rect 38200 3689 38209 3723
rect 38209 3689 38243 3723
rect 38243 3689 38252 3723
rect 38200 3680 38252 3689
rect 23020 3612 23072 3664
rect 24768 3612 24820 3664
rect 25596 3544 25648 3596
rect 25780 3587 25832 3596
rect 25780 3553 25789 3587
rect 25789 3553 25823 3587
rect 25823 3553 25832 3587
rect 25780 3544 25832 3553
rect 27252 3612 27304 3664
rect 30564 3612 30616 3664
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 13728 3476 13780 3528
rect 16764 3476 16816 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 27896 3476 27948 3528
rect 11336 3451 11388 3460
rect 11336 3417 11345 3451
rect 11345 3417 11379 3451
rect 11379 3417 11388 3451
rect 11336 3408 11388 3417
rect 14648 3408 14700 3460
rect 15200 3408 15252 3460
rect 16304 3451 16356 3460
rect 16304 3417 16313 3451
rect 16313 3417 16347 3451
rect 16347 3417 16356 3451
rect 16304 3408 16356 3417
rect 17224 3408 17276 3460
rect 18972 3408 19024 3460
rect 19064 3408 19116 3460
rect 20536 3408 20588 3460
rect 20720 3408 20772 3460
rect 22652 3451 22704 3460
rect 22652 3417 22661 3451
rect 22661 3417 22695 3451
rect 22695 3417 22704 3451
rect 22652 3408 22704 3417
rect 23940 3408 23992 3460
rect 14096 3340 14148 3392
rect 18788 3340 18840 3392
rect 21824 3340 21876 3392
rect 23112 3340 23164 3392
rect 23204 3340 23256 3392
rect 26148 3408 26200 3460
rect 27712 3340 27764 3392
rect 27988 3408 28040 3460
rect 30748 3587 30800 3596
rect 30748 3553 30757 3587
rect 30757 3553 30791 3587
rect 30791 3553 30800 3587
rect 30748 3544 30800 3553
rect 30932 3587 30984 3596
rect 30932 3553 30941 3587
rect 30941 3553 30975 3587
rect 30975 3553 30984 3587
rect 32588 3587 32640 3596
rect 30932 3544 30984 3553
rect 32588 3553 32597 3587
rect 32597 3553 32631 3587
rect 32631 3553 32640 3587
rect 32588 3544 32640 3553
rect 34336 3544 34388 3596
rect 35256 3587 35308 3596
rect 35256 3553 35265 3587
rect 35265 3553 35299 3587
rect 35299 3553 35308 3587
rect 35256 3544 35308 3553
rect 38476 3544 38528 3596
rect 29736 3476 29788 3528
rect 29644 3408 29696 3460
rect 37924 3476 37976 3528
rect 33140 3408 33192 3460
rect 33968 3408 34020 3460
rect 34060 3408 34112 3460
rect 30288 3340 30340 3392
rect 30748 3340 30800 3392
rect 35348 3408 35400 3460
rect 36636 3451 36688 3460
rect 36636 3417 36645 3451
rect 36645 3417 36679 3451
rect 36679 3417 36688 3451
rect 36636 3408 36688 3417
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 3240 3068 3292 3120
rect 5172 3136 5224 3188
rect 6460 3136 6512 3188
rect 9312 3136 9364 3188
rect 9404 3136 9456 3188
rect 12900 3136 12952 3188
rect 12992 3136 13044 3188
rect 16304 3136 16356 3188
rect 4804 3068 4856 3120
rect 5540 3068 5592 3120
rect 7472 3068 7524 3120
rect 7840 3068 7892 3120
rect 8852 3068 8904 3120
rect 10876 3068 10928 3120
rect 14832 3068 14884 3120
rect 4252 3043 4304 3052
rect 1032 2864 1084 2916
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 11060 3000 11112 3052
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 17776 3136 17828 3188
rect 18052 3136 18104 3188
rect 19248 3136 19300 3188
rect 17040 3068 17092 3120
rect 21824 3136 21876 3188
rect 21916 3136 21968 3188
rect 22560 3136 22612 3188
rect 20076 3068 20128 3120
rect 21272 3111 21324 3120
rect 21272 3077 21281 3111
rect 21281 3077 21315 3111
rect 21315 3077 21324 3111
rect 21272 3068 21324 3077
rect 22192 3068 22244 3120
rect 22928 3068 22980 3120
rect 24492 3111 24544 3120
rect 24492 3077 24501 3111
rect 24501 3077 24535 3111
rect 24535 3077 24544 3111
rect 24492 3068 24544 3077
rect 24952 3068 25004 3120
rect 26332 3068 26384 3120
rect 27068 3068 27120 3120
rect 28724 3068 28776 3120
rect 31300 3136 31352 3188
rect 32680 3068 32732 3120
rect 34428 3068 34480 3120
rect 34612 3111 34664 3120
rect 34612 3077 34621 3111
rect 34621 3077 34655 3111
rect 34655 3077 34664 3111
rect 34612 3068 34664 3077
rect 34796 3068 34848 3120
rect 4896 2932 4948 2984
rect 6736 2932 6788 2984
rect 9312 2975 9364 2984
rect 9312 2941 9321 2975
rect 9321 2941 9355 2975
rect 9355 2941 9364 2975
rect 9312 2932 9364 2941
rect 9588 2975 9640 2984
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 10968 2932 11020 2984
rect 940 2796 992 2848
rect 6920 2864 6972 2916
rect 6000 2796 6052 2848
rect 9404 2796 9456 2848
rect 11612 2864 11664 2916
rect 13084 2864 13136 2916
rect 16028 2864 16080 2916
rect 16764 2932 16816 2984
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 17224 2932 17276 2984
rect 21640 3000 21692 3052
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 23848 3000 23900 3052
rect 24216 3043 24268 3052
rect 24216 3009 24225 3043
rect 24225 3009 24259 3043
rect 24259 3009 24268 3043
rect 24216 3000 24268 3009
rect 26424 3043 26476 3052
rect 26424 3009 26433 3043
rect 26433 3009 26467 3043
rect 26467 3009 26476 3043
rect 26424 3000 26476 3009
rect 36360 3043 36412 3052
rect 20812 2932 20864 2984
rect 22284 2975 22336 2984
rect 11428 2796 11480 2848
rect 12256 2796 12308 2848
rect 17684 2796 17736 2848
rect 17776 2796 17828 2848
rect 18972 2864 19024 2916
rect 20720 2864 20772 2916
rect 21088 2864 21140 2916
rect 22284 2941 22293 2975
rect 22293 2941 22327 2975
rect 22327 2941 22336 2975
rect 22284 2932 22336 2941
rect 23480 2932 23532 2984
rect 25964 2975 26016 2984
rect 18236 2796 18288 2848
rect 19248 2796 19300 2848
rect 20904 2796 20956 2848
rect 24124 2864 24176 2916
rect 24032 2796 24084 2848
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 27160 2975 27212 2984
rect 27160 2941 27169 2975
rect 27169 2941 27203 2975
rect 27203 2941 27212 2975
rect 27160 2932 27212 2941
rect 27436 2932 27488 2984
rect 27988 2932 28040 2984
rect 28632 2932 28684 2984
rect 29644 2975 29696 2984
rect 29644 2941 29653 2975
rect 29653 2941 29687 2975
rect 29687 2941 29696 2975
rect 29644 2932 29696 2941
rect 29920 2975 29972 2984
rect 29920 2941 29929 2975
rect 29929 2941 29963 2975
rect 29963 2941 29972 2975
rect 29920 2932 29972 2941
rect 31484 2932 31536 2984
rect 32312 2975 32364 2984
rect 32312 2941 32321 2975
rect 32321 2941 32355 2975
rect 32355 2941 32364 2975
rect 32312 2932 32364 2941
rect 33600 2932 33652 2984
rect 26976 2796 27028 2848
rect 27160 2796 27212 2848
rect 29644 2796 29696 2848
rect 30380 2796 30432 2848
rect 31576 2796 31628 2848
rect 36360 3009 36369 3043
rect 36369 3009 36403 3043
rect 36403 3009 36412 3043
rect 36360 3000 36412 3009
rect 37740 3043 37792 3052
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 34152 2864 34204 2916
rect 34060 2839 34112 2848
rect 34060 2805 34069 2839
rect 34069 2805 34103 2839
rect 34103 2805 34112 2839
rect 34060 2796 34112 2805
rect 34796 2796 34848 2848
rect 37464 2796 37516 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4528 2592 4580 2644
rect 4988 2592 5040 2644
rect 6184 2592 6236 2644
rect 2320 2567 2372 2576
rect 2320 2533 2329 2567
rect 2329 2533 2363 2567
rect 2363 2533 2372 2567
rect 2320 2524 2372 2533
rect 9404 2592 9456 2644
rect 11704 2592 11756 2644
rect 16580 2592 16632 2644
rect 16672 2592 16724 2644
rect 5816 2456 5868 2508
rect 6368 2456 6420 2508
rect 6736 2456 6788 2508
rect 7196 2456 7248 2508
rect 7472 2456 7524 2508
rect 9312 2456 9364 2508
rect 11060 2456 11112 2508
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 15200 2456 15252 2508
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 11152 2388 11204 2440
rect 4988 2363 5040 2372
rect 4988 2329 4997 2363
rect 4997 2329 5031 2363
rect 5031 2329 5040 2363
rect 4988 2320 5040 2329
rect 5080 2363 5132 2372
rect 5080 2329 5089 2363
rect 5089 2329 5123 2363
rect 5123 2329 5132 2363
rect 5080 2320 5132 2329
rect 5356 2320 5408 2372
rect 6920 2252 6972 2304
rect 9588 2320 9640 2372
rect 12532 2320 12584 2372
rect 13728 2363 13780 2372
rect 13728 2329 13737 2363
rect 13737 2329 13771 2363
rect 13771 2329 13780 2363
rect 13728 2320 13780 2329
rect 14464 2363 14516 2372
rect 14464 2329 14473 2363
rect 14473 2329 14507 2363
rect 14507 2329 14516 2363
rect 14464 2320 14516 2329
rect 29460 2592 29512 2644
rect 34244 2592 34296 2644
rect 16856 2499 16908 2508
rect 16856 2465 16865 2499
rect 16865 2465 16899 2499
rect 16899 2465 16908 2499
rect 16856 2456 16908 2465
rect 20168 2456 20220 2508
rect 20904 2456 20956 2508
rect 23572 2456 23624 2508
rect 23848 2456 23900 2508
rect 29644 2456 29696 2508
rect 32312 2499 32364 2508
rect 32312 2465 32321 2499
rect 32321 2465 32355 2499
rect 32355 2465 32364 2499
rect 32312 2456 32364 2465
rect 35532 2456 35584 2508
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 37648 2456 37700 2508
rect 12072 2252 12124 2304
rect 17592 2320 17644 2372
rect 18880 2363 18932 2372
rect 18880 2329 18889 2363
rect 18889 2329 18923 2363
rect 18923 2329 18932 2363
rect 18880 2320 18932 2329
rect 17224 2252 17276 2304
rect 21364 2320 21416 2372
rect 22284 2320 22336 2372
rect 23296 2320 23348 2372
rect 23664 2320 23716 2372
rect 20720 2252 20772 2304
rect 23756 2295 23808 2304
rect 23756 2261 23765 2295
rect 23765 2261 23799 2295
rect 23799 2261 23808 2295
rect 23756 2252 23808 2261
rect 24124 2320 24176 2372
rect 24860 2363 24912 2372
rect 24860 2329 24869 2363
rect 24869 2329 24903 2363
rect 24903 2329 24912 2363
rect 24860 2320 24912 2329
rect 27436 2363 27488 2372
rect 27436 2329 27445 2363
rect 27445 2329 27479 2363
rect 27479 2329 27488 2363
rect 27436 2320 27488 2329
rect 29920 2320 29972 2372
rect 30012 2363 30064 2372
rect 30012 2329 30021 2363
rect 30021 2329 30055 2363
rect 30055 2329 30064 2363
rect 30012 2320 30064 2329
rect 31300 2320 31352 2372
rect 28356 2252 28408 2304
rect 34704 2320 34756 2372
rect 36452 2320 36504 2372
rect 36636 2295 36688 2304
rect 36636 2261 36645 2295
rect 36645 2261 36679 2295
rect 36679 2261 36688 2295
rect 36636 2252 36688 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 4068 2048 4120 2100
rect 22652 2048 22704 2100
rect 23756 2048 23808 2100
rect 24768 2048 24820 2100
rect 29920 2048 29972 2100
rect 32772 2048 32824 2100
rect 2688 1980 2740 2032
rect 5080 1980 5132 2032
rect 6920 1980 6972 2032
rect 10324 1980 10376 2032
rect 10692 1980 10744 2032
rect 13728 1980 13780 2032
rect 17132 1980 17184 2032
rect 17224 1980 17276 2032
rect 26700 1980 26752 2032
rect 34060 1980 34112 2032
rect 3792 1912 3844 1964
rect 11704 1912 11756 1964
rect 14464 1912 14516 1964
rect 16580 1912 16632 1964
rect 16672 1912 16724 1964
rect 14096 1844 14148 1896
rect 17592 1844 17644 1896
rect 21364 1912 21416 1964
rect 22284 1844 22336 1896
rect 9588 1776 9640 1828
rect 18236 1776 18288 1828
rect 27620 1912 27672 1964
rect 28448 1912 28500 1964
rect 36636 2048 36688 2100
rect 39028 1776 39080 1828
rect 3148 1708 3200 1760
rect 18512 1708 18564 1760
rect 11336 1640 11388 1692
rect 18880 1640 18932 1692
rect 16580 1572 16632 1624
rect 23756 1572 23808 1624
rect 29644 1572 29696 1624
rect 37004 1572 37056 1624
rect 20 1300 72 1352
rect 2504 1300 2556 1352
<< metal2 >>
rect 18 39200 74 39800
rect 662 39200 718 39800
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5170 39200 5226 39800
rect 5814 39200 5870 39800
rect 7102 39200 7158 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 9678 39200 9734 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14186 39200 14242 39800
rect 15474 39200 15530 39800
rect 16118 39200 16174 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 18694 39200 18750 39800
rect 19982 39200 20038 39800
rect 20626 39200 20682 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25134 39200 25190 39800
rect 25778 39200 25834 39800
rect 27066 39200 27122 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 32 37330 60 39200
rect 20 37324 72 37330
rect 20 37266 72 37272
rect 676 36378 704 39200
rect 1320 36922 1348 39200
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 2608 37210 2636 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 1308 36916 1360 36922
rect 1308 36858 1360 36864
rect 1596 36825 1624 37198
rect 2608 37182 2820 37210
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2884 36922 2912 38791
rect 3146 38176 3202 38185
rect 3146 38111 3202 38120
rect 2964 37324 3016 37330
rect 2964 37266 3016 37272
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 1582 36816 1638 36825
rect 1582 36751 1638 36760
rect 2320 36780 2372 36786
rect 2320 36722 2372 36728
rect 664 36372 716 36378
rect 664 36314 716 36320
rect 1676 36168 1728 36174
rect 1674 36136 1676 36145
rect 1728 36136 1730 36145
rect 1674 36071 1730 36080
rect 2228 36100 2280 36106
rect 2228 36042 2280 36048
rect 1860 35692 1912 35698
rect 1860 35634 1912 35640
rect 1768 35488 1820 35494
rect 1766 35456 1768 35465
rect 1820 35456 1822 35465
rect 1766 35391 1822 35400
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1780 34105 1808 34546
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 1766 33416 1822 33425
rect 1766 33351 1768 33360
rect 1820 33351 1822 33360
rect 1768 33322 1820 33328
rect 1872 32366 1900 35634
rect 2044 33448 2096 33454
rect 2044 33390 2096 33396
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1860 32360 1912 32366
rect 1860 32302 1912 32308
rect 1596 32065 1624 32302
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 846 27024 902 27033
rect 846 26959 902 26968
rect 860 4826 888 26959
rect 1688 23866 1716 31758
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 31385 1808 31622
rect 1766 31376 1822 31385
rect 1766 31311 1822 31320
rect 1768 30728 1820 30734
rect 1766 30696 1768 30705
rect 1820 30696 1822 30705
rect 1766 30631 1822 30640
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1780 29345 1808 29446
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1768 29028 1820 29034
rect 1768 28970 1820 28976
rect 1780 28665 1808 28970
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1872 28150 1900 32302
rect 1860 28144 1912 28150
rect 1860 28086 1912 28092
rect 1768 27328 1820 27334
rect 1766 27296 1768 27305
rect 1820 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1780 26625 1808 26930
rect 1766 26616 1822 26625
rect 1766 26551 1822 26560
rect 1766 25256 1822 25265
rect 1766 25191 1822 25200
rect 1780 25158 1808 25191
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1768 24812 1820 24818
rect 1768 24754 1820 24760
rect 1780 24585 1808 24754
rect 1860 24608 1912 24614
rect 1766 24576 1822 24585
rect 1860 24550 1912 24556
rect 1766 24511 1822 24520
rect 1872 24206 1900 24550
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1780 23905 1808 24142
rect 1766 23896 1822 23905
rect 1676 23860 1728 23866
rect 1766 23831 1822 23840
rect 1676 23802 1728 23808
rect 940 23044 992 23050
rect 940 22986 992 22992
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 664 4004 716 4010
rect 664 3946 716 3952
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 32 800 60 1294
rect 676 800 704 3946
rect 952 2854 980 22986
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1768 21888 1820 21894
rect 1766 21856 1768 21865
rect 1820 21856 1822 21865
rect 1766 21791 1822 21800
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 1780 20505 1808 20742
rect 1766 20496 1822 20505
rect 1872 20466 1900 24142
rect 1952 22160 2004 22166
rect 1952 22102 2004 22108
rect 1766 20431 1822 20440
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1584 19848 1636 19854
rect 1582 19816 1584 19825
rect 1636 19816 1638 19825
rect 1582 19751 1638 19760
rect 1780 19378 1808 20198
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1768 19168 1820 19174
rect 1766 19136 1768 19145
rect 1820 19136 1822 19145
rect 1766 19071 1822 19080
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 1584 17128 1636 17134
rect 1582 17096 1584 17105
rect 1636 17096 1638 17105
rect 1582 17031 1638 17040
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1124 14816 1176 14822
rect 1124 14758 1176 14764
rect 1032 11280 1084 11286
rect 1032 11222 1084 11228
rect 1044 2922 1072 11222
rect 1136 5234 1164 14758
rect 1504 12900 1532 16390
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1688 15065 1716 15370
rect 1674 15056 1730 15065
rect 1674 14991 1730 15000
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1780 14278 1808 14311
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1872 13841 1900 15370
rect 1858 13832 1914 13841
rect 1858 13767 1914 13776
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 13025 1624 13262
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1964 12918 1992 22102
rect 2056 13462 2084 33390
rect 2240 16522 2268 36042
rect 2332 35834 2360 36722
rect 2412 36712 2464 36718
rect 2412 36654 2464 36660
rect 2320 35828 2372 35834
rect 2320 35770 2372 35776
rect 2424 23866 2452 36654
rect 2976 36174 3004 37266
rect 3056 37256 3108 37262
rect 3056 37198 3108 37204
rect 3068 36922 3096 37198
rect 3160 36922 3188 38111
rect 3252 37262 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 4632 37126 4660 37726
rect 5184 37262 5212 39200
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 3056 36916 3108 36922
rect 3056 36858 3108 36864
rect 3148 36916 3200 36922
rect 3148 36858 3200 36864
rect 3988 36718 4016 37062
rect 3976 36712 4028 36718
rect 3976 36654 4028 36660
rect 5092 36650 5120 37198
rect 5828 37126 5856 39200
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 5356 37120 5408 37126
rect 5356 37062 5408 37068
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 5080 36644 5132 36650
rect 5080 36586 5132 36592
rect 5368 36582 5396 37062
rect 5448 36848 5500 36854
rect 5448 36790 5500 36796
rect 5356 36576 5408 36582
rect 5356 36518 5408 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2688 36168 2740 36174
rect 2688 36110 2740 36116
rect 2964 36168 3016 36174
rect 2964 36110 3016 36116
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 2608 29714 2636 34682
rect 2700 32570 2728 36110
rect 5460 36106 5488 36790
rect 5448 36100 5500 36106
rect 5448 36042 5500 36048
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4620 33516 4672 33522
rect 4620 33458 4672 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 2688 32564 2740 32570
rect 2688 32506 2740 32512
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30938 4660 33458
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 2596 29708 2648 29714
rect 2596 29650 2648 29656
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2608 23497 2636 23666
rect 2594 23488 2650 23497
rect 2594 23423 2650 23432
rect 4080 23322 4108 27406
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 5460 22094 5488 36042
rect 5816 36032 5868 36038
rect 5816 35974 5868 35980
rect 6460 36032 6512 36038
rect 6460 35974 6512 35980
rect 5828 33522 5856 35974
rect 5816 33516 5868 33522
rect 5816 33458 5868 33464
rect 6472 31890 6500 35974
rect 6460 31884 6512 31890
rect 6460 31826 6512 31832
rect 6092 31816 6144 31822
rect 6092 31758 6144 31764
rect 6000 25152 6052 25158
rect 6000 25094 6052 25100
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5552 23118 5580 24006
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5368 22066 5488 22094
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 2318 18592 2374 18601
rect 2318 18527 2374 18536
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2332 14618 2360 18527
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 1952 12912 2004 12918
rect 1504 12872 1624 12900
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 1320 5710 1348 9658
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 8265 1440 9522
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 1124 5228 1176 5234
rect 1124 5170 1176 5176
rect 1308 5024 1360 5030
rect 1308 4966 1360 4972
rect 1032 2916 1084 2922
rect 1032 2858 1084 2864
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 1320 800 1348 4966
rect 1412 4146 1440 8026
rect 1504 6322 1532 10134
rect 1596 8090 1624 12872
rect 1952 12854 2004 12860
rect 3988 12850 4016 13126
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 1688 12345 1716 12786
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 1768 11008 1820 11014
rect 1766 10976 1768 10985
rect 1820 10976 1822 10985
rect 1766 10911 1822 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10305 1808 10610
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1780 9625 1808 9998
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7585 1808 7686
rect 1766 7576 1822 7585
rect 1766 7511 1822 7520
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1766 6216 1822 6225
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 1858 5944 1914 5953
rect 1858 5879 1914 5888
rect 1872 5846 1900 5879
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1492 5568 1544 5574
rect 1688 5545 1716 5578
rect 1492 5510 1544 5516
rect 1674 5536 1730 5545
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1504 1465 1532 5510
rect 1674 5471 1730 5480
rect 1964 4622 1992 8298
rect 2148 7478 2176 9998
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2240 9042 2268 9454
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2240 7290 2268 8978
rect 2148 7262 2268 7290
rect 2148 6798 2176 7262
rect 2226 7168 2282 7177
rect 2226 7103 2282 7112
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1688 2825 1716 4490
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3505 1808 3878
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1674 2816 1730 2825
rect 1674 2751 1730 2760
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 18 200 74 800
rect 662 200 718 800
rect 1306 200 1362 800
rect 1872 785 1900 4490
rect 1950 3632 2006 3641
rect 1950 3567 2006 3576
rect 1964 3534 1992 3567
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 2056 3466 2084 6598
rect 2148 5545 2176 6734
rect 2134 5536 2190 5545
rect 2134 5471 2190 5480
rect 2240 4826 2268 7103
rect 2332 5234 2360 11494
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10062 2544 10406
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2226 3496 2282 3505
rect 2044 3460 2096 3466
rect 2226 3431 2282 3440
rect 2044 3402 2096 3408
rect 2240 3194 2268 3431
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2318 2680 2374 2689
rect 2318 2615 2374 2624
rect 2332 2582 2360 2615
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 2424 2446 2452 9862
rect 2608 8974 2636 10066
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2608 8498 2636 8910
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2700 7834 2728 9318
rect 2792 7936 2820 10610
rect 2976 10266 3004 10610
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 8430 2912 9998
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2792 7908 2912 7936
rect 2700 7806 2820 7834
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 5114 2544 7686
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2596 6792 2648 6798
rect 2594 6760 2596 6769
rect 2648 6760 2650 6769
rect 2594 6695 2650 6704
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2608 5914 2636 6258
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2700 5778 2728 7142
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2516 5086 2728 5114
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2516 1358 2544 4966
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 2608 800 2636 3334
rect 2700 2038 2728 5086
rect 2792 4214 2820 7806
rect 2884 4865 2912 7908
rect 2976 7410 3004 10202
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3068 8809 3096 8842
rect 3054 8800 3110 8809
rect 3054 8735 3110 8744
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2870 4856 2926 4865
rect 2870 4791 2926 4800
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2976 4078 3004 6870
rect 3068 6390 3096 7822
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3160 6322 3188 11290
rect 3252 9586 3280 11494
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3344 10538 3372 10678
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 8498 3280 9114
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3252 5710 3280 8298
rect 3344 7993 3372 9318
rect 3330 7984 3386 7993
rect 3330 7919 3386 7928
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3344 6390 3372 7686
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3054 4720 3110 4729
rect 3054 4655 3110 4664
rect 3068 4622 3096 4655
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3252 4010 3280 4422
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3602 2820 3878
rect 3344 3670 3372 5306
rect 3436 5166 3464 10406
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 7449 3556 8774
rect 3514 7440 3570 7449
rect 3514 7375 3570 7384
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 5302 3556 7142
rect 3620 7002 3648 10406
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3620 4185 3648 6054
rect 3712 4282 3740 8230
rect 3804 8022 3832 12582
rect 3896 12345 3924 12718
rect 4080 12481 4108 20742
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4986 15600 5042 15609
rect 4986 15535 5042 15544
rect 5000 15502 5028 15535
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4066 12472 4122 12481
rect 4214 12475 4522 12484
rect 4066 12407 4122 12416
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 10169 4108 11086
rect 4632 11014 4660 11630
rect 4908 11082 4936 12582
rect 5000 11218 5028 15438
rect 5092 13705 5120 17138
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5078 13696 5134 13705
rect 5078 13631 5134 13640
rect 5184 13326 5212 15846
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5092 12442 5120 12786
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 4632 9586 4660 10610
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3896 7410 3924 9386
rect 4080 9110 4108 9386
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3988 7546 4016 8842
rect 4250 8664 4306 8673
rect 4250 8599 4306 8608
rect 4264 8498 4292 8599
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7750 4108 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4632 7585 4660 9318
rect 4724 8809 4752 9522
rect 4710 8800 4766 8809
rect 4710 8735 4766 8744
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4724 8090 4752 8570
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4618 7576 4674 7585
rect 3976 7540 4028 7546
rect 4816 7562 4844 9862
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 7970 4936 9454
rect 5000 8265 5028 9998
rect 4986 8256 5042 8265
rect 4986 8191 5042 8200
rect 4908 7942 5028 7970
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4618 7511 4674 7520
rect 4724 7534 4844 7562
rect 3976 7482 4028 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2688 2032 2740 2038
rect 2688 1974 2740 1980
rect 3160 1766 3188 2382
rect 3148 1760 3200 1766
rect 3148 1702 3200 1708
rect 3252 800 3280 3062
rect 3804 1970 3832 7346
rect 4172 7188 4200 7346
rect 4540 7313 4568 7346
rect 4620 7336 4672 7342
rect 4526 7304 4582 7313
rect 4620 7278 4672 7284
rect 4526 7239 4582 7248
rect 4080 7160 4200 7188
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3882 6624 3938 6633
rect 3882 6559 3938 6568
rect 3896 5846 3924 6559
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3988 5030 4016 6734
rect 4080 6322 4108 7160
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4172 6202 4200 6938
rect 4252 6792 4304 6798
rect 4304 6752 4476 6780
rect 4252 6734 4304 6740
rect 4250 6352 4306 6361
rect 4250 6287 4252 6296
rect 4304 6287 4306 6296
rect 4252 6258 4304 6264
rect 4080 6174 4200 6202
rect 4080 5896 4108 6174
rect 4448 6118 4476 6752
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4252 5908 4304 5914
rect 4080 5868 4200 5896
rect 4172 5642 4200 5868
rect 4252 5850 4304 5856
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4264 5817 4292 5850
rect 4250 5808 4306 5817
rect 4250 5743 4306 5752
rect 4264 5710 4292 5743
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3976 5024 4028 5030
rect 4448 5012 4476 5850
rect 4632 5166 4660 7278
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4448 4984 4660 5012
rect 3976 4966 4028 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4706 4660 4984
rect 4540 4678 4660 4706
rect 4540 4622 4568 4678
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4526 4312 4582 4321
rect 4526 4247 4582 4256
rect 4540 4214 4568 4247
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 3976 4072 4028 4078
rect 3974 4040 3976 4049
rect 4160 4072 4212 4078
rect 4028 4040 4030 4049
rect 3974 3975 4030 3984
rect 4080 4020 4160 4026
rect 4080 4014 4212 4020
rect 4080 3998 4200 4014
rect 4080 3618 4108 3998
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4724 3738 4752 7534
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4816 6866 4844 7414
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5846 4844 6190
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4816 4282 4844 4490
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4080 3602 4292 3618
rect 4080 3596 4304 3602
rect 4080 3590 4252 3596
rect 4252 3538 4304 3544
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 3233 4016 3470
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3974 3224 4030 3233
rect 3974 3159 4030 3168
rect 4080 2106 4108 3334
rect 4264 3058 4292 3538
rect 4908 3466 4936 7822
rect 5000 6202 5028 7942
rect 5092 7410 5120 11018
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5078 7032 5134 7041
rect 5078 6967 5080 6976
rect 5132 6967 5134 6976
rect 5080 6938 5132 6944
rect 5078 6896 5134 6905
rect 5078 6831 5134 6840
rect 5092 6798 5120 6831
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5000 6174 5120 6202
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4816 2961 4844 3062
rect 4908 2990 4936 3402
rect 4896 2984 4948 2990
rect 4802 2952 4858 2961
rect 5000 2961 5028 6054
rect 5092 3369 5120 6174
rect 5184 5302 5212 11154
rect 5276 10554 5304 16594
rect 5368 11529 5396 22066
rect 5552 22030 5580 22374
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5460 17202 5488 19314
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5828 16522 5856 17138
rect 5816 16516 5868 16522
rect 5816 16458 5868 16464
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 15366 5488 16390
rect 5908 15428 5960 15434
rect 5908 15370 5960 15376
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5920 14482 5948 15370
rect 6012 15026 6040 25094
rect 6104 18222 6132 31758
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 6380 28762 6408 29582
rect 6368 28756 6420 28762
rect 6368 28698 6420 28704
rect 6460 23656 6512 23662
rect 6460 23598 6512 23604
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 14074 5948 14282
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 12238 5488 13874
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 5276 10526 5396 10554
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5276 5012 5304 10406
rect 5368 10062 5396 10526
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5460 9586 5488 12174
rect 5552 10674 5580 13398
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6012 12306 6040 12378
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9722 5580 9862
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 9489 5580 9522
rect 5538 9480 5594 9489
rect 5538 9415 5594 9424
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8566 5488 9318
rect 5538 9072 5594 9081
rect 5538 9007 5594 9016
rect 5552 8974 5580 9007
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5354 8120 5410 8129
rect 5354 8055 5356 8064
rect 5408 8055 5410 8064
rect 5356 8026 5408 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5356 7880 5408 7886
rect 5354 7848 5356 7857
rect 5408 7848 5410 7857
rect 5354 7783 5410 7792
rect 5460 7274 5488 7890
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5552 6746 5580 8774
rect 5644 7410 5672 10678
rect 5736 8838 5764 12106
rect 6012 11762 6040 12242
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5828 11218 5856 11630
rect 6104 11234 6132 14758
rect 6196 11665 6224 19926
rect 6472 18850 6500 23598
rect 6564 19242 6592 37198
rect 6920 36712 6972 36718
rect 6920 36654 6972 36660
rect 6932 31346 6960 36654
rect 7116 36174 7144 39200
rect 7760 37126 7788 39200
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7852 36854 7880 37198
rect 7840 36848 7892 36854
rect 7840 36790 7892 36796
rect 9048 36786 9076 39200
rect 9692 37262 9720 39200
rect 10336 37330 10364 39200
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 10508 37188 10560 37194
rect 10508 37130 10560 37136
rect 10692 37188 10744 37194
rect 10692 37130 10744 37136
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 10324 36780 10376 36786
rect 10324 36722 10376 36728
rect 9036 36576 9088 36582
rect 9036 36518 9088 36524
rect 9404 36576 9456 36582
rect 9404 36518 9456 36524
rect 7104 36168 7156 36174
rect 7104 36110 7156 36116
rect 8944 33312 8996 33318
rect 8944 33254 8996 33260
rect 6920 31340 6972 31346
rect 6920 31282 6972 31288
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6656 28218 6684 29106
rect 6748 28558 6776 30534
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 7392 26926 7420 31078
rect 8956 30802 8984 33254
rect 9048 31822 9076 36518
rect 9128 31952 9180 31958
rect 9128 31894 9180 31900
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 8944 30796 8996 30802
rect 8944 30738 8996 30744
rect 9140 29646 9168 31894
rect 9416 31822 9444 36518
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 9496 29776 9548 29782
rect 9496 29718 9548 29724
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9140 28626 9168 29582
rect 9324 29306 9352 29582
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7484 27538 7512 28358
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 7564 27396 7616 27402
rect 7564 27338 7616 27344
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20602 6868 20878
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6472 18822 6592 18850
rect 6564 18766 6592 18822
rect 6552 18760 6604 18766
rect 6550 18728 6552 18737
rect 6604 18728 6606 18737
rect 6550 18663 6606 18672
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6564 14346 6592 14554
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6182 11656 6238 11665
rect 6182 11591 6238 11600
rect 5816 11212 5868 11218
rect 6104 11206 6224 11234
rect 5816 11154 5868 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5920 10849 5948 11018
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5906 10840 5962 10849
rect 5816 10804 5868 10810
rect 5906 10775 5962 10784
rect 5816 10746 5868 10752
rect 5828 10470 5856 10746
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5816 10056 5868 10062
rect 5814 10024 5816 10033
rect 5868 10024 5870 10033
rect 5814 9959 5870 9968
rect 5908 9648 5960 9654
rect 5906 9616 5908 9625
rect 5960 9616 5962 9625
rect 5906 9551 5962 9560
rect 5908 9512 5960 9518
rect 5828 9472 5908 9500
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5828 7818 5856 9472
rect 5908 9454 5960 9460
rect 6012 9364 6040 10950
rect 5920 9336 6040 9364
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5552 6718 5672 6746
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5368 6118 5396 6598
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5460 5642 5488 6122
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5368 5166 5396 5578
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5276 4984 5488 5012
rect 5078 3360 5134 3369
rect 5078 3295 5134 3304
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4896 2926 4948 2932
rect 4986 2952 5042 2961
rect 4802 2887 4858 2896
rect 4986 2887 5042 2896
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4158 2544 4214 2553
rect 4158 2479 4214 2488
rect 4172 2446 4200 2479
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 4540 800 4568 2586
rect 5000 2378 5028 2586
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 5092 2038 5120 2314
rect 5080 2032 5132 2038
rect 5080 1974 5132 1980
rect 5184 800 5212 3130
rect 5460 2774 5488 4984
rect 5552 3126 5580 6598
rect 5644 5302 5672 6718
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5630 5128 5686 5137
rect 5630 5063 5632 5072
rect 5684 5063 5686 5072
rect 5632 5034 5684 5040
rect 5736 5001 5764 7754
rect 5828 5846 5856 7754
rect 5920 6390 5948 9336
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5722 4992 5778 5001
rect 5722 4927 5778 4936
rect 5736 3720 5764 4927
rect 6012 4146 6040 8910
rect 6104 8401 6132 11086
rect 6196 9217 6224 11206
rect 6288 10266 6316 11766
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6366 10976 6422 10985
rect 6366 10911 6422 10920
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9897 6316 9998
rect 6274 9888 6330 9897
rect 6274 9823 6330 9832
rect 6380 9738 6408 10911
rect 6472 9761 6500 11086
rect 6288 9710 6408 9738
rect 6458 9752 6514 9761
rect 6182 9208 6238 9217
rect 6182 9143 6238 9152
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6090 8392 6146 8401
rect 6090 8327 6146 8336
rect 6196 8242 6224 8978
rect 6288 8378 6316 9710
rect 6458 9687 6514 9696
rect 6366 9616 6422 9625
rect 6366 9551 6422 9560
rect 6380 9042 6408 9551
rect 6564 9330 6592 11630
rect 6656 11121 6684 20266
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6748 17882 6776 18294
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7024 17270 7052 17478
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6748 15570 6776 17070
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6748 14890 6776 15506
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6840 14074 6868 16118
rect 6932 15094 6960 16390
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7024 15638 7052 15846
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7024 14958 7052 15370
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6642 11112 6698 11121
rect 6642 11047 6698 11056
rect 6748 10033 6776 12582
rect 7024 12434 7052 13874
rect 7300 13734 7328 24890
rect 7392 16658 7420 26862
rect 7576 26586 7604 27338
rect 8312 27130 8340 28018
rect 8484 27396 8536 27402
rect 8484 27338 8536 27344
rect 8496 27305 8524 27338
rect 8482 27296 8538 27305
rect 8482 27231 8538 27240
rect 8300 27124 8352 27130
rect 8300 27066 8352 27072
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 8496 26314 8524 27231
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 9508 25294 9536 29718
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9588 28008 9640 28014
rect 9588 27950 9640 27956
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 8208 24676 8260 24682
rect 8208 24618 8260 24624
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22710 7788 22918
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7852 22506 7880 23054
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 8220 22166 8248 24618
rect 9416 24274 9444 24686
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8404 22234 8432 22510
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8864 22094 8892 23054
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 8496 22066 8892 22094
rect 8496 22030 8524 22066
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7576 19514 7604 20402
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7392 14074 7420 15370
rect 7668 14822 7696 18158
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 6932 12406 7052 12434
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6734 10024 6790 10033
rect 6644 9988 6696 9994
rect 6734 9959 6790 9968
rect 6644 9930 6696 9936
rect 6656 9500 6684 9930
rect 6840 9654 6868 11562
rect 6932 10713 6960 12406
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6918 10704 6974 10713
rect 6918 10639 6974 10648
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 9722 6960 10542
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6828 9512 6880 9518
rect 6656 9472 6828 9500
rect 6828 9454 6880 9460
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6736 9376 6788 9382
rect 6564 9302 6684 9330
rect 6736 9318 6788 9324
rect 6656 9092 6684 9302
rect 6748 9217 6776 9318
rect 6734 9208 6790 9217
rect 6734 9143 6790 9152
rect 6564 9064 6684 9092
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6472 8922 6500 8978
rect 6380 8906 6500 8922
rect 6368 8900 6500 8906
rect 6420 8894 6500 8900
rect 6368 8842 6420 8848
rect 6564 8548 6592 9064
rect 6828 8560 6880 8566
rect 6366 8528 6422 8537
rect 6564 8520 6828 8548
rect 6828 8502 6880 8508
rect 6366 8463 6368 8472
rect 6420 8463 6422 8472
rect 6368 8434 6420 8440
rect 6828 8424 6880 8430
rect 6288 8350 6684 8378
rect 6828 8366 6880 8372
rect 6368 8288 6420 8294
rect 6196 8214 6316 8242
rect 6368 8230 6420 8236
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6104 7546 6132 7754
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6196 6798 6224 8026
rect 6288 7177 6316 8214
rect 6380 7342 6408 8230
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6552 7200 6604 7206
rect 6274 7168 6330 7177
rect 6552 7142 6604 7148
rect 6274 7103 6330 7112
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6012 4010 6040 4082
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5908 3732 5960 3738
rect 5736 3692 5908 3720
rect 5908 3674 5960 3680
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5998 2952 6054 2961
rect 5998 2887 6054 2896
rect 6012 2854 6040 2887
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5368 2746 5488 2774
rect 5368 2378 5396 2746
rect 6196 2650 6224 5170
rect 6288 3466 6316 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6366 5672 6422 5681
rect 6366 5607 6368 5616
rect 6420 5607 6422 5616
rect 6368 5578 6420 5584
rect 6380 4049 6408 5578
rect 6366 4040 6422 4049
rect 6366 3975 6422 3984
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6380 2514 6408 3975
rect 6472 3194 6500 6394
rect 6564 6322 6592 7142
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6564 5642 6592 5782
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6656 4758 6684 8350
rect 6840 7818 6868 8366
rect 6932 8362 6960 9386
rect 7024 8974 7052 12310
rect 7116 10606 7144 12650
rect 7208 12238 7236 13262
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7194 11792 7250 11801
rect 7194 11727 7196 11736
rect 7248 11727 7250 11736
rect 7196 11698 7248 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 10742 7236 11494
rect 7300 11354 7328 12854
rect 7392 12714 7420 13874
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7392 11286 7420 11766
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7024 8430 7052 8910
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6932 7324 6960 8298
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 7024 7721 7052 7890
rect 7010 7712 7066 7721
rect 7010 7647 7066 7656
rect 7012 7336 7064 7342
rect 6932 7296 7012 7324
rect 6748 6254 6776 7278
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6322 6868 6734
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6826 6216 6882 6225
rect 6826 6151 6828 6160
rect 6880 6151 6882 6160
rect 6828 6122 6880 6128
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6656 4321 6684 4694
rect 6748 4622 6776 5646
rect 6828 5364 6880 5370
rect 6932 5352 6960 7296
rect 7012 7278 7064 7284
rect 7010 5536 7066 5545
rect 7010 5471 7066 5480
rect 7024 5370 7052 5471
rect 6880 5324 6960 5352
rect 7012 5364 7064 5370
rect 6828 5306 6880 5312
rect 7012 5306 7064 5312
rect 7010 5264 7066 5273
rect 7010 5199 7066 5208
rect 7024 5166 7052 5199
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6642 4312 6698 4321
rect 6642 4247 6698 4256
rect 6748 4078 6776 4558
rect 7116 4214 7144 10134
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 8276 7236 9998
rect 7300 9450 7328 10678
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7392 8537 7420 10406
rect 7484 10266 7512 14214
rect 7576 12434 7604 14282
rect 7576 12406 7696 12434
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7576 11082 7604 12038
rect 7668 11354 7696 12406
rect 7760 11762 7788 17614
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7668 10810 7696 11154
rect 7760 10985 7788 11222
rect 7852 11218 7880 14894
rect 7944 11393 7972 19994
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8312 18426 8340 18702
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8036 15201 8064 18226
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17270 8156 18158
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8220 17270 8248 17478
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8220 15570 8248 17002
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 15706 8340 16594
rect 8496 16250 8524 19450
rect 8588 19378 8616 19654
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 17746 8616 18566
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8208 15564 8260 15570
rect 8128 15524 8208 15552
rect 8022 15192 8078 15201
rect 8022 15127 8078 15136
rect 8036 13938 8064 15127
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 7930 11384 7986 11393
rect 7930 11319 7986 11328
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7746 10976 7802 10985
rect 7746 10911 7802 10920
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7470 10160 7526 10169
rect 7470 10095 7526 10104
rect 7564 10124 7616 10130
rect 7378 8528 7434 8537
rect 7378 8463 7434 8472
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7208 8248 7328 8276
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 5166 7236 7686
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3534 6776 4014
rect 7300 3618 7328 8248
rect 7392 7954 7420 8298
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 6089 7420 7754
rect 7378 6080 7434 6089
rect 7378 6015 7434 6024
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7392 5370 7420 5578
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7208 3602 7328 3618
rect 7196 3596 7328 3602
rect 7248 3590 7328 3596
rect 7196 3538 7248 3544
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6748 2990 6776 3470
rect 7484 3126 7512 10095
rect 7668 10112 7696 10746
rect 7616 10084 7696 10112
rect 7564 10066 7616 10072
rect 7576 7478 7604 10066
rect 7654 10024 7710 10033
rect 7654 9959 7656 9968
rect 7708 9959 7710 9968
rect 7656 9930 7708 9936
rect 7748 9648 7800 9654
rect 7852 9636 7880 11154
rect 8036 9738 8064 12650
rect 7800 9608 7880 9636
rect 7944 9710 8064 9738
rect 7944 9625 7972 9710
rect 8024 9648 8076 9654
rect 7930 9616 7986 9625
rect 7748 9590 7800 9596
rect 7760 8378 7788 9590
rect 8024 9590 8076 9596
rect 7930 9551 7986 9560
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 9110 7972 9454
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7668 8362 7788 8378
rect 7656 8356 7788 8362
rect 7708 8350 7788 8356
rect 7656 8298 7708 8304
rect 7746 8256 7802 8265
rect 7746 8191 7802 8200
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 6866 7604 7278
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7760 6746 7788 8191
rect 7852 8129 7880 8842
rect 7930 8392 7986 8401
rect 7930 8327 7986 8336
rect 7838 8120 7894 8129
rect 7838 8055 7894 8064
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7852 7857 7880 7890
rect 7838 7848 7894 7857
rect 7838 7783 7894 7792
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7041 7880 7686
rect 7838 7032 7894 7041
rect 7838 6967 7894 6976
rect 7838 6896 7894 6905
rect 7838 6831 7894 6840
rect 7668 6718 7788 6746
rect 7852 6730 7880 6831
rect 7840 6724 7892 6730
rect 7562 5536 7618 5545
rect 7562 5471 7618 5480
rect 7576 4554 7604 5471
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3738 7604 3878
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7562 3496 7618 3505
rect 7562 3431 7564 3440
rect 7616 3431 7618 3440
rect 7564 3402 7616 3408
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6748 2514 6776 2926
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5828 800 5856 2450
rect 6932 2394 6960 2858
rect 7194 2816 7250 2825
rect 7194 2751 7250 2760
rect 7208 2514 7236 2751
rect 7484 2514 7512 3062
rect 7668 2825 7696 6718
rect 7840 6666 7892 6672
rect 7746 6488 7802 6497
rect 7746 6423 7802 6432
rect 7760 6390 7788 6423
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7852 5574 7880 5850
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7760 4690 7788 5510
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7852 5001 7880 5034
rect 7838 4992 7894 5001
rect 7838 4927 7894 4936
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7838 3360 7894 3369
rect 7838 3295 7894 3304
rect 7852 3126 7880 3295
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7654 2816 7710 2825
rect 7944 2774 7972 8327
rect 8036 8022 8064 9590
rect 8128 9042 8156 15524
rect 8208 15506 8260 15512
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8220 14482 8248 14894
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8312 14074 8340 15030
rect 8404 14074 8432 16118
rect 8588 16046 8616 17682
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8496 14482 8524 15098
rect 8588 14550 8616 15982
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8404 12782 8432 13330
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8496 12434 8524 14418
rect 8680 14396 8708 15982
rect 8588 14368 8708 14396
rect 8588 13258 8616 14368
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8496 12406 8616 12434
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8312 10742 8340 12038
rect 8404 11830 8432 12038
rect 8496 11937 8524 12174
rect 8482 11928 8538 11937
rect 8482 11863 8538 11872
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8484 11688 8536 11694
rect 8588 11676 8616 12406
rect 8536 11648 8616 11676
rect 8484 11630 8536 11636
rect 8300 10736 8352 10742
rect 8206 10704 8262 10713
rect 8300 10678 8352 10684
rect 8206 10639 8262 10648
rect 8220 9738 8248 10639
rect 8404 10606 8432 11630
rect 8496 11014 8524 11630
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8496 10130 8524 10950
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8390 9888 8446 9897
rect 8390 9823 8446 9832
rect 8220 9710 8340 9738
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8022 7440 8078 7449
rect 8022 7375 8078 7384
rect 8036 3754 8064 7375
rect 8128 5137 8156 8570
rect 8220 8362 8248 9114
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8206 6896 8262 6905
rect 8206 6831 8262 6840
rect 8220 5710 8248 6831
rect 8312 6746 8340 9710
rect 8404 9489 8432 9823
rect 8576 9512 8628 9518
rect 8390 9480 8446 9489
rect 8446 9438 8524 9466
rect 8576 9454 8628 9460
rect 8390 9415 8446 9424
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8404 7478 8432 9143
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8496 6882 8524 9438
rect 8588 8566 8616 9454
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8588 7818 8616 8502
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8588 7721 8616 7754
rect 8574 7712 8630 7721
rect 8574 7647 8630 7656
rect 8496 6854 8616 6882
rect 8312 6718 8524 6746
rect 8496 6662 8524 6718
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8298 5808 8354 5817
rect 8298 5743 8300 5752
rect 8352 5743 8354 5752
rect 8300 5714 8352 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8404 5370 8432 6598
rect 8588 6474 8616 6854
rect 8496 6446 8616 6474
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8312 5166 8340 5306
rect 8300 5160 8352 5166
rect 8114 5128 8170 5137
rect 8300 5102 8352 5108
rect 8114 5063 8170 5072
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8220 4010 8248 4762
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8496 3942 8524 6446
rect 8680 5846 8708 13738
rect 8772 9654 8800 17614
rect 8864 13977 8892 22066
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8850 13968 8906 13977
rect 8850 13903 8906 13912
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8772 8838 8800 9386
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8864 8430 8892 12854
rect 8956 12434 8984 18158
rect 9416 18086 9444 22510
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9404 18080 9456 18086
rect 9508 18057 9536 25230
rect 9600 24750 9628 27950
rect 9692 26994 9720 29038
rect 9784 28762 9812 29446
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9784 27674 9812 28698
rect 9864 28144 9916 28150
rect 9864 28086 9916 28092
rect 9772 27668 9824 27674
rect 9772 27610 9824 27616
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9784 27130 9812 27406
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9692 26518 9720 26930
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9876 25158 9904 28086
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9600 24614 9628 24686
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9692 18630 9720 24822
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9404 18022 9456 18028
rect 9494 18048 9550 18057
rect 9324 17610 9352 18022
rect 9494 17983 9550 17992
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9048 16454 9076 17546
rect 9416 16726 9444 17750
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9692 17354 9720 17546
rect 9600 17338 9720 17354
rect 9600 17332 9732 17338
rect 9600 17326 9680 17332
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9048 14618 9076 15642
rect 9232 15570 9260 16458
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9048 12918 9076 14554
rect 9232 13870 9260 15506
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9128 13320 9180 13326
rect 9126 13288 9128 13297
rect 9180 13288 9182 13297
rect 9126 13223 9182 13232
rect 9232 12986 9260 13806
rect 9324 13530 9352 14282
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9416 13410 9444 16662
rect 9600 16572 9628 17326
rect 9680 17274 9732 17280
rect 9784 17270 9812 19382
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 16697 9720 17138
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9600 16544 9720 16572
rect 9692 14482 9720 16544
rect 9784 15434 9812 16934
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9772 14952 9824 14958
rect 9770 14920 9772 14929
rect 9824 14920 9826 14929
rect 9770 14855 9826 14864
rect 9876 14600 9904 24346
rect 10336 23866 10364 36722
rect 10520 26382 10548 37130
rect 10704 36922 10732 37130
rect 10968 37120 11020 37126
rect 10968 37062 11020 37068
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10980 31890 11008 37062
rect 11624 36922 11652 39200
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 12268 37210 12296 39200
rect 12992 37256 13044 37262
rect 11612 36916 11664 36922
rect 11612 36858 11664 36864
rect 12176 35894 12204 37198
rect 12268 37182 12480 37210
rect 12992 37198 13044 37204
rect 12452 37126 12480 37182
rect 12440 37120 12492 37126
rect 12440 37062 12492 37068
rect 12900 36712 12952 36718
rect 12900 36654 12952 36660
rect 12176 35866 12296 35894
rect 10968 31884 11020 31890
rect 10968 31826 11020 31832
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10704 29850 10732 30670
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 11612 30660 11664 30666
rect 11612 30602 11664 30608
rect 11072 30394 11100 30602
rect 11060 30388 11112 30394
rect 11060 30330 11112 30336
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 10704 27130 10732 27950
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10612 24750 10640 26454
rect 10704 25294 10732 26930
rect 10796 26790 10824 27338
rect 10888 26994 10916 28698
rect 10980 27538 11008 29582
rect 11164 29170 11192 29718
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 10968 27532 11020 27538
rect 10968 27474 11020 27480
rect 11072 27130 11100 28494
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10796 26586 10824 26726
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10704 24954 10732 25230
rect 10692 24948 10744 24954
rect 10692 24890 10744 24896
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10612 24410 10640 24686
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9968 22098 9996 23598
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10152 22574 10180 23258
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 10152 22098 10180 22510
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10152 21146 10180 21898
rect 10244 21690 10272 22646
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10336 21894 10364 22374
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10322 21720 10378 21729
rect 10232 21684 10284 21690
rect 10322 21655 10378 21664
rect 10232 21626 10284 21632
rect 10336 21554 10364 21655
rect 10520 21554 10548 23666
rect 10612 22710 10640 24006
rect 10796 23594 10824 26318
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10876 25764 10928 25770
rect 10876 25706 10928 25712
rect 10888 25498 10916 25706
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10980 25294 11008 25774
rect 11164 25702 11192 29106
rect 11242 26480 11298 26489
rect 11242 26415 11298 26424
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10784 23588 10836 23594
rect 10784 23530 10836 23536
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10796 23118 10824 23190
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10520 20806 10548 21490
rect 10704 20874 10732 21558
rect 10784 21412 10836 21418
rect 10784 21354 10836 21360
rect 10692 20868 10744 20874
rect 10692 20810 10744 20816
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10152 18970 10180 19382
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10152 16046 10180 18022
rect 10612 17678 10640 18022
rect 10600 17672 10652 17678
rect 10598 17640 10600 17649
rect 10652 17640 10654 17649
rect 10598 17575 10654 17584
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10244 16425 10272 16458
rect 10230 16416 10286 16425
rect 10230 16351 10286 16360
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10140 16040 10192 16046
rect 10138 16008 10140 16017
rect 10192 16008 10194 16017
rect 10138 15943 10194 15952
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15065 9996 15506
rect 10140 15088 10192 15094
rect 9954 15056 10010 15065
rect 10010 15014 10088 15042
rect 10140 15030 10192 15036
rect 9954 14991 10010 15000
rect 10060 14618 10088 15014
rect 9784 14572 9904 14600
rect 10048 14612 10100 14618
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9508 13530 9536 13942
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9416 13382 9536 13410
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9126 12880 9182 12889
rect 9126 12815 9128 12824
rect 9180 12815 9182 12824
rect 9128 12786 9180 12792
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 8956 12406 9076 12434
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8850 7576 8906 7585
rect 8850 7511 8906 7520
rect 8758 6896 8814 6905
rect 8758 6831 8814 6840
rect 8772 6390 8800 6831
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8758 6080 8814 6089
rect 8758 6015 8814 6024
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8680 4486 8708 5782
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8772 4298 8800 6015
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8680 4270 8800 4298
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8036 3726 8156 3754
rect 8128 3670 8156 3726
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8588 3398 8616 4218
rect 8680 3505 8708 4270
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3602 8800 3878
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8666 3496 8722 3505
rect 8666 3431 8722 3440
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8864 3126 8892 7511
rect 8956 4690 8984 8978
rect 9048 8906 9076 12406
rect 9310 11928 9366 11937
rect 9310 11863 9366 11872
rect 9324 11626 9352 11863
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 9738 9168 11086
rect 9416 10810 9444 12582
rect 9508 11801 9536 13382
rect 9600 12646 9628 13806
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9692 12434 9720 14418
rect 9600 12406 9720 12434
rect 9600 12306 9628 12406
rect 9678 12336 9734 12345
rect 9588 12300 9640 12306
rect 9678 12271 9680 12280
rect 9588 12242 9640 12248
rect 9732 12271 9734 12280
rect 9680 12242 9732 12248
rect 9678 12200 9734 12209
rect 9784 12186 9812 14572
rect 10048 14554 10100 14560
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10060 13326 10088 14010
rect 10152 13530 10180 15030
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9784 12158 9904 12186
rect 9678 12135 9734 12144
rect 9692 11830 9720 12135
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 11898 9812 12038
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9680 11824 9732 11830
rect 9494 11792 9550 11801
rect 9680 11766 9732 11772
rect 9494 11727 9550 11736
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9140 9710 9260 9738
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 7274 9076 8842
rect 9140 7750 9168 9590
rect 9232 7954 9260 9710
rect 9416 9518 9444 9998
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9110 9444 9454
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9416 8498 9444 9046
rect 9508 8786 9536 11727
rect 9680 11620 9732 11626
rect 9732 11580 9812 11608
rect 9680 11562 9732 11568
rect 9678 10704 9734 10713
rect 9678 10639 9734 10648
rect 9692 10606 9720 10639
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 8906 9628 10406
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9508 8758 9628 8786
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9310 8392 9366 8401
rect 9310 8327 9366 8336
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9140 6118 9168 7686
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9232 5658 9260 7890
rect 9324 6905 9352 8327
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 7342 9444 7822
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9310 6896 9366 6905
rect 9416 6866 9444 7278
rect 9310 6831 9312 6840
rect 9364 6831 9366 6840
rect 9404 6860 9456 6866
rect 9312 6802 9364 6808
rect 9404 6802 9456 6808
rect 9324 6771 9352 6802
rect 9416 6458 9444 6802
rect 9494 6488 9550 6497
rect 9404 6452 9456 6458
rect 9494 6423 9496 6432
rect 9404 6394 9456 6400
rect 9548 6423 9550 6432
rect 9496 6394 9548 6400
rect 9416 5778 9444 6394
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9232 5630 9536 5658
rect 9036 5296 9088 5302
rect 9128 5296 9180 5302
rect 9036 5238 9088 5244
rect 9126 5264 9128 5273
rect 9180 5264 9182 5273
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8942 4176 8998 4185
rect 8942 4111 8944 4120
rect 8996 4111 8998 4120
rect 8944 4082 8996 4088
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 7654 2751 7710 2760
rect 7760 2746 7972 2774
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 6932 2366 7144 2394
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 2038 6960 2246
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 7116 800 7144 2366
rect 7760 800 7788 2746
rect 9048 800 9076 5238
rect 9126 5199 9182 5208
rect 9140 4434 9168 5199
rect 9220 5160 9272 5166
rect 9404 5160 9456 5166
rect 9220 5102 9272 5108
rect 9402 5128 9404 5137
rect 9456 5128 9458 5137
rect 9232 4554 9260 5102
rect 9402 5063 9458 5072
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9140 4406 9260 4434
rect 9232 3602 9260 4406
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9324 3194 9352 3402
rect 9402 3224 9458 3233
rect 9312 3188 9364 3194
rect 9402 3159 9404 3168
rect 9312 3130 9364 3136
rect 9456 3159 9458 3168
rect 9404 3130 9456 3136
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9324 2514 9352 2926
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9416 2650 9444 2790
rect 9508 2774 9536 5630
rect 9600 3466 9628 8758
rect 9692 8294 9720 10542
rect 9784 10441 9812 11580
rect 9876 11014 9904 12158
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9770 10432 9826 10441
rect 9770 10367 9826 10376
rect 9876 10130 9904 10950
rect 9968 10742 9996 12582
rect 10060 12306 10088 13262
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10152 11898 10180 12854
rect 10244 12442 10272 16118
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10244 11898 10272 12271
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10138 11656 10194 11665
rect 10060 11354 10088 11630
rect 10138 11591 10140 11600
rect 10192 11591 10194 11600
rect 10140 11562 10192 11568
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10046 11112 10102 11121
rect 10152 11082 10180 11290
rect 10046 11047 10102 11056
rect 10140 11076 10192 11082
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9784 8634 9812 8842
rect 9876 8673 9904 9687
rect 9968 8906 9996 10542
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9862 8664 9918 8673
rect 9772 8628 9824 8634
rect 9862 8599 9918 8608
rect 9772 8570 9824 8576
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9692 6730 9720 7103
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9784 5896 9812 8366
rect 9876 6730 9904 8599
rect 10060 8276 10088 11047
rect 10140 11018 10192 11024
rect 10152 8430 10180 11018
rect 10230 10976 10286 10985
rect 10230 10911 10286 10920
rect 10244 10606 10272 10911
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10230 8936 10286 8945
rect 10230 8871 10286 8880
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 9954 8256 10010 8265
rect 10060 8248 10180 8276
rect 9954 8191 10010 8200
rect 9968 7478 9996 8191
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9876 6474 9904 6666
rect 9876 6446 9996 6474
rect 9968 6390 9996 6446
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9784 5868 9996 5896
rect 9770 5808 9826 5817
rect 9770 5743 9772 5752
rect 9824 5743 9826 5752
rect 9772 5714 9824 5720
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 4690 9720 5510
rect 9784 4826 9812 5714
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4826 9904 4966
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9600 2990 9628 3402
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9968 2774 9996 5868
rect 10048 3596 10100 3602
rect 10152 3584 10180 8248
rect 10244 5642 10272 8871
rect 10336 6390 10364 16186
rect 10428 14090 10456 16934
rect 10520 16046 10548 17206
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10428 14062 10548 14090
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10428 7478 10456 13942
rect 10520 12481 10548 14062
rect 10506 12472 10562 12481
rect 10506 12407 10562 12416
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10520 10577 10548 12242
rect 10612 11665 10640 16458
rect 10704 14958 10732 20810
rect 10796 16182 10824 21354
rect 10980 19786 11008 25230
rect 11256 24274 11284 26415
rect 11348 26382 11376 29106
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11532 28490 11560 28902
rect 11428 28484 11480 28490
rect 11428 28426 11480 28432
rect 11520 28484 11572 28490
rect 11520 28426 11572 28432
rect 11440 28082 11468 28426
rect 11428 28076 11480 28082
rect 11428 28018 11480 28024
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11060 24132 11112 24138
rect 11060 24074 11112 24080
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11072 23798 11100 24074
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 11256 23322 11284 24074
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11164 21622 11192 21898
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11256 21418 11284 22646
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10980 19514 11008 19722
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11164 18698 11192 20742
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 17270 10916 17478
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10980 16726 11008 17138
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10796 11830 10824 16118
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10506 10568 10562 10577
rect 10506 10503 10562 10512
rect 10506 9616 10562 9625
rect 10506 9551 10562 9560
rect 10520 7818 10548 9551
rect 10598 9344 10654 9353
rect 10598 9279 10654 9288
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10612 7698 10640 9279
rect 10520 7670 10640 7698
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10100 3556 10180 3584
rect 10048 3538 10100 3544
rect 9508 2746 9628 2774
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9600 2378 9628 2746
rect 9692 2746 9996 2774
rect 10520 2774 10548 7670
rect 10598 6760 10654 6769
rect 10704 6730 10732 11562
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10598 6695 10600 6704
rect 10652 6695 10654 6704
rect 10692 6724 10744 6730
rect 10600 6666 10652 6672
rect 10692 6666 10744 6672
rect 10690 6352 10746 6361
rect 10690 6287 10746 6296
rect 10704 6186 10732 6287
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10796 5148 10824 10746
rect 10888 8906 10916 13262
rect 10980 9654 11008 16390
rect 11072 13433 11100 16934
rect 11058 13424 11114 13433
rect 11058 13359 11114 13368
rect 11058 12064 11114 12073
rect 11058 11999 11114 12008
rect 11072 11626 11100 11999
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11058 11384 11114 11393
rect 11058 11319 11114 11328
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 8945 11008 9318
rect 10966 8936 11022 8945
rect 10876 8900 10928 8906
rect 10966 8871 11022 8880
rect 10876 8842 10928 8848
rect 10874 8800 10930 8809
rect 10874 8735 10930 8744
rect 10888 7188 10916 8735
rect 11072 8022 11100 11319
rect 11164 9908 11192 18090
rect 11256 11354 11284 18634
rect 11348 15473 11376 26318
rect 11440 24410 11468 28018
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11532 18426 11560 27270
rect 11624 23730 11652 30602
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12176 30138 12204 30194
rect 12084 30110 12204 30138
rect 11888 28960 11940 28966
rect 11808 28908 11888 28914
rect 11808 28902 11940 28908
rect 11808 28886 11928 28902
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11716 24857 11744 28018
rect 11808 26382 11836 28886
rect 12084 28082 12112 30110
rect 12268 29034 12296 35866
rect 12808 30796 12860 30802
rect 12808 30738 12860 30744
rect 12256 29028 12308 29034
rect 12256 28970 12308 28976
rect 12440 28484 12492 28490
rect 12440 28426 12492 28432
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 11992 26858 12020 27814
rect 12176 26994 12204 27814
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12268 27062 12296 27406
rect 12256 27056 12308 27062
rect 12256 26998 12308 27004
rect 12348 27056 12400 27062
rect 12348 26998 12400 27004
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 11980 26852 12032 26858
rect 11980 26794 12032 26800
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11702 24848 11758 24857
rect 11702 24783 11758 24792
rect 11612 23724 11664 23730
rect 11612 23666 11664 23672
rect 11624 19922 11652 23666
rect 11808 23118 11836 26318
rect 11888 25832 11940 25838
rect 11888 25774 11940 25780
rect 11900 25498 11928 25774
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11992 25362 12020 26794
rect 12360 26518 12388 26998
rect 12348 26512 12400 26518
rect 12348 26454 12400 26460
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 11980 25152 12032 25158
rect 12360 25106 12388 25638
rect 12452 25378 12480 28426
rect 12716 28008 12768 28014
rect 12716 27950 12768 27956
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12544 25974 12572 27338
rect 12728 26450 12756 27950
rect 12820 26489 12848 30738
rect 12912 28558 12940 36654
rect 13004 30938 13032 37198
rect 13360 37188 13412 37194
rect 13360 37130 13412 37136
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 13372 29646 13400 37130
rect 13556 37126 13584 39200
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 14200 36786 14228 39200
rect 15488 37330 15516 39200
rect 15476 37324 15528 37330
rect 15476 37266 15528 37272
rect 16132 37262 16160 39200
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 16120 37256 16172 37262
rect 16120 37198 16172 37204
rect 14188 36780 14240 36786
rect 14188 36722 14240 36728
rect 15764 36378 15792 37198
rect 16776 36786 16804 39200
rect 16856 37324 16908 37330
rect 16856 37266 16908 37272
rect 16764 36780 16816 36786
rect 16764 36722 16816 36728
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 16120 36100 16172 36106
rect 16120 36042 16172 36048
rect 14464 31952 14516 31958
rect 14464 31894 14516 31900
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13832 30326 13860 31282
rect 14476 31278 14504 31894
rect 14740 31816 14792 31822
rect 14740 31758 14792 31764
rect 14464 31272 14516 31278
rect 14464 31214 14516 31220
rect 14476 30326 14504 31214
rect 13820 30320 13872 30326
rect 13820 30262 13872 30268
rect 14464 30320 14516 30326
rect 14464 30262 14516 30268
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13636 29572 13688 29578
rect 13636 29514 13688 29520
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12806 26480 12862 26489
rect 12716 26444 12768 26450
rect 12912 26450 12940 28358
rect 13176 28008 13228 28014
rect 13176 27950 13228 27956
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 12806 26415 12862 26424
rect 12900 26444 12952 26450
rect 12716 26386 12768 26392
rect 12900 26386 12952 26392
rect 12808 26308 12860 26314
rect 12808 26250 12860 26256
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12452 25350 12572 25378
rect 11980 25094 12032 25100
rect 11992 24562 12020 25094
rect 12268 25078 12388 25106
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 11992 24534 12112 24562
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11704 23044 11756 23050
rect 11704 22986 11756 22992
rect 11716 22166 11744 22986
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 11716 21962 11744 22102
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11716 21690 11744 21898
rect 11808 21690 11836 21898
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11716 21457 11744 21490
rect 11702 21448 11758 21457
rect 11702 21383 11758 21392
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11716 19786 11744 20198
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11808 19446 11836 21286
rect 11992 19446 12020 24346
rect 12084 24138 12112 24534
rect 12176 24342 12204 24822
rect 12164 24336 12216 24342
rect 12164 24278 12216 24284
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 21418 12112 23462
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 12176 18358 12204 22374
rect 12268 19334 12296 25078
rect 12544 24274 12572 25350
rect 12348 24268 12400 24274
rect 12532 24268 12584 24274
rect 12400 24228 12480 24256
rect 12348 24210 12400 24216
rect 12348 22160 12400 22166
rect 12348 22102 12400 22108
rect 12360 20262 12388 22102
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12346 19952 12402 19961
rect 12346 19887 12348 19896
rect 12400 19887 12402 19896
rect 12348 19858 12400 19864
rect 12268 19306 12388 19334
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 17134 11468 17614
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11440 16590 11468 17070
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11440 16153 11468 16526
rect 11426 16144 11482 16153
rect 11426 16079 11482 16088
rect 11334 15464 11390 15473
rect 11334 15399 11390 15408
rect 11532 12617 11560 17478
rect 11716 17338 11744 17750
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11808 17134 11836 17546
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16561 11836 17070
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12268 16794 12296 17002
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 16584 12216 16590
rect 11794 16552 11850 16561
rect 12164 16526 12216 16532
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 11794 16487 11850 16496
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11518 12608 11574 12617
rect 11518 12543 11574 12552
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11348 11082 11376 12378
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11532 10962 11560 12174
rect 11440 10934 11560 10962
rect 11334 10840 11390 10849
rect 11334 10775 11390 10784
rect 11244 9920 11296 9926
rect 11164 9880 11244 9908
rect 11244 9862 11296 9868
rect 11256 8634 11284 9862
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11150 8528 11206 8537
rect 11150 8463 11206 8472
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11072 7342 11100 7958
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10888 7160 11100 7188
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6322 11008 6734
rect 11072 6338 11100 7160
rect 11164 6458 11192 8463
rect 11348 7886 11376 10775
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11256 7478 11284 7686
rect 11348 7546 11376 7686
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11334 6488 11390 6497
rect 11152 6452 11204 6458
rect 11334 6423 11390 6432
rect 11152 6394 11204 6400
rect 10968 6316 11020 6322
rect 11072 6310 11284 6338
rect 10968 6258 11020 6264
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 5160 11020 5166
rect 10796 5120 10968 5148
rect 10968 5102 11020 5108
rect 10980 4457 11008 5102
rect 11072 5030 11100 5510
rect 11256 5386 11284 6310
rect 11348 6118 11376 6423
rect 11440 6390 11468 10934
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9500 11560 9998
rect 11624 9654 11652 13670
rect 11808 13002 11836 16390
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12084 15450 12112 16118
rect 12176 15570 12204 16526
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12268 15502 12296 16526
rect 11900 15422 12112 15450
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11900 14074 11928 15422
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11808 12974 11928 13002
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12753 11744 12786
rect 11702 12744 11758 12753
rect 11702 12679 11758 12688
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11716 12170 11744 12271
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11716 11354 11744 11863
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11900 9602 11928 12974
rect 11992 12442 12020 14486
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11978 12200 12034 12209
rect 11978 12135 11980 12144
rect 12032 12135 12034 12144
rect 11980 12106 12032 12112
rect 12084 11830 12112 15302
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11992 10266 12020 10746
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11978 10024 12034 10033
rect 11978 9959 11980 9968
rect 12032 9959 12034 9968
rect 11980 9930 12032 9936
rect 11900 9574 12020 9602
rect 11704 9512 11756 9518
rect 11532 9472 11704 9500
rect 11756 9472 11836 9500
rect 11704 9454 11756 9460
rect 11808 9042 11836 9472
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 8809 11560 8842
rect 11518 8800 11574 8809
rect 11518 8735 11574 8744
rect 11808 8498 11836 8978
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11440 5846 11468 6326
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11426 5672 11482 5681
rect 11426 5607 11482 5616
rect 11256 5358 11376 5386
rect 11060 5024 11112 5030
rect 11112 4984 11192 5012
rect 11060 4966 11112 4972
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10966 4448 11022 4457
rect 10966 4383 11022 4392
rect 11072 4078 11100 4558
rect 10784 4072 10836 4078
rect 10782 4040 10784 4049
rect 11060 4072 11112 4078
rect 10836 4040 10838 4049
rect 11060 4014 11112 4020
rect 10782 3975 10838 3984
rect 10796 2961 10824 3975
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10888 3126 10916 3606
rect 11072 3534 11100 4014
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 11072 3058 11100 3470
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2984 11020 2990
rect 10782 2952 10838 2961
rect 10968 2926 11020 2932
rect 10782 2887 10838 2896
rect 10980 2825 11008 2926
rect 10966 2816 11022 2825
rect 10520 2746 10732 2774
rect 10966 2751 11022 2760
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9600 1834 9628 2314
rect 9588 1828 9640 1834
rect 9588 1770 9640 1776
rect 9692 800 9720 2746
rect 10704 2038 10732 2746
rect 11072 2514 11100 2994
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11164 2446 11192 4984
rect 11348 3466 11376 5358
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 10324 2032 10376 2038
rect 10324 1974 10376 1980
rect 10692 2032 10744 2038
rect 10692 1974 10744 1980
rect 10336 800 10364 1974
rect 11348 1698 11376 3402
rect 11440 2854 11468 5607
rect 11532 5216 11560 7822
rect 11624 7177 11652 8434
rect 11900 8294 11928 8502
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11610 7168 11666 7177
rect 11610 7103 11666 7112
rect 11716 6866 11744 7822
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 7206 11836 7346
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11886 7032 11942 7041
rect 11886 6967 11888 6976
rect 11940 6967 11942 6976
rect 11888 6938 11940 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 5846 11652 6598
rect 11716 6322 11744 6802
rect 11992 6730 12020 9574
rect 12084 8922 12112 11494
rect 12176 10554 12204 14214
rect 12268 11082 12296 15302
rect 12360 13954 12388 19306
rect 12452 17134 12480 24228
rect 12532 24210 12584 24216
rect 12530 21584 12586 21593
rect 12530 21519 12532 21528
rect 12584 21519 12586 21528
rect 12532 21490 12584 21496
rect 12532 21072 12584 21078
rect 12532 21014 12584 21020
rect 12544 19310 12572 21014
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12636 18970 12664 25978
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12728 21622 12756 24754
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12820 20602 12848 26250
rect 12912 26081 12940 26386
rect 12898 26072 12954 26081
rect 12898 26007 12954 26016
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 13004 25158 13032 25978
rect 13096 25906 13124 26454
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 13096 25809 13124 25842
rect 13082 25800 13138 25809
rect 13082 25735 13138 25744
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 13188 23746 13216 27950
rect 13556 27606 13584 27950
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 13648 27538 13676 29514
rect 14004 29504 14056 29510
rect 14004 29446 14056 29452
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13832 27674 13860 28086
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13740 25498 13768 25638
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13280 24750 13308 25230
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13280 24410 13308 24550
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 12912 23718 13216 23746
rect 12912 23526 12940 23718
rect 12900 23520 12952 23526
rect 12900 23462 12952 23468
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13004 22642 13032 23462
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12912 21078 12940 22102
rect 13004 22030 13032 22578
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 13096 21486 13124 21898
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 13096 20534 13124 21422
rect 13280 20534 13308 24210
rect 13372 22710 13400 24550
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 13464 22094 13492 24754
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13740 22778 13768 24142
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23798 13860 24006
rect 13820 23792 13872 23798
rect 13820 23734 13872 23740
rect 13924 23322 13952 28018
rect 14016 26926 14044 29446
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14464 28484 14516 28490
rect 14464 28426 14516 28432
rect 14188 28416 14240 28422
rect 14188 28358 14240 28364
rect 14372 28416 14424 28422
rect 14372 28358 14424 28364
rect 14096 27396 14148 27402
rect 14096 27338 14148 27344
rect 14108 26994 14136 27338
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 14016 23202 14044 24754
rect 14108 23254 14136 25434
rect 14200 25430 14228 28358
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14188 25424 14240 25430
rect 14188 25366 14240 25372
rect 14200 25226 14228 25366
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 13924 23174 14044 23202
rect 14096 23248 14148 23254
rect 14096 23190 14148 23196
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13740 22681 13768 22714
rect 13726 22672 13782 22681
rect 13726 22607 13782 22616
rect 13372 22066 13492 22094
rect 13820 22092 13872 22098
rect 13372 21593 13400 22066
rect 13820 22034 13872 22040
rect 13452 22024 13504 22030
rect 13504 21984 13584 22012
rect 13452 21966 13504 21972
rect 13358 21584 13414 21593
rect 13358 21519 13414 21528
rect 13372 20777 13400 21519
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13464 20942 13492 21014
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13358 20768 13414 20777
rect 13358 20703 13414 20712
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12714 19952 12770 19961
rect 12714 19887 12770 19896
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12728 18358 12756 19887
rect 12912 19378 12940 20402
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12806 18184 12862 18193
rect 12806 18119 12862 18128
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16794 12756 17070
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12452 14414 12480 15438
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12360 13926 12480 13954
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12360 12186 12388 13806
rect 12452 12889 12480 13926
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 13530 12572 13738
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12438 12880 12494 12889
rect 12438 12815 12494 12824
rect 12544 12306 12572 12922
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12360 12170 12480 12186
rect 12360 12164 12492 12170
rect 12360 12158 12440 12164
rect 12440 12106 12492 12112
rect 12348 11688 12400 11694
rect 12544 11676 12572 12242
rect 12636 12186 12664 16390
rect 12728 12306 12756 16390
rect 12820 16182 12848 18119
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12636 12158 12756 12186
rect 12400 11648 12572 11676
rect 12624 11688 12676 11694
rect 12622 11656 12624 11665
rect 12676 11656 12678 11665
rect 12348 11630 12400 11636
rect 12452 11354 12480 11648
rect 12622 11591 12678 11600
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12452 10658 12480 11290
rect 12624 10736 12676 10742
rect 12622 10704 12624 10713
rect 12676 10704 12678 10713
rect 12440 10652 12492 10658
rect 12622 10639 12678 10648
rect 12440 10594 12492 10600
rect 12176 10526 12572 10554
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12268 9110 12296 9930
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12084 8906 12296 8922
rect 12084 8900 12308 8906
rect 12084 8894 12256 8900
rect 12256 8842 12308 8848
rect 12360 8378 12388 10202
rect 12438 9888 12494 9897
rect 12438 9823 12494 9832
rect 12452 9518 12480 9823
rect 12544 9654 12572 10526
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12438 8664 12494 8673
rect 12438 8599 12440 8608
rect 12492 8599 12494 8608
rect 12440 8570 12492 8576
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12176 8350 12388 8378
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7002 12112 7754
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12084 6390 12112 6598
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11716 5778 11744 6258
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5234 11744 5714
rect 11704 5228 11756 5234
rect 11532 5188 11652 5216
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4554 11560 5034
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11624 4486 11652 5188
rect 11704 5170 11756 5176
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11336 1692 11388 1698
rect 11336 1634 11388 1640
rect 11624 800 11652 2858
rect 12176 2774 12204 8350
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12360 8248 12480 8276
rect 12268 7274 12296 8230
rect 12360 7954 12388 8248
rect 12452 7954 12480 8248
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12360 6866 12388 7278
rect 12438 7032 12494 7041
rect 12438 6967 12440 6976
rect 12492 6967 12494 6976
rect 12440 6938 12492 6944
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12084 2746 12204 2774
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11716 1970 11744 2586
rect 12084 2310 12112 2746
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 11704 1964 11756 1970
rect 11704 1906 11756 1912
rect 12268 800 12296 2790
rect 12544 2378 12572 8502
rect 12622 6896 12678 6905
rect 12622 6831 12678 6840
rect 12636 5302 12664 6831
rect 12728 5642 12756 12158
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12820 4554 12848 15846
rect 12912 14929 12940 18294
rect 13004 17610 13032 19654
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13096 16454 13124 20470
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13188 19514 13216 19926
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13280 17921 13308 19450
rect 13266 17912 13322 17921
rect 13266 17847 13322 17856
rect 13372 17082 13400 20402
rect 13188 17054 13400 17082
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12990 16144 13046 16153
rect 12990 16079 12992 16088
rect 13044 16079 13046 16088
rect 12992 16050 13044 16056
rect 12898 14920 12954 14929
rect 12898 14855 12954 14864
rect 12912 14822 12940 14855
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12898 14512 12954 14521
rect 12898 14447 12954 14456
rect 12912 14414 12940 14447
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12898 14240 12954 14249
rect 12898 14175 12954 14184
rect 12912 13274 12940 14175
rect 13004 13938 13032 16050
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13096 13870 13124 14894
rect 13188 13954 13216 17054
rect 13464 16726 13492 20878
rect 13556 18850 13584 21984
rect 13832 21894 13860 22034
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13648 20913 13676 20946
rect 13634 20904 13690 20913
rect 13634 20839 13690 20848
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13648 19553 13676 19790
rect 13634 19544 13690 19553
rect 13634 19479 13690 19488
rect 13556 18822 13676 18850
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 15348 13400 16390
rect 13464 15502 13492 16526
rect 13556 16182 13584 16934
rect 13648 16561 13676 18822
rect 13924 18358 13952 23174
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14108 20890 14136 23054
rect 14108 20862 14228 20890
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 16658 13768 17478
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13634 16552 13690 16561
rect 13634 16487 13690 16496
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 16250 13676 16390
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15910 13676 16050
rect 13636 15904 13688 15910
rect 13832 15858 13860 16662
rect 13636 15846 13688 15852
rect 13740 15830 13860 15858
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13372 15320 13492 15348
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13280 14249 13308 14350
rect 13266 14240 13322 14249
rect 13266 14175 13322 14184
rect 13360 14000 13412 14006
rect 13188 13926 13308 13954
rect 13360 13942 13412 13948
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12992 13388 13044 13394
rect 13096 13376 13124 13806
rect 13044 13348 13124 13376
rect 12992 13330 13044 13336
rect 12912 13246 13032 13274
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12912 8566 12940 12543
rect 13004 12434 13032 13246
rect 13096 12986 13124 13348
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13082 12880 13138 12889
rect 13082 12815 13138 12824
rect 13096 12782 13124 12815
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13280 12434 13308 13926
rect 13372 13462 13400 13942
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13004 12406 13124 12434
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 13004 7818 13032 12242
rect 13096 10062 13124 12406
rect 13188 12406 13308 12434
rect 13464 12434 13492 15320
rect 13634 13560 13690 13569
rect 13634 13495 13690 13504
rect 13648 13326 13676 13495
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13464 12406 13584 12434
rect 13188 10606 13216 12406
rect 13358 12336 13414 12345
rect 13358 12271 13414 12280
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13188 9382 13216 10542
rect 13280 10062 13308 11630
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13372 9874 13400 12271
rect 13450 10704 13506 10713
rect 13450 10639 13506 10648
rect 13464 10606 13492 10639
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13280 9846 13400 9874
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8022 13124 8842
rect 13176 8832 13228 8838
rect 13174 8800 13176 8809
rect 13228 8800 13230 8809
rect 13174 8735 13230 8744
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12992 7812 13044 7818
rect 12992 7754 13044 7760
rect 13082 6896 13138 6905
rect 13082 6831 13138 6840
rect 13096 6798 13124 6831
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13280 5302 13308 9846
rect 13360 8968 13412 8974
rect 13412 8928 13492 8956
rect 13360 8910 13412 8916
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 13372 4078 13400 6734
rect 13464 4214 13492 8928
rect 13556 7954 13584 12406
rect 13634 12336 13690 12345
rect 13634 12271 13636 12280
rect 13688 12271 13690 12280
rect 13636 12242 13688 12248
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 9654 13676 10950
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13740 8906 13768 15830
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 14006 13860 15302
rect 14016 14958 14044 19654
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13924 12434 13952 14418
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 12918 14044 14282
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 13832 12406 13952 12434
rect 13832 10674 13860 12406
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13924 11393 13952 11494
rect 13910 11384 13966 11393
rect 13910 11319 13966 11328
rect 14016 11218 14044 11494
rect 14108 11354 14136 20742
rect 14200 12434 14228 20862
rect 14292 19514 14320 26930
rect 14384 26450 14412 28358
rect 14476 27402 14504 28426
rect 14568 27606 14596 28494
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14568 27282 14596 27542
rect 14476 27254 14596 27282
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14476 26330 14504 27254
rect 14556 27056 14608 27062
rect 14556 26998 14608 27004
rect 14568 26586 14596 26998
rect 14556 26580 14608 26586
rect 14556 26522 14608 26528
rect 14384 26302 14504 26330
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14384 17626 14412 26302
rect 14568 25838 14596 26318
rect 14556 25832 14608 25838
rect 14556 25774 14608 25780
rect 14464 25764 14516 25770
rect 14464 25706 14516 25712
rect 14476 25226 14504 25706
rect 14554 25392 14610 25401
rect 14554 25327 14610 25336
rect 14464 25220 14516 25226
rect 14464 25162 14516 25168
rect 14568 25106 14596 25327
rect 14476 25078 14596 25106
rect 14476 23866 14504 25078
rect 14660 24698 14688 29242
rect 14752 28490 14780 31758
rect 14832 31272 14884 31278
rect 14832 31214 14884 31220
rect 14844 30802 14872 31214
rect 14924 31136 14976 31142
rect 14924 31078 14976 31084
rect 14936 30870 14964 31078
rect 14924 30864 14976 30870
rect 14924 30806 14976 30812
rect 14832 30796 14884 30802
rect 14832 30738 14884 30744
rect 14936 30122 14964 30806
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15108 30184 15160 30190
rect 15108 30126 15160 30132
rect 14924 30116 14976 30122
rect 14924 30058 14976 30064
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 14844 28626 14872 29038
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14740 28484 14792 28490
rect 14740 28426 14792 28432
rect 14844 28218 14872 28562
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14844 26466 14872 26726
rect 14936 26586 14964 30058
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 15028 29170 15056 29990
rect 15120 29714 15148 30126
rect 15396 29850 15424 30670
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 16040 29850 16068 30262
rect 16132 30258 16160 36042
rect 16868 35894 16896 37266
rect 18064 37262 18092 39200
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 17040 36576 17092 36582
rect 17040 36518 17092 36524
rect 16868 35866 16988 35894
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 16304 30116 16356 30122
rect 16304 30058 16356 30064
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 15120 28490 15148 29446
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 15304 28490 15332 28970
rect 15660 28960 15712 28966
rect 15660 28902 15712 28908
rect 15016 28484 15068 28490
rect 15016 28426 15068 28432
rect 15108 28484 15160 28490
rect 15108 28426 15160 28432
rect 15292 28484 15344 28490
rect 15292 28426 15344 28432
rect 15028 27606 15056 28426
rect 15672 28014 15700 28902
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15660 28008 15712 28014
rect 15660 27950 15712 27956
rect 15672 27878 15700 27950
rect 15660 27872 15712 27878
rect 15660 27814 15712 27820
rect 15016 27600 15068 27606
rect 15016 27542 15068 27548
rect 15764 27470 15792 28358
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14844 26438 14964 26466
rect 14660 24670 14780 24698
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14476 22098 14504 22986
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 20262 14504 21422
rect 14568 20398 14596 24278
rect 14660 23798 14688 24550
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 14660 21622 14688 23122
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14660 18902 14688 21558
rect 14752 20942 14780 24670
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14752 19718 14780 20878
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14384 17598 14688 17626
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17105 14412 17478
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14370 17096 14426 17105
rect 14370 17031 14426 17040
rect 14476 16697 14504 17138
rect 14462 16688 14518 16697
rect 14462 16623 14518 16632
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14292 16046 14320 16186
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 15706 14596 15982
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14660 15586 14688 17598
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14568 15558 14688 15586
rect 14292 13258 14320 15506
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14200 12406 14320 12434
rect 14292 11558 14320 12406
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14108 11257 14136 11290
rect 14094 11248 14150 11257
rect 14004 11212 14056 11218
rect 14094 11183 14150 11192
rect 14004 11154 14056 11160
rect 14280 11144 14332 11150
rect 14384 11132 14412 15370
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14476 14521 14504 14962
rect 14462 14512 14518 14521
rect 14462 14447 14518 14456
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 12918 14504 13670
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14332 11104 14412 11132
rect 14280 11086 14332 11092
rect 14292 10810 14320 11086
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14476 10742 14504 12718
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 13818 10568 13874 10577
rect 13818 10503 13874 10512
rect 13832 9674 13860 10503
rect 14002 10432 14058 10441
rect 14002 10367 14058 10376
rect 13832 9646 13952 9674
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13544 7948 13596 7954
rect 13596 7908 13676 7936
rect 13544 7890 13596 7896
rect 13542 7032 13598 7041
rect 13542 6967 13598 6976
rect 13556 6798 13584 6967
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13648 5166 13676 7908
rect 13924 7886 13952 9646
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 7002 13768 7210
rect 13818 7168 13874 7177
rect 13818 7103 13874 7112
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13832 6458 13860 7103
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13726 5400 13782 5409
rect 13726 5335 13782 5344
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13740 4865 13768 5335
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13726 4856 13782 4865
rect 13726 4791 13782 4800
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3194 13032 3878
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12912 2938 12940 3130
rect 12912 2922 13124 2938
rect 12912 2916 13136 2922
rect 12912 2910 13084 2916
rect 13084 2858 13136 2864
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 13556 800 13584 4422
rect 13740 3534 13768 4791
rect 13832 4690 13860 5102
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13924 4593 13952 7822
rect 14016 5001 14044 10367
rect 14094 9888 14150 9897
rect 14094 9823 14150 9832
rect 14108 8362 14136 9823
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14200 6662 14228 9046
rect 14292 8634 14320 9454
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6730 14320 7346
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14108 6254 14136 6598
rect 14292 6458 14320 6666
rect 14280 6452 14332 6458
rect 14200 6412 14280 6440
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14108 5098 14136 5578
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14002 4992 14058 5001
rect 14002 4927 14058 4936
rect 14096 4616 14148 4622
rect 13910 4584 13966 4593
rect 14096 4558 14148 4564
rect 13910 4519 13966 4528
rect 14108 4185 14136 4558
rect 14200 4282 14228 6412
rect 14280 6394 14332 6400
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4622 14320 5102
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14094 4176 14150 4185
rect 14094 4111 14150 4120
rect 14096 3936 14148 3942
rect 14292 3924 14320 4558
rect 14148 3896 14320 3924
rect 14096 3878 14148 3884
rect 14292 3602 14320 3896
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13740 2038 13768 2314
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 14108 1902 14136 3334
rect 14292 3058 14320 3538
rect 14280 3052 14332 3058
rect 14200 3012 14280 3040
rect 14200 2514 14228 3012
rect 14280 2994 14332 3000
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14384 2394 14412 10610
rect 14568 10248 14596 15558
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14476 10220 14596 10248
rect 14476 7478 14504 10220
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14568 9586 14596 10066
rect 14660 9926 14688 14214
rect 14752 11937 14780 19314
rect 14844 17134 14872 20334
rect 14936 17746 14964 26438
rect 15028 25838 15056 26862
rect 15120 26382 15148 27066
rect 15384 26920 15436 26926
rect 15384 26862 15436 26868
rect 15396 26518 15424 26862
rect 15384 26512 15436 26518
rect 15384 26454 15436 26460
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 15016 25832 15068 25838
rect 15016 25774 15068 25780
rect 15120 24682 15148 25910
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 24698 15424 24754
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15212 24670 15424 24698
rect 15212 24562 15240 24670
rect 15120 24534 15240 24562
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15014 24440 15070 24449
rect 15014 24375 15016 24384
rect 15068 24375 15070 24384
rect 15016 24346 15068 24352
rect 15120 24290 15148 24534
rect 15028 24262 15148 24290
rect 15028 22094 15056 24262
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15120 22710 15148 24074
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 15212 22574 15240 23258
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15028 22066 15148 22094
rect 15120 19786 15148 22066
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15212 21486 15240 22034
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15304 20534 15332 24550
rect 15488 22094 15516 27270
rect 15672 25838 15700 27338
rect 15764 26518 15792 27406
rect 15856 27033 15884 29106
rect 16120 28960 16172 28966
rect 16120 28902 16172 28908
rect 16132 28778 16160 28902
rect 16132 28750 16252 28778
rect 16028 28688 16080 28694
rect 16080 28636 16160 28642
rect 16028 28630 16160 28636
rect 16040 28614 16160 28630
rect 16224 28626 16252 28750
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15842 27024 15898 27033
rect 15842 26959 15844 26968
rect 15896 26959 15898 26968
rect 15844 26930 15896 26936
rect 15948 26858 15976 27338
rect 15936 26852 15988 26858
rect 15936 26794 15988 26800
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15752 26512 15804 26518
rect 15752 26454 15804 26460
rect 15856 26330 15884 26726
rect 15764 26302 15884 26330
rect 16040 26314 16068 28358
rect 16028 26308 16080 26314
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15672 23322 15700 25774
rect 15764 25158 15792 26302
rect 16028 26250 16080 26256
rect 16132 25702 16160 28614
rect 16212 28620 16264 28626
rect 16212 28562 16264 28568
rect 16316 28150 16344 30058
rect 16396 28960 16448 28966
rect 16396 28902 16448 28908
rect 16304 28144 16356 28150
rect 16304 28086 16356 28092
rect 16316 27538 16344 28086
rect 16304 27532 16356 27538
rect 16304 27474 16356 27480
rect 16120 25696 16172 25702
rect 16120 25638 16172 25644
rect 16132 25294 16160 25638
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15396 22066 15516 22094
rect 15396 21146 15424 22066
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15016 19712 15068 19718
rect 15212 19666 15240 20334
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15580 19854 15608 19994
rect 15384 19848 15436 19854
rect 15568 19848 15620 19854
rect 15384 19790 15436 19796
rect 15474 19816 15530 19825
rect 15016 19654 15068 19660
rect 15028 19446 15056 19654
rect 15120 19638 15240 19666
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 15120 18358 15148 19638
rect 15396 19378 15424 19790
rect 15568 19790 15620 19796
rect 15474 19751 15476 19760
rect 15528 19751 15530 19760
rect 15476 19722 15528 19728
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14936 15706 14964 16390
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15028 15450 15056 17818
rect 15120 17814 15148 18294
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15212 17270 15240 19314
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15384 17808 15436 17814
rect 15384 17750 15436 17756
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16454 15148 16934
rect 15304 16697 15332 17478
rect 15290 16688 15346 16697
rect 15290 16623 15346 16632
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15212 15570 15240 16526
rect 15396 16425 15424 17750
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15382 16416 15438 16425
rect 15382 16351 15438 16360
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 14936 15422 15056 15450
rect 14936 14906 14964 15422
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14844 14878 14964 14906
rect 14844 13870 14872 14878
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14844 13297 14872 13806
rect 14830 13288 14886 13297
rect 14830 13223 14886 13232
rect 14830 12472 14886 12481
rect 14830 12407 14886 12416
rect 14738 11928 14794 11937
rect 14738 11863 14794 11872
rect 14844 11830 14872 12407
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14556 9580 14608 9586
rect 14608 9540 14688 9568
rect 14556 9522 14608 9528
rect 14556 9036 14608 9042
rect 14660 9024 14688 9540
rect 14608 8996 14688 9024
rect 14556 8978 14608 8984
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 8809 14596 8842
rect 14554 8800 14610 8809
rect 14554 8735 14610 8744
rect 14568 8294 14596 8735
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14660 7886 14688 8996
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14660 7478 14688 7822
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14476 7002 14504 7414
rect 14752 7313 14780 11766
rect 14936 11082 14964 14758
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14830 10976 14886 10985
rect 14830 10911 14886 10920
rect 14844 9654 14872 10911
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 14924 9376 14976 9382
rect 14830 9344 14886 9353
rect 14924 9318 14976 9324
rect 14830 9279 14886 9288
rect 14738 7304 14794 7313
rect 14738 7239 14794 7248
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14752 6322 14780 7142
rect 14844 6390 14872 9279
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5574 14780 6258
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14568 2774 14596 5238
rect 14646 4312 14702 4321
rect 14646 4247 14702 4256
rect 14660 3466 14688 4247
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14844 3126 14872 6054
rect 14936 4214 14964 9318
rect 15028 8906 15056 15302
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15120 14006 15148 14894
rect 15212 14414 15240 15506
rect 15384 15428 15436 15434
rect 15488 15416 15516 17614
rect 15580 15586 15608 18702
rect 15672 18426 15700 22646
rect 15764 22094 15792 25094
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 24274 15976 24550
rect 15936 24268 15988 24274
rect 15936 24210 15988 24216
rect 15844 24064 15896 24070
rect 15844 24006 15896 24012
rect 15856 23032 15884 24006
rect 15948 23662 15976 24210
rect 16040 24138 16068 25094
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 15948 23186 15976 23598
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 15936 23044 15988 23050
rect 15856 23004 15936 23032
rect 15936 22986 15988 22992
rect 16408 22094 16436 28902
rect 16592 25378 16620 31282
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16776 28558 16804 29514
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 16868 28218 16896 28358
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16960 28082 16988 35866
rect 17052 29646 17080 36518
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 17144 31414 17172 33798
rect 17132 31408 17184 31414
rect 17132 31350 17184 31356
rect 17316 30048 17368 30054
rect 17316 29990 17368 29996
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 17328 28762 17356 29990
rect 18616 29850 18644 37198
rect 18708 37126 18736 39200
rect 19996 37346 20024 39200
rect 19432 37324 19484 37330
rect 19996 37318 20116 37346
rect 19432 37266 19484 37272
rect 18696 37120 18748 37126
rect 18696 37062 18748 37068
rect 18880 36780 18932 36786
rect 18880 36722 18932 36728
rect 18892 30326 18920 36722
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19352 32502 19380 32710
rect 19340 32496 19392 32502
rect 19340 32438 19392 32444
rect 18880 30320 18932 30326
rect 18880 30262 18932 30268
rect 18604 29844 18656 29850
rect 18604 29786 18656 29792
rect 18234 29744 18290 29753
rect 18234 29679 18290 29688
rect 18248 29646 18276 29679
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18696 29504 18748 29510
rect 18696 29446 18748 29452
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17776 28484 17828 28490
rect 17776 28426 17828 28432
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 16960 27962 16988 28018
rect 17788 28014 17816 28426
rect 17868 28144 17920 28150
rect 17868 28086 17920 28092
rect 16868 27934 16988 27962
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 16868 27674 16896 27934
rect 16948 27872 17000 27878
rect 16948 27814 17000 27820
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16500 25350 16620 25378
rect 16500 24954 16528 25350
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23089 16528 23530
rect 16486 23080 16542 23089
rect 16486 23015 16542 23024
rect 16592 22982 16620 25162
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 15764 22066 15884 22094
rect 16408 22066 16528 22094
rect 15856 21486 15884 22066
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16316 21690 16344 21898
rect 16394 21720 16450 21729
rect 16304 21684 16356 21690
rect 16394 21655 16396 21664
rect 16304 21626 16356 21632
rect 16448 21655 16450 21664
rect 16396 21626 16448 21632
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15948 20992 15976 21490
rect 15764 20964 15976 20992
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15672 16969 15700 17070
rect 15658 16960 15714 16969
rect 15658 16895 15714 16904
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 16250 15700 16458
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15580 15558 15700 15586
rect 15436 15388 15516 15416
rect 15384 15370 15436 15376
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 14074 15332 14214
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 13326 15240 13670
rect 15396 13530 15424 15030
rect 15488 15026 15516 15388
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15488 13326 15516 14350
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15476 13320 15528 13326
rect 15580 13297 15608 15302
rect 15476 13262 15528 13268
rect 15566 13288 15622 13297
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15212 11558 15240 12242
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 11144 15160 11150
rect 15160 11092 15240 11098
rect 15108 11086 15240 11092
rect 15120 11070 15240 11086
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15028 5642 15056 6258
rect 15120 6118 15148 6666
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15106 5400 15162 5409
rect 15106 5335 15162 5344
rect 15120 5302 15148 5335
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 15106 4992 15162 5001
rect 15106 4927 15162 4936
rect 15120 4554 15148 4927
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15106 4312 15162 4321
rect 15106 4247 15162 4256
rect 15120 4214 15148 4247
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15212 3466 15240 11070
rect 15304 9994 15332 13262
rect 15566 13223 15622 13232
rect 15672 12322 15700 15558
rect 15396 12294 15700 12322
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15290 8392 15346 8401
rect 15290 8327 15346 8336
rect 15304 7954 15332 8327
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 5522 15332 7890
rect 15396 6934 15424 12294
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15672 11898 15700 12106
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15474 11384 15530 11393
rect 15474 11319 15476 11328
rect 15528 11319 15530 11328
rect 15476 11290 15528 11296
rect 15474 11248 15530 11257
rect 15474 11183 15476 11192
rect 15528 11183 15530 11192
rect 15476 11154 15528 11160
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 10266 15700 10406
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15764 8809 15792 20964
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15948 20058 15976 20810
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15844 19984 15896 19990
rect 15842 19952 15844 19961
rect 15896 19952 15898 19961
rect 15842 19887 15898 19896
rect 16132 18766 16160 20402
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 19378 16436 20198
rect 16304 19372 16356 19378
rect 16304 19314 16356 19320
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16040 17542 16068 18566
rect 16132 17678 16160 18566
rect 16120 17672 16172 17678
rect 16172 17632 16252 17660
rect 16120 17614 16172 17620
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15856 16697 15884 17478
rect 16224 16794 16252 17632
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15842 16688 15898 16697
rect 15842 16623 15898 16632
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16028 16040 16080 16046
rect 15948 16000 16028 16028
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 15162 15884 15438
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15856 14362 15884 15098
rect 15948 14482 15976 16000
rect 16028 15982 16080 15988
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15856 14334 15976 14362
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 12434 15884 14214
rect 15948 13734 15976 14334
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15948 12646 15976 12922
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15856 12406 15976 12434
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 9518 15884 11494
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15842 9208 15898 9217
rect 15842 9143 15898 9152
rect 15750 8800 15806 8809
rect 15750 8735 15806 8744
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15568 7948 15620 7954
rect 15488 7908 15568 7936
rect 15488 7818 15516 7908
rect 15568 7890 15620 7896
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15764 7546 15792 8026
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15304 5494 15424 5522
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14568 2746 14872 2774
rect 14200 2366 14412 2394
rect 14464 2372 14516 2378
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 14200 800 14228 2366
rect 14464 2314 14516 2320
rect 14476 1970 14504 2314
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14844 800 14872 2746
rect 15200 2508 15252 2514
rect 15396 2496 15424 5494
rect 15856 4554 15884 9143
rect 15948 8673 15976 12406
rect 15934 8664 15990 8673
rect 15934 8599 15990 8608
rect 16040 7410 16068 14214
rect 16132 9738 16160 16594
rect 16224 16046 16252 16730
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16212 15360 16264 15366
rect 16210 15328 16212 15337
rect 16264 15328 16266 15337
rect 16210 15263 16266 15272
rect 16316 14278 16344 19314
rect 16500 17921 16528 22066
rect 16592 18834 16620 22918
rect 16684 21622 16712 24754
rect 16776 24750 16804 27406
rect 16960 27402 16988 27814
rect 17880 27674 17908 28086
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 16948 27396 17000 27402
rect 16948 27338 17000 27344
rect 16960 27062 16988 27338
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 17592 27056 17644 27062
rect 17592 26998 17644 27004
rect 16960 26450 16988 26998
rect 17408 26512 17460 26518
rect 17144 26472 17408 26500
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 17144 25770 17172 26472
rect 17408 26454 17460 26460
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17132 25764 17184 25770
rect 17132 25706 17184 25712
rect 16856 25424 16908 25430
rect 16856 25366 16908 25372
rect 16868 25226 16896 25366
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 17040 25220 17092 25226
rect 17040 25162 17092 25168
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16868 24274 16896 25162
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 17052 24138 17080 25162
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17040 24132 17092 24138
rect 16960 24092 17040 24120
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16868 22094 16896 23462
rect 16960 22166 16988 24092
rect 17040 24074 17092 24080
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 16776 22066 16896 22094
rect 16776 21962 16804 22066
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16776 20262 16804 20470
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16486 17912 16542 17921
rect 16592 17882 16620 18770
rect 16486 17847 16488 17856
rect 16540 17847 16542 17856
rect 16580 17876 16632 17882
rect 16488 17818 16540 17824
rect 16580 17818 16632 17824
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16592 17626 16620 17682
rect 16500 17610 16620 17626
rect 16488 17604 16620 17610
rect 16540 17598 16620 17604
rect 16488 17546 16540 17552
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16408 15502 16436 16662
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 14822 16436 15438
rect 16500 15162 16528 17546
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16500 13938 16528 14350
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16302 13696 16358 13705
rect 16224 13394 16252 13670
rect 16302 13631 16358 13640
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16224 12170 16252 13126
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16132 9710 16252 9738
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16132 9489 16160 9590
rect 16224 9518 16252 9710
rect 16212 9512 16264 9518
rect 16118 9480 16174 9489
rect 16212 9454 16264 9460
rect 16118 9415 16174 9424
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16026 7304 16082 7313
rect 16026 7239 16082 7248
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 16040 3369 16068 7239
rect 16132 6934 16160 8298
rect 16224 8022 16252 9454
rect 16316 8566 16344 13631
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16394 12880 16450 12889
rect 16394 12815 16450 12824
rect 16408 10130 16436 12815
rect 16500 11937 16528 13194
rect 16486 11928 16542 11937
rect 16486 11863 16542 11872
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 8566 16436 10066
rect 16500 9518 16528 10610
rect 16592 9586 16620 14350
rect 16684 11558 16712 19790
rect 16776 16182 16804 20198
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16868 17338 16896 17546
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16868 16017 16896 17138
rect 16960 16794 16988 22102
rect 17052 21146 17080 23666
rect 17144 23186 17172 24686
rect 17236 24154 17264 26250
rect 17328 26042 17356 26250
rect 17604 26042 17632 26998
rect 18708 26926 18736 29446
rect 19444 28694 19472 37266
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19996 36922 20024 37198
rect 20088 37126 20116 37318
rect 20640 37210 20668 39200
rect 21284 37262 21312 39200
rect 21180 37256 21232 37262
rect 20640 37182 20760 37210
rect 21180 37198 21232 37204
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 20732 37126 20760 37182
rect 20076 37120 20128 37126
rect 20076 37062 20128 37068
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20352 35760 20404 35766
rect 20352 35702 20404 35708
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20364 32502 20392 35702
rect 19984 32496 20036 32502
rect 19984 32438 20036 32444
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19352 28082 19380 28494
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 18064 26314 18092 26726
rect 18052 26308 18104 26314
rect 18052 26250 18104 26256
rect 17682 26072 17738 26081
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 17592 26036 17644 26042
rect 17682 26007 17684 26016
rect 17592 25978 17644 25984
rect 17736 26007 17738 26016
rect 17684 25978 17736 25984
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 24449 17356 24686
rect 17314 24440 17370 24449
rect 17314 24375 17370 24384
rect 17236 24126 17356 24154
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17236 21706 17264 22578
rect 17328 22098 17356 24126
rect 17420 23730 17448 25842
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17512 23050 17540 23462
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17420 22234 17448 22986
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 17236 21678 17356 21706
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17144 21146 17172 21286
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 17052 20534 17080 20742
rect 17236 20602 17264 21558
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 17328 19417 17356 21678
rect 17420 21486 17448 21898
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 20058 17540 20810
rect 17604 20806 17632 24686
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17788 23798 17816 24210
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17682 20904 17738 20913
rect 17682 20839 17684 20848
rect 17736 20839 17738 20848
rect 17684 20810 17736 20816
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17788 20380 17816 23734
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17880 21962 17908 22374
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 18064 21010 18092 26250
rect 18248 24290 18276 26862
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18340 24750 18368 25094
rect 18524 24993 18552 25094
rect 18510 24984 18566 24993
rect 18510 24919 18566 24928
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18328 24744 18380 24750
rect 18432 24721 18460 24754
rect 18328 24686 18380 24692
rect 18418 24712 18474 24721
rect 18418 24647 18474 24656
rect 18248 24274 18368 24290
rect 18236 24268 18368 24274
rect 18288 24262 18368 24268
rect 18236 24210 18288 24216
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18248 23866 18276 24074
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18340 23338 18368 24262
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18432 23730 18460 24074
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18432 23497 18460 23666
rect 18418 23488 18474 23497
rect 18418 23423 18474 23432
rect 18340 23310 18460 23338
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17868 20392 17920 20398
rect 17788 20352 17868 20380
rect 17868 20334 17920 20340
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 20058 17816 20198
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17408 19440 17460 19446
rect 17314 19408 17370 19417
rect 17408 19382 17460 19388
rect 17314 19343 17370 19352
rect 17420 18970 17448 19382
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16854 16008 16910 16017
rect 16854 15943 16910 15952
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16776 11257 16804 15846
rect 16868 15502 16896 15846
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16948 14816 17000 14822
rect 17052 14793 17080 17138
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17328 16182 17356 16390
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 16948 14758 17000 14764
rect 17038 14784 17094 14793
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 13938 16896 14418
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16868 13394 16896 13874
rect 16960 13705 16988 14758
rect 17038 14719 17094 14728
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 16946 13696 17002 13705
rect 16946 13631 17002 13640
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16868 12850 16896 13330
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 17144 12434 17172 14350
rect 17236 13258 17264 14826
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17328 12434 17356 15302
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17420 13705 17448 13942
rect 17406 13696 17462 13705
rect 17406 13631 17462 13640
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17052 12406 17172 12434
rect 17236 12406 17356 12434
rect 16762 11248 16818 11257
rect 16762 11183 16818 11192
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 11121 16988 11154
rect 16946 11112 17002 11121
rect 16946 11047 17002 11056
rect 16856 10056 16908 10062
rect 16670 10024 16726 10033
rect 16856 9998 16908 10004
rect 16670 9959 16726 9968
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16488 9512 16540 9518
rect 16684 9466 16712 9959
rect 16488 9454 16540 9460
rect 16592 9438 16712 9466
rect 16764 9444 16816 9450
rect 16592 9194 16620 9438
rect 16764 9386 16816 9392
rect 16500 9166 16620 9194
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16500 8276 16528 9166
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 8634 16620 8978
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16776 8378 16804 9386
rect 16868 8974 16896 9998
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16946 8936 17002 8945
rect 16868 8634 16896 8910
rect 16946 8871 17002 8880
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16868 8430 16896 8570
rect 16408 8248 16528 8276
rect 16684 8350 16804 8378
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16302 8120 16358 8129
rect 16302 8055 16358 8064
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16316 7886 16344 8055
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16408 7274 16436 8248
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16118 5536 16174 5545
rect 16118 5471 16174 5480
rect 16132 5302 16160 5471
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16224 5114 16252 7142
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16316 5778 16344 6190
rect 16408 5846 16436 7210
rect 16500 6390 16528 7754
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16592 6390 16620 7686
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16578 5808 16634 5817
rect 16304 5772 16356 5778
rect 16578 5743 16634 5752
rect 16304 5714 16356 5720
rect 16592 5710 16620 5743
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16302 5400 16358 5409
rect 16302 5335 16358 5344
rect 16132 5086 16252 5114
rect 16316 5098 16344 5335
rect 16304 5092 16356 5098
rect 16026 3360 16082 3369
rect 16026 3295 16082 3304
rect 16040 2922 16068 3295
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 15252 2468 15424 2496
rect 15200 2450 15252 2456
rect 16132 800 16160 5086
rect 16304 5034 16356 5040
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4826 16252 4966
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16316 4282 16344 5034
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16592 4486 16620 4694
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16304 4072 16356 4078
rect 16302 4040 16304 4049
rect 16356 4040 16358 4049
rect 16302 3975 16358 3984
rect 16592 3670 16620 4422
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16316 3194 16344 3402
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16684 2774 16712 8350
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 7342 16804 8230
rect 16868 7954 16896 8366
rect 16960 8090 16988 8871
rect 17052 8276 17080 12406
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17144 12073 17172 12106
rect 17130 12064 17186 12073
rect 17130 11999 17186 12008
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17144 10810 17172 11222
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17144 9586 17172 10746
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17130 8936 17186 8945
rect 17130 8871 17132 8880
rect 17184 8871 17186 8880
rect 17132 8842 17184 8848
rect 17144 8430 17172 8842
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17052 8248 17172 8276
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16960 7449 16988 7482
rect 16946 7440 17002 7449
rect 16946 7375 17002 7384
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6866 16896 7278
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 7002 16988 7142
rect 16948 6996 17000 7002
rect 17052 6984 17080 7822
rect 17144 7750 17172 8248
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 7206 17172 7686
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17052 6956 17172 6984
rect 16948 6938 17000 6944
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16776 5250 16804 6666
rect 16868 5778 16896 6802
rect 17052 6254 17080 6802
rect 17144 6254 17172 6956
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17236 5778 17264 12406
rect 17420 12238 17448 12650
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 9178 17356 9318
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17406 9072 17462 9081
rect 17512 9042 17540 19790
rect 17880 18442 17908 20334
rect 18156 19786 18184 22374
rect 18340 22234 18368 22578
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18328 22228 18380 22234
rect 18328 22170 18380 22176
rect 18248 20398 18276 22170
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 18050 19544 18106 19553
rect 18050 19479 18106 19488
rect 18064 18766 18092 19479
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17880 18414 18184 18442
rect 18156 18358 18184 18414
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17604 10033 17632 18226
rect 18064 17338 18092 18294
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17696 14006 17724 15642
rect 17788 15570 17816 15642
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17788 15026 17816 15506
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17880 14328 17908 16934
rect 17972 16522 18000 17002
rect 18156 16538 18184 17478
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 18064 16510 18184 16538
rect 17972 16046 18000 16458
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17972 15638 18000 15982
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17960 14340 18012 14346
rect 17880 14300 17960 14328
rect 17960 14282 18012 14288
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 18064 13682 18092 16510
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 16182 18184 16390
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17696 13654 18092 13682
rect 17590 10024 17646 10033
rect 17590 9959 17646 9968
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 9042 17632 9454
rect 17406 9007 17462 9016
rect 17500 9036 17552 9042
rect 17420 7585 17448 9007
rect 17500 8978 17552 8984
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17406 7576 17462 7585
rect 17406 7511 17408 7520
rect 17460 7511 17462 7520
rect 17408 7482 17460 7488
rect 17420 7451 17448 7482
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6934 17540 7142
rect 17604 7041 17632 8978
rect 17590 7032 17646 7041
rect 17590 6967 17646 6976
rect 17500 6928 17552 6934
rect 17406 6896 17462 6905
rect 17500 6870 17552 6876
rect 17406 6831 17462 6840
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 16776 5222 16896 5250
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16776 3534 16804 5102
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 2990 16804 3470
rect 16868 3108 16896 5222
rect 17144 5166 17172 5714
rect 17420 5642 17448 6831
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17144 4690 17172 5102
rect 17236 4826 17264 5578
rect 17604 5001 17632 6190
rect 17696 5817 17724 13654
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17776 13388 17828 13394
rect 17828 13348 17908 13376
rect 17776 13330 17828 13336
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 12918 17816 13126
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17788 7546 17816 12854
rect 17880 12306 17908 13348
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17880 10810 17908 12242
rect 17972 11694 18000 12378
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18064 10470 18092 13466
rect 18156 11354 18184 15302
rect 18248 13802 18276 20198
rect 18328 18216 18380 18222
rect 18326 18184 18328 18193
rect 18380 18184 18382 18193
rect 18326 18119 18382 18128
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 17270 18368 18022
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18432 17134 18460 23310
rect 18524 19310 18552 24006
rect 18616 21554 18644 26318
rect 18708 22094 18736 26862
rect 18800 26586 18828 26998
rect 18788 26580 18840 26586
rect 18788 26522 18840 26528
rect 18786 26480 18842 26489
rect 18786 26415 18842 26424
rect 18800 26314 18828 26415
rect 18788 26308 18840 26314
rect 18788 26250 18840 26256
rect 18984 25945 19012 28018
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 19260 26858 19288 27338
rect 19352 27334 19380 27814
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 18970 25936 19026 25945
rect 18970 25871 19026 25880
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18892 23798 18920 24006
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 18708 22066 18828 22094
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18616 20806 18644 21490
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18616 18970 18644 19382
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18616 18086 18644 18770
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18708 16833 18736 17614
rect 18694 16824 18750 16833
rect 18694 16759 18750 16768
rect 18602 16688 18658 16697
rect 18602 16623 18604 16632
rect 18656 16623 18658 16632
rect 18604 16594 18656 16600
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18432 15337 18460 15438
rect 18418 15328 18474 15337
rect 18418 15263 18474 15272
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18340 12918 18368 15030
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18432 12434 18460 13806
rect 18524 13530 18552 16526
rect 18800 16046 18828 22066
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18892 20534 18920 21286
rect 18880 20528 18932 20534
rect 18880 20470 18932 20476
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18892 19242 18920 19722
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18892 18902 18920 19178
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18984 15722 19012 25871
rect 19076 22438 19104 26794
rect 19260 26518 19288 26794
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 19260 25838 19288 26454
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19248 25832 19300 25838
rect 19154 25800 19210 25809
rect 19248 25774 19300 25780
rect 19154 25735 19210 25744
rect 19168 24818 19196 25735
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19168 22250 19196 24754
rect 19076 22222 19196 22250
rect 19076 20505 19104 22222
rect 19352 22094 19380 26386
rect 19444 22778 19472 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19524 26852 19576 26858
rect 19524 26794 19576 26800
rect 19536 26314 19564 26794
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19708 24676 19760 24682
rect 19708 24618 19760 24624
rect 19614 24576 19670 24585
rect 19614 24511 19670 24520
rect 19628 24138 19656 24511
rect 19720 24206 19748 24618
rect 19890 24440 19946 24449
rect 19890 24375 19946 24384
rect 19904 24342 19932 24375
rect 19892 24336 19944 24342
rect 19892 24278 19944 24284
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19536 23050 19564 23734
rect 19904 23225 19932 23802
rect 19890 23216 19946 23225
rect 19890 23151 19946 23160
rect 19524 23044 19576 23050
rect 19524 22986 19576 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22778 20024 32438
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 20088 26450 20116 28562
rect 20168 26512 20220 26518
rect 20166 26480 20168 26489
rect 20220 26480 20222 26489
rect 20076 26444 20128 26450
rect 20166 26415 20222 26424
rect 20076 26386 20128 26392
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20076 25968 20128 25974
rect 20076 25910 20128 25916
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 19536 22273 19564 22578
rect 20088 22386 20116 25910
rect 19996 22358 20116 22386
rect 19522 22264 19578 22273
rect 19522 22199 19578 22208
rect 19892 22094 19944 22098
rect 19352 22092 19944 22094
rect 19352 22066 19892 22092
rect 19892 22034 19944 22040
rect 19432 22024 19484 22030
rect 19338 21992 19394 22001
rect 19432 21966 19484 21972
rect 19338 21927 19394 21936
rect 19352 21622 19380 21927
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19248 21548 19300 21554
rect 19444 21536 19472 21966
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21690 20024 22358
rect 20074 22128 20130 22137
rect 20074 22063 20130 22072
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19616 21548 19668 21554
rect 19444 21508 19616 21536
rect 19248 21490 19300 21496
rect 19616 21490 19668 21496
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 19062 20496 19118 20505
rect 19062 20431 19118 20440
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 18616 15694 19012 15722
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18432 12406 18552 12434
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18142 11248 18198 11257
rect 18142 11183 18198 11192
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17880 8129 17908 10406
rect 18050 9752 18106 9761
rect 18050 9687 18106 9696
rect 17866 8120 17922 8129
rect 17866 8055 17922 8064
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17972 6118 18000 6666
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17682 5808 17738 5817
rect 17682 5743 17738 5752
rect 18064 5302 18092 9687
rect 18156 5642 18184 11183
rect 18248 9518 18276 11834
rect 18340 10606 18368 12038
rect 18524 11830 18552 12406
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18420 10600 18472 10606
rect 18616 10588 18644 15694
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 15337 18920 15438
rect 18878 15328 18934 15337
rect 18878 15263 18934 15272
rect 18696 15088 18748 15094
rect 18984 15042 19012 15506
rect 19076 15065 19104 18702
rect 18696 15030 18748 15036
rect 18708 14618 18736 15030
rect 18800 15014 19012 15042
rect 19062 15056 19118 15065
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 14074 18736 14214
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18800 14006 18828 15014
rect 19062 14991 19118 15000
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18892 14346 18920 14894
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18708 11558 18736 13738
rect 18786 13288 18842 13297
rect 18786 13223 18842 13232
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11014 18736 11494
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18800 10826 18828 13223
rect 18892 12102 18920 14010
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18472 10560 18644 10588
rect 18708 10798 18828 10826
rect 18420 10542 18472 10548
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 9178 18276 9318
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18248 8265 18276 9114
rect 18234 8256 18290 8265
rect 18234 8191 18290 8200
rect 18340 7750 18368 10406
rect 18432 10130 18460 10542
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 9489 18460 9522
rect 18512 9512 18564 9518
rect 18418 9480 18474 9489
rect 18512 9454 18564 9460
rect 18418 9415 18474 9424
rect 18524 8974 18552 9454
rect 18512 8968 18564 8974
rect 18510 8936 18512 8945
rect 18564 8936 18566 8945
rect 18510 8871 18566 8880
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18234 6216 18290 6225
rect 18234 6151 18290 6160
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 17314 4992 17370 5001
rect 17314 4927 17370 4936
rect 17590 4992 17646 5001
rect 17590 4927 17646 4936
rect 17328 4826 17356 4927
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17236 4570 17264 4626
rect 17052 4554 17264 4570
rect 17040 4548 17264 4554
rect 17092 4542 17264 4548
rect 17406 4584 17462 4593
rect 17406 4519 17408 4528
rect 17040 4490 17092 4496
rect 17460 4519 17462 4528
rect 17408 4490 17460 4496
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17500 3936 17552 3942
rect 17498 3904 17500 3913
rect 17684 3936 17736 3942
rect 17552 3904 17554 3913
rect 17684 3878 17736 3884
rect 17498 3839 17554 3848
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 17040 3120 17092 3126
rect 16868 3080 17040 3108
rect 17040 3062 17092 3068
rect 17236 2990 17264 3402
rect 16764 2984 16816 2990
rect 17132 2984 17184 2990
rect 16816 2932 16896 2938
rect 16764 2926 16896 2932
rect 17132 2926 17184 2932
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 16776 2910 16896 2926
rect 16776 2861 16804 2910
rect 16684 2746 16804 2774
rect 16670 2680 16726 2689
rect 16580 2644 16632 2650
rect 16670 2615 16672 2624
rect 16580 2586 16632 2592
rect 16724 2615 16726 2624
rect 16672 2586 16724 2592
rect 16592 2530 16620 2586
rect 16592 2502 16712 2530
rect 16684 1970 16712 2502
rect 16580 1964 16632 1970
rect 16580 1906 16632 1912
rect 16672 1964 16724 1970
rect 16672 1906 16724 1912
rect 16592 1630 16620 1906
rect 16580 1624 16632 1630
rect 16580 1566 16632 1572
rect 16776 800 16804 2746
rect 16868 2514 16896 2910
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17144 2038 17172 2926
rect 17696 2854 17724 3878
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17788 2854 17816 3130
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17972 2774 18000 4082
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18064 3194 18092 4014
rect 18248 3534 18276 6151
rect 18340 4690 18368 7414
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18432 4078 18460 8366
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18524 7886 18552 7958
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18510 7576 18566 7585
rect 18510 7511 18566 7520
rect 18524 7342 18552 7511
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18340 3670 18368 4014
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17972 2746 18092 2774
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17236 2038 17264 2246
rect 17132 2032 17184 2038
rect 17132 1974 17184 1980
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 17604 1902 17632 2314
rect 17592 1896 17644 1902
rect 17592 1838 17644 1844
rect 18064 800 18092 2746
rect 18248 1834 18276 2790
rect 18236 1828 18288 1834
rect 18236 1770 18288 1776
rect 18524 1766 18552 6598
rect 18616 5930 18644 9687
rect 18708 7478 18736 10798
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18800 6882 18828 10474
rect 18892 10198 18920 10950
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18892 9382 18920 9522
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18984 8566 19012 14894
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 11830 19104 14758
rect 19168 14074 19196 20742
rect 19260 14346 19288 21490
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19446 19380 19654
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19444 18850 19472 21286
rect 19628 20806 19656 21490
rect 19812 21350 19840 21626
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19904 20874 19932 21422
rect 19892 20868 19944 20874
rect 19892 20810 19944 20816
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 20810
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 20088 20482 20116 22063
rect 20180 22001 20208 26250
rect 20272 25294 20300 28630
rect 20364 28626 20392 32438
rect 21192 30938 21220 37198
rect 22480 36922 22508 37198
rect 22572 37126 22600 39200
rect 23216 37262 23244 39200
rect 23848 37324 23900 37330
rect 23848 37266 23900 37272
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 22560 37120 22612 37126
rect 22560 37062 22612 37068
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 21180 30932 21232 30938
rect 21180 30874 21232 30880
rect 21824 30388 21876 30394
rect 21824 30330 21876 30336
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 20640 29102 20668 29242
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20628 29096 20680 29102
rect 20628 29038 20680 29044
rect 20916 28966 20944 29106
rect 21468 28994 21496 29582
rect 21836 29238 21864 30330
rect 21916 30320 21968 30326
rect 21916 30262 21968 30268
rect 21928 29850 21956 30262
rect 22112 30190 22140 31078
rect 22100 30184 22152 30190
rect 22100 30126 22152 30132
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 21824 29232 21876 29238
rect 21824 29174 21876 29180
rect 22112 28994 22140 30126
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 21468 28966 21680 28994
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 21272 28960 21324 28966
rect 21272 28902 21324 28908
rect 20352 28620 20404 28626
rect 20352 28562 20404 28568
rect 21284 28490 21312 28902
rect 21364 28620 21416 28626
rect 21364 28562 21416 28568
rect 21272 28484 21324 28490
rect 21272 28426 21324 28432
rect 21376 28370 21404 28562
rect 21284 28342 21404 28370
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20352 27532 20404 27538
rect 20352 27474 20404 27480
rect 20364 27130 20392 27474
rect 20352 27124 20404 27130
rect 20352 27066 20404 27072
rect 20260 25288 20312 25294
rect 20258 25256 20260 25265
rect 20312 25256 20314 25265
rect 20258 25191 20314 25200
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20272 23118 20300 24346
rect 20364 23474 20392 27066
rect 20456 27062 20484 27814
rect 20444 27056 20496 27062
rect 20444 26998 20496 27004
rect 20640 25480 20668 28018
rect 20720 27668 20772 27674
rect 20720 27610 20772 27616
rect 20732 26926 20760 27610
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20824 26042 20852 27338
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20456 25452 20668 25480
rect 20456 24313 20484 25452
rect 20626 25392 20682 25401
rect 20626 25327 20682 25336
rect 20640 25294 20668 25327
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20442 24304 20498 24313
rect 20548 24274 20576 25162
rect 20720 24744 20772 24750
rect 20640 24692 20720 24698
rect 20640 24686 20772 24692
rect 20640 24670 20760 24686
rect 20442 24239 20498 24248
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20456 23905 20484 24142
rect 20442 23896 20498 23905
rect 20442 23831 20498 23840
rect 20548 23662 20576 24210
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20364 23446 20576 23474
rect 20350 23352 20406 23361
rect 20350 23287 20406 23296
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20272 22137 20300 22170
rect 20258 22128 20314 22137
rect 20258 22063 20314 22072
rect 20166 21992 20222 22001
rect 20166 21927 20222 21936
rect 20258 20904 20314 20913
rect 20258 20839 20314 20848
rect 19996 20454 20116 20482
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19352 18834 19472 18850
rect 19340 18828 19472 18834
rect 19392 18822 19472 18828
rect 19340 18770 19392 18776
rect 19536 18680 19564 18906
rect 19904 18698 19932 18906
rect 19352 18652 19564 18680
rect 19892 18692 19944 18698
rect 19352 17610 19380 18652
rect 19892 18634 19944 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19892 18352 19944 18358
rect 19890 18320 19892 18329
rect 19944 18320 19946 18329
rect 19890 18255 19946 18264
rect 19432 18080 19484 18086
rect 19430 18048 19432 18057
rect 19484 18048 19486 18057
rect 19430 17983 19486 17992
rect 19524 17672 19576 17678
rect 19576 17620 19932 17626
rect 19524 17614 19932 17620
rect 19340 17604 19392 17610
rect 19536 17598 19932 17614
rect 19340 17546 19392 17552
rect 19904 17542 19932 17598
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19352 16182 19380 16526
rect 19904 16522 19932 16730
rect 19892 16516 19944 16522
rect 19892 16458 19944 16464
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19340 16176 19392 16182
rect 19444 16153 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19340 16118 19392 16124
rect 19430 16144 19486 16153
rect 19430 16079 19486 16088
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15502 19656 15846
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 15144 19380 15370
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19352 15116 19564 15144
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19430 14784 19486 14793
rect 19352 14618 19380 14758
rect 19430 14719 19486 14728
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19340 14408 19392 14414
rect 19444 14396 19472 14719
rect 19392 14368 19472 14396
rect 19340 14350 19392 14356
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19536 14278 19564 15116
rect 19996 14278 20024 20454
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20088 19310 20116 20334
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 20180 18329 20208 19926
rect 20166 18320 20222 18329
rect 20076 18284 20128 18290
rect 20166 18255 20222 18264
rect 20076 18226 20128 18232
rect 20088 18170 20116 18226
rect 20088 18142 20208 18170
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20088 17270 20116 18022
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16028 20116 17070
rect 20180 16182 20208 18142
rect 20272 16561 20300 20839
rect 20364 19530 20392 23287
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20456 19666 20484 23054
rect 20548 22094 20576 23446
rect 20640 22710 20668 24670
rect 20720 24132 20772 24138
rect 20720 24074 20772 24080
rect 20732 23798 20760 24074
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20732 23497 20760 23598
rect 20718 23488 20774 23497
rect 20718 23423 20774 23432
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20548 22066 20668 22094
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 20913 20576 21490
rect 20534 20904 20590 20913
rect 20534 20839 20590 20848
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 19802 20576 20742
rect 20640 19990 20668 22066
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20628 19848 20680 19854
rect 20548 19796 20628 19802
rect 20548 19790 20680 19796
rect 20548 19774 20668 19790
rect 20456 19638 20576 19666
rect 20364 19502 20484 19530
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20364 18154 20392 19382
rect 20352 18148 20404 18154
rect 20352 18090 20404 18096
rect 20456 17354 20484 19502
rect 20364 17326 20484 17354
rect 20258 16552 20314 16561
rect 20258 16487 20314 16496
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20168 16176 20220 16182
rect 20272 16153 20300 16390
rect 20168 16118 20220 16124
rect 20258 16144 20314 16153
rect 20258 16079 20314 16088
rect 20088 16000 20208 16028
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20088 15502 20116 15642
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20180 15434 20208 16000
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19340 14000 19392 14006
rect 19338 13968 19340 13977
rect 19392 13968 19394 13977
rect 19338 13903 19394 13912
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19432 13864 19484 13870
rect 19628 13841 19656 13874
rect 19996 13870 20024 14214
rect 19984 13864 20036 13870
rect 19432 13806 19484 13812
rect 19614 13832 19670 13841
rect 19352 13002 19380 13806
rect 19260 12974 19380 13002
rect 19154 12744 19210 12753
rect 19154 12679 19156 12688
rect 19208 12679 19210 12688
rect 19156 12650 19208 12656
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 19260 9874 19288 12974
rect 19338 12744 19394 12753
rect 19444 12730 19472 13806
rect 19984 13806 20036 13812
rect 19614 13767 19670 13776
rect 19628 13326 19656 13767
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19708 12776 19760 12782
rect 19444 12702 19656 12730
rect 19708 12718 19760 12724
rect 19338 12679 19394 12688
rect 19352 12646 19380 12679
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19076 9846 19288 9874
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 19076 8294 19104 9846
rect 19352 9674 19380 12582
rect 19430 12472 19486 12481
rect 19628 12442 19656 12702
rect 19720 12646 19748 12718
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19430 12407 19432 12416
rect 19484 12407 19486 12416
rect 19616 12436 19668 12442
rect 19432 12378 19484 12384
rect 19996 12434 20024 13126
rect 20088 12617 20116 15302
rect 20180 14618 20208 15370
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20272 14396 20300 15846
rect 20364 15745 20392 17326
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20350 15736 20406 15745
rect 20350 15671 20406 15680
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20180 14368 20300 14396
rect 20074 12608 20130 12617
rect 20074 12543 20130 12552
rect 19616 12378 19668 12384
rect 19904 12406 20024 12434
rect 20074 12472 20130 12481
rect 20074 12407 20130 12416
rect 19904 12345 19932 12406
rect 19984 12368 20036 12374
rect 19890 12336 19946 12345
rect 19432 12300 19484 12306
rect 19984 12310 20036 12316
rect 19890 12271 19946 12280
rect 19432 12242 19484 12248
rect 19444 11898 19472 12242
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19444 11218 19472 11834
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 11218 19748 11494
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 9926 19932 10406
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19352 9646 19472 9674
rect 19248 9512 19300 9518
rect 19246 9480 19248 9489
rect 19300 9480 19302 9489
rect 19246 9415 19302 9424
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8974 19380 9318
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 8566 19380 8910
rect 19444 8906 19472 9646
rect 19890 9480 19946 9489
rect 19890 9415 19946 9424
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19628 9178 19656 9318
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19432 8900 19484 8906
rect 19904 8888 19932 9415
rect 19996 9042 20024 12310
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19904 8860 20024 8888
rect 19432 8842 19484 8848
rect 19444 8634 19472 8842
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19154 8392 19210 8401
rect 19154 8327 19210 8336
rect 19168 8294 19196 8327
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19352 7954 19380 8502
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19444 7818 19472 8230
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 18984 7177 19012 7754
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7426 20024 8860
rect 19352 7398 20024 7426
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 18878 7032 18934 7041
rect 18878 6967 18934 6976
rect 18708 6854 18828 6882
rect 18708 6236 18736 6854
rect 18788 6792 18840 6798
rect 18892 6780 18920 6967
rect 18840 6752 18920 6780
rect 19156 6792 19208 6798
rect 18788 6734 18840 6740
rect 19352 6746 19380 7398
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19156 6734 19208 6740
rect 19168 6497 19196 6734
rect 19260 6718 19380 6746
rect 19154 6488 19210 6497
rect 19154 6423 19210 6432
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18892 6254 18920 6326
rect 18788 6248 18840 6254
rect 18708 6208 18788 6236
rect 18788 6190 18840 6196
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18800 6066 18828 6190
rect 18800 6038 19104 6066
rect 18616 5902 19012 5930
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18616 2258 18644 4150
rect 18708 3670 18736 4558
rect 18800 4214 18828 5714
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18892 5370 18920 5578
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18892 4593 18920 4626
rect 18878 4584 18934 4593
rect 18878 4519 18934 4528
rect 18788 4208 18840 4214
rect 18788 4150 18840 4156
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18800 3398 18828 3674
rect 18984 3466 19012 5902
rect 19076 5302 19104 6038
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 19260 4622 19288 6718
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18984 2922 19012 3402
rect 19076 3369 19104 3402
rect 19062 3360 19118 3369
rect 19062 3295 19118 3304
rect 19260 3194 19288 3470
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18972 2916 19024 2922
rect 18972 2858 19024 2864
rect 19260 2854 19288 3130
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 18616 2230 18736 2258
rect 18512 1760 18564 1766
rect 18512 1702 18564 1708
rect 18708 800 18736 2230
rect 18892 1698 18920 2314
rect 18880 1692 18932 1698
rect 18880 1634 18932 1640
rect 19352 800 19380 6598
rect 19444 5030 19472 7210
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19800 6452 19852 6458
rect 19852 6412 20024 6440
rect 19800 6394 19852 6400
rect 19996 5574 20024 6412
rect 20088 6390 20116 12407
rect 20180 7954 20208 14368
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12986 20300 13262
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20364 12617 20392 15302
rect 20350 12608 20406 12617
rect 20350 12543 20406 12552
rect 20456 12481 20484 17138
rect 20548 16969 20576 19638
rect 20534 16960 20590 16969
rect 20534 16895 20590 16904
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20548 16522 20576 16730
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 14822 20576 16050
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 13326 20576 14758
rect 20640 14113 20668 19774
rect 20732 19242 20760 23423
rect 20824 20874 20852 25774
rect 20916 24886 20944 26862
rect 20904 24880 20956 24886
rect 20904 24822 20956 24828
rect 21008 23118 21036 28018
rect 21178 27840 21234 27849
rect 21178 27775 21234 27784
rect 21192 26790 21220 27775
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20916 21457 20944 21490
rect 20902 21448 20958 21457
rect 20902 21383 20958 21392
rect 20916 21350 20944 21383
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 21008 21185 21036 23054
rect 20994 21176 21050 21185
rect 20994 21111 21050 21120
rect 21100 21026 21128 25638
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 21192 24138 21220 25094
rect 21284 24274 21312 28342
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21560 27606 21588 28018
rect 21548 27600 21600 27606
rect 21548 27542 21600 27548
rect 21364 26784 21416 26790
rect 21364 26726 21416 26732
rect 21376 26314 21404 26726
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21468 25226 21496 25638
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 21284 22574 21312 24210
rect 21652 23118 21680 28966
rect 21928 28966 22140 28994
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21836 27606 21864 28358
rect 21824 27600 21876 27606
rect 21824 27542 21876 27548
rect 21836 27402 21864 27542
rect 21824 27396 21876 27402
rect 21824 27338 21876 27344
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 21192 22166 21220 22442
rect 21180 22160 21232 22166
rect 21180 22102 21232 22108
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21284 21622 21312 21898
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 20916 20998 21128 21026
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20916 20466 20944 20998
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20916 20369 20944 20402
rect 20902 20360 20958 20369
rect 20902 20295 20958 20304
rect 20994 19952 21050 19961
rect 20994 19887 21050 19896
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20916 19446 20944 19654
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 18193 20760 18566
rect 20718 18184 20774 18193
rect 20718 18119 20774 18128
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20732 17610 20760 18022
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20824 17610 20852 17818
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20732 17066 20760 17546
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20824 17082 20852 17206
rect 20720 17060 20772 17066
rect 20824 17054 20944 17082
rect 20720 17002 20772 17008
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20824 16794 20852 16934
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20732 15434 20760 15574
rect 20824 15502 20852 16730
rect 20916 16454 20944 17054
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20902 15736 20958 15745
rect 20902 15671 20958 15680
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20824 15026 20852 15438
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20626 14104 20682 14113
rect 20626 14039 20682 14048
rect 20720 14000 20772 14006
rect 20718 13968 20720 13977
rect 20772 13968 20774 13977
rect 20718 13903 20774 13912
rect 20824 13841 20852 14962
rect 20810 13832 20866 13841
rect 20810 13767 20866 13776
rect 20718 13560 20774 13569
rect 20718 13495 20720 13504
rect 20772 13495 20774 13504
rect 20720 13466 20772 13472
rect 20916 13394 20944 15671
rect 21008 13784 21036 19887
rect 21100 19446 21128 20810
rect 21088 19440 21140 19446
rect 21088 19382 21140 19388
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 21100 17882 21128 18294
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21086 15736 21142 15745
rect 21086 15671 21142 15680
rect 21100 15473 21128 15671
rect 21086 15464 21142 15473
rect 21086 15399 21142 15408
rect 21192 13802 21220 21490
rect 21284 17134 21312 21558
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21180 13796 21232 13802
rect 21008 13756 21128 13784
rect 20994 13696 21050 13705
rect 20994 13631 21050 13640
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20902 13288 20958 13297
rect 20902 13223 20958 13232
rect 20536 13184 20588 13190
rect 20534 13152 20536 13161
rect 20812 13184 20864 13190
rect 20588 13152 20590 13161
rect 20534 13087 20590 13096
rect 20718 13152 20774 13161
rect 20812 13126 20864 13132
rect 20718 13087 20774 13096
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20548 12753 20576 12786
rect 20534 12744 20590 12753
rect 20534 12679 20590 12688
rect 20442 12472 20498 12481
rect 20442 12407 20498 12416
rect 20258 12200 20314 12209
rect 20534 12200 20590 12209
rect 20258 12135 20314 12144
rect 20444 12164 20496 12170
rect 20272 11830 20300 12135
rect 20534 12135 20590 12144
rect 20444 12106 20496 12112
rect 20456 11898 20484 12106
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20272 11218 20300 11766
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20442 10976 20498 10985
rect 20442 10911 20498 10920
rect 20350 10704 20406 10713
rect 20350 10639 20406 10648
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20166 7440 20222 7449
rect 20166 7375 20168 7384
rect 20220 7375 20222 7384
rect 20168 7346 20220 7352
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19996 4622 20024 5510
rect 20180 5114 20208 7142
rect 20272 6497 20300 9862
rect 20364 9586 20392 10639
rect 20456 10062 20484 10911
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20442 9888 20498 9897
rect 20442 9823 20498 9832
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20364 7002 20392 7346
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20456 6905 20484 9823
rect 20548 7041 20576 12135
rect 20626 11656 20682 11665
rect 20626 11591 20682 11600
rect 20640 7274 20668 11591
rect 20732 11082 20760 13087
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20824 10742 20852 13126
rect 20812 10736 20864 10742
rect 20718 10704 20774 10713
rect 20812 10678 20864 10684
rect 20718 10639 20774 10648
rect 20732 7478 20760 10639
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9586 20852 9998
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20824 9042 20852 9522
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20824 7546 20852 8026
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20534 7032 20590 7041
rect 20534 6967 20590 6976
rect 20628 6928 20680 6934
rect 20442 6896 20498 6905
rect 20628 6870 20680 6876
rect 20442 6831 20498 6840
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20258 6488 20314 6497
rect 20456 6458 20484 6666
rect 20258 6423 20314 6432
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20364 5710 20392 6258
rect 20640 6254 20668 6870
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20548 5914 20576 6190
rect 20732 6118 20760 6734
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20732 5778 20760 6054
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20352 5704 20404 5710
rect 20824 5658 20852 7142
rect 20352 5646 20404 5652
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20732 5630 20852 5658
rect 20088 5086 20208 5114
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19430 4448 19486 4457
rect 19430 4383 19486 4392
rect 19444 3738 19472 4383
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20088 3126 20116 5086
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 20180 2514 20208 4490
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3602 20300 3878
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20456 2774 20484 5578
rect 20732 3466 20760 5630
rect 20916 5522 20944 13223
rect 21008 11257 21036 13631
rect 21100 12918 21128 13756
rect 21180 13738 21232 13744
rect 21284 13530 21312 14554
rect 21376 14074 21404 22578
rect 21546 21040 21602 21049
rect 21546 20975 21602 20984
rect 21560 20942 21588 20975
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21652 20806 21680 23054
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21560 20602 21588 20742
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19786 21496 20198
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21454 17912 21510 17921
rect 21454 17847 21456 17856
rect 21508 17847 21510 17856
rect 21456 17818 21508 17824
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 16522 21496 17478
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 21100 11540 21128 12854
rect 21192 12782 21220 13262
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21192 12442 21220 12718
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21376 11778 21404 14010
rect 21284 11750 21404 11778
rect 21284 11694 21312 11750
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21100 11512 21312 11540
rect 20994 11248 21050 11257
rect 20994 11183 21050 11192
rect 21008 10010 21036 11183
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21100 10130 21128 10746
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21008 9982 21128 10010
rect 20996 9648 21048 9654
rect 20994 9616 20996 9625
rect 21048 9616 21050 9625
rect 20994 9551 21050 9560
rect 21100 8430 21128 9982
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 8430 21220 8774
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21100 8294 21128 8366
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21178 8120 21234 8129
rect 20996 8084 21048 8090
rect 21178 8055 21234 8064
rect 20996 8026 21048 8032
rect 21008 7342 21036 8026
rect 21192 7954 21220 8055
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21192 7857 21220 7890
rect 21178 7848 21234 7857
rect 21178 7783 21234 7792
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 21086 7304 21142 7313
rect 21086 7239 21142 7248
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21008 5642 21036 6598
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 20824 5494 20944 5522
rect 20824 4146 20852 5494
rect 21100 5370 21128 7239
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 21192 5250 21220 7783
rect 21284 7750 21312 11512
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21100 5222 21220 5250
rect 21284 5234 21312 7686
rect 21376 6662 21404 11630
rect 21468 10713 21496 14894
rect 21560 14074 21588 17614
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21560 12345 21588 12650
rect 21652 12481 21680 18702
rect 21744 17542 21772 23598
rect 21836 21554 21864 25842
rect 21928 23798 21956 28966
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 22020 28082 22048 28698
rect 22756 28558 22784 29582
rect 22836 29028 22888 29034
rect 22836 28970 22888 28976
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22374 27976 22430 27985
rect 22374 27911 22430 27920
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22204 27713 22232 27814
rect 22190 27704 22246 27713
rect 22190 27639 22246 27648
rect 22008 27396 22060 27402
rect 22008 27338 22060 27344
rect 22020 26042 22048 27338
rect 22388 26994 22416 27911
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 22020 25226 22048 25978
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 22020 23594 22048 25162
rect 22376 23792 22428 23798
rect 22204 23752 22376 23780
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21836 19378 21864 20946
rect 21928 20874 21956 22918
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21928 19922 21956 20810
rect 22020 20777 22048 21490
rect 22006 20768 22062 20777
rect 22006 20703 22062 20712
rect 22112 19990 22140 22442
rect 22204 21690 22232 23752
rect 22376 23734 22428 23740
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22376 23044 22428 23050
rect 22376 22986 22428 22992
rect 22388 22574 22416 22986
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21729 22324 21830
rect 22282 21720 22338 21729
rect 22192 21684 22244 21690
rect 22282 21655 22338 21664
rect 22192 21626 22244 21632
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22204 20534 22232 21286
rect 22296 20874 22324 21286
rect 22284 20868 22336 20874
rect 22284 20810 22336 20816
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22284 20528 22336 20534
rect 22284 20470 22336 20476
rect 22296 20330 22324 20470
rect 22388 20398 22416 22510
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 22374 19816 22430 19825
rect 22374 19751 22376 19760
rect 22428 19751 22430 19760
rect 22376 19722 22428 19728
rect 22100 19440 22152 19446
rect 22098 19408 22100 19417
rect 22152 19408 22154 19417
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 22008 19372 22060 19378
rect 22098 19343 22154 19352
rect 22008 19314 22060 19320
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21744 16726 21772 17206
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21836 15994 21864 19314
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21928 17610 21956 18566
rect 21916 17604 21968 17610
rect 21916 17546 21968 17552
rect 22020 16182 22048 19314
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 16522 22232 18022
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 21836 15966 21956 15994
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21744 14414 21772 14962
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21638 12472 21694 12481
rect 21638 12407 21694 12416
rect 21546 12336 21602 12345
rect 21546 12271 21602 12280
rect 21454 10704 21510 10713
rect 21454 10639 21510 10648
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21468 6361 21496 9454
rect 21744 8566 21772 14214
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21836 7750 21864 15846
rect 21928 12646 21956 15966
rect 22204 14482 22232 16050
rect 22296 15570 22324 18702
rect 22480 16182 22508 23258
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22572 21457 22600 22510
rect 22756 22094 22784 28494
rect 22848 27062 22876 28970
rect 22940 28218 22968 37062
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 23032 29646 23060 36654
rect 23584 36378 23612 36722
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23480 36304 23532 36310
rect 23480 36246 23532 36252
rect 23492 35630 23520 36246
rect 23480 35624 23532 35630
rect 23480 35566 23532 35572
rect 23492 30258 23520 35566
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23112 30184 23164 30190
rect 23112 30126 23164 30132
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 23124 28506 23152 30126
rect 23204 29708 23256 29714
rect 23204 29650 23256 29656
rect 23032 28478 23152 28506
rect 22928 28212 22980 28218
rect 22928 28154 22980 28160
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22928 26308 22980 26314
rect 22928 26250 22980 26256
rect 22848 24750 22876 26250
rect 22940 25770 22968 26250
rect 22928 25764 22980 25770
rect 22928 25706 22980 25712
rect 23032 25650 23060 28478
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 23124 25974 23152 28358
rect 23112 25968 23164 25974
rect 23112 25910 23164 25916
rect 23112 25764 23164 25770
rect 23112 25706 23164 25712
rect 22940 25622 23060 25650
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22664 22066 22784 22094
rect 22558 21448 22614 21457
rect 22558 21383 22614 21392
rect 22572 20534 22600 21383
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22572 19718 22600 20334
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 16182 22600 17478
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22572 14890 22600 15574
rect 22560 14884 22612 14890
rect 22560 14826 22612 14832
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21928 10470 21956 12582
rect 22020 11218 22048 13738
rect 22112 13410 22140 13806
rect 22112 13394 22232 13410
rect 22112 13388 22244 13394
rect 22112 13382 22192 13388
rect 22192 13330 22244 13336
rect 22204 13138 22232 13330
rect 22112 13110 22232 13138
rect 22112 11762 22140 13110
rect 22296 12434 22324 14010
rect 22388 13530 22416 14486
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22388 12617 22416 12718
rect 22374 12608 22430 12617
rect 22374 12543 22430 12552
rect 22296 12406 22416 12434
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22112 11218 22140 11698
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 22388 9654 22416 12406
rect 22480 12170 22508 14282
rect 22572 12594 22600 14554
rect 22664 13394 22692 22066
rect 22744 22024 22796 22030
rect 22742 21992 22744 22001
rect 22796 21992 22798 22001
rect 22742 21927 22798 21936
rect 22756 21690 22784 21927
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22848 21185 22876 24686
rect 22940 23186 22968 25622
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 23032 24138 23060 24686
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 23124 23508 23152 25706
rect 23216 23769 23244 29650
rect 23584 29646 23612 36314
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23388 29504 23440 29510
rect 23388 29446 23440 29452
rect 23296 28416 23348 28422
rect 23296 28358 23348 28364
rect 23308 28150 23336 28358
rect 23296 28144 23348 28150
rect 23296 28086 23348 28092
rect 23400 28014 23428 29446
rect 23480 29232 23532 29238
rect 23480 29174 23532 29180
rect 23492 28966 23520 29174
rect 23676 29102 23704 29990
rect 23768 29238 23796 29990
rect 23756 29232 23808 29238
rect 23756 29174 23808 29180
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23388 28008 23440 28014
rect 23388 27950 23440 27956
rect 23400 25838 23428 27950
rect 23676 27674 23704 29038
rect 23768 28218 23796 29038
rect 23756 28212 23808 28218
rect 23756 28154 23808 28160
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23492 26897 23520 27406
rect 23478 26888 23534 26897
rect 23478 26823 23534 26832
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23202 23760 23258 23769
rect 23202 23695 23258 23704
rect 23204 23656 23256 23662
rect 23202 23624 23204 23633
rect 23256 23624 23258 23633
rect 23202 23559 23258 23568
rect 23124 23480 23244 23508
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22834 21176 22890 21185
rect 22834 21111 22890 21120
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22848 19378 22876 20266
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22940 18680 22968 21830
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19786 23060 20198
rect 23020 19780 23072 19786
rect 23020 19722 23072 19728
rect 23018 19680 23074 19689
rect 23018 19615 23074 19624
rect 23032 19446 23060 19615
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23216 18834 23244 23480
rect 23308 23322 23336 23802
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23294 21176 23350 21185
rect 23294 21111 23350 21120
rect 23308 20874 23336 21111
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 23400 19378 23428 25774
rect 23572 25220 23624 25226
rect 23572 25162 23624 25168
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 22710 23520 24550
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23492 20913 23520 22102
rect 23584 22098 23612 25162
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23676 23118 23704 23462
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23768 22386 23796 27950
rect 23860 24682 23888 37266
rect 24032 37256 24084 37262
rect 24032 37198 24084 37204
rect 24504 37210 24532 39200
rect 24044 36922 24072 37198
rect 24400 37188 24452 37194
rect 24504 37182 24624 37210
rect 24400 37130 24452 37136
rect 24032 36916 24084 36922
rect 24032 36858 24084 36864
rect 24216 36780 24268 36786
rect 24216 36722 24268 36728
rect 24228 35834 24256 36722
rect 24216 35828 24268 35834
rect 24216 35770 24268 35776
rect 24412 30734 24440 37130
rect 24596 37126 24624 37182
rect 25148 37126 25176 39200
rect 25792 37262 25820 39200
rect 26516 37324 26568 37330
rect 26516 37266 26568 37272
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 26056 37188 26108 37194
rect 26056 37130 26108 37136
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 26068 32910 26096 37130
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 25228 32768 25280 32774
rect 25228 32710 25280 32716
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24858 30152 24914 30161
rect 24858 30087 24914 30096
rect 24872 30054 24900 30087
rect 24860 30048 24912 30054
rect 24860 29990 24912 29996
rect 25240 29714 25268 32710
rect 25596 30660 25648 30666
rect 25596 30602 25648 30608
rect 25504 30184 25556 30190
rect 25504 30126 25556 30132
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25516 29578 25544 30126
rect 25320 29572 25372 29578
rect 25320 29514 25372 29520
rect 25504 29572 25556 29578
rect 25504 29514 25556 29520
rect 24032 29504 24084 29510
rect 24032 29446 24084 29452
rect 23940 29232 23992 29238
rect 23940 29174 23992 29180
rect 23952 27470 23980 29174
rect 24044 28490 24072 29446
rect 25332 29306 25360 29514
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 24216 28552 24268 28558
rect 24216 28494 24268 28500
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 24032 28484 24084 28490
rect 24032 28426 24084 28432
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 24122 27432 24178 27441
rect 24122 27367 24178 27376
rect 24136 26314 24164 27367
rect 24228 26353 24256 28494
rect 25044 28484 25096 28490
rect 25044 28426 25096 28432
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24584 28008 24636 28014
rect 24584 27950 24636 27956
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24214 26344 24270 26353
rect 24124 26308 24176 26314
rect 24214 26279 24270 26288
rect 24124 26250 24176 26256
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23848 24676 23900 24682
rect 23848 24618 23900 24624
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23860 23633 23888 24074
rect 23846 23624 23902 23633
rect 23846 23559 23902 23568
rect 23952 23322 23980 24754
rect 24044 23338 24072 25774
rect 24228 25294 24256 26279
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 24216 24880 24268 24886
rect 24216 24822 24268 24828
rect 24228 24410 24256 24822
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 24124 24336 24176 24342
rect 24124 24278 24176 24284
rect 24136 24138 24164 24278
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 24320 23798 24348 24618
rect 24308 23792 24360 23798
rect 24214 23760 24270 23769
rect 24308 23734 24360 23740
rect 24214 23695 24216 23704
rect 24268 23695 24270 23704
rect 24216 23666 24268 23672
rect 23940 23316 23992 23322
rect 24044 23310 24256 23338
rect 23940 23258 23992 23264
rect 24032 23248 24084 23254
rect 24032 23190 24084 23196
rect 23676 22358 23796 22386
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23572 21616 23624 21622
rect 23570 21584 23572 21593
rect 23624 21584 23626 21593
rect 23570 21519 23626 21528
rect 23478 20904 23534 20913
rect 23478 20839 23534 20848
rect 23676 20058 23704 22358
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23768 21486 23796 22170
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23768 20534 23796 21422
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23768 19922 23796 20470
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19446 23704 19654
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23020 18692 23072 18698
rect 22940 18652 23020 18680
rect 23020 18634 23072 18640
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 22742 16960 22798 16969
rect 22742 16895 22798 16904
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22572 12566 22692 12594
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22572 11801 22600 12378
rect 22664 12238 22692 12566
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22558 11792 22614 11801
rect 22558 11727 22614 11736
rect 22572 10538 22600 11727
rect 22652 11212 22704 11218
rect 22756 11200 22784 16895
rect 22704 11172 22784 11200
rect 22652 11154 22704 11160
rect 22560 10532 22612 10538
rect 22560 10474 22612 10480
rect 22756 10130 22784 11172
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22848 9654 22876 18566
rect 23676 18426 23704 18566
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23020 18080 23072 18086
rect 23018 18048 23020 18057
rect 23072 18048 23074 18057
rect 23018 17983 23074 17992
rect 23020 16516 23072 16522
rect 23020 16458 23072 16464
rect 23032 15638 23060 16458
rect 23112 15972 23164 15978
rect 23112 15914 23164 15920
rect 23124 15881 23152 15914
rect 23110 15872 23166 15881
rect 23110 15807 23166 15816
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22940 13462 22968 14894
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22020 8838 22048 9522
rect 22284 9376 22336 9382
rect 22112 9336 22284 9364
rect 22112 9178 22140 9336
rect 22284 9318 22336 9324
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22100 9036 22152 9042
rect 22204 9024 22232 9114
rect 22152 8996 22232 9024
rect 22100 8978 22152 8984
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21560 7002 21588 7278
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21454 6352 21510 6361
rect 21454 6287 21510 6296
rect 21272 5228 21324 5234
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20916 4010 20944 4558
rect 21008 4282 21036 5102
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20548 3108 20576 3402
rect 20548 3080 20852 3108
rect 20824 2990 20852 3080
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20456 2746 20668 2774
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20640 800 20668 2746
rect 20732 2310 20760 2858
rect 20916 2854 20944 3946
rect 21100 2922 21128 5222
rect 21272 5170 21324 5176
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21192 4826 21220 4966
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21284 4554 21312 4762
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21468 4185 21496 4422
rect 21454 4176 21510 4185
rect 21454 4111 21510 4120
rect 21270 3224 21326 3233
rect 21270 3159 21326 3168
rect 21284 3126 21312 3159
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20916 2514 20944 2790
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 21376 1970 21404 2314
rect 21364 1964 21416 1970
rect 21364 1906 21416 1912
rect 21284 870 21404 898
rect 21284 800 21312 870
rect 1858 776 1914 785
rect 1858 711 1914 720
rect 2594 200 2650 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 5170 200 5226 800
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12254 200 12310 800
rect 13542 200 13598 800
rect 14186 200 14242 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 18694 200 18750 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21270 200 21326 800
rect 21376 762 21404 870
rect 21560 762 21588 4422
rect 21652 3058 21680 6938
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21744 5846 21772 6122
rect 21822 6080 21878 6089
rect 21822 6015 21878 6024
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21836 4214 21864 6015
rect 21824 4208 21876 4214
rect 21824 4150 21876 4156
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21730 3768 21786 3777
rect 21730 3703 21786 3712
rect 21744 3602 21772 3703
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21836 3398 21864 4014
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21822 3224 21878 3233
rect 21928 3194 21956 8434
rect 22020 7954 22048 8774
rect 22282 8256 22338 8265
rect 22282 8191 22338 8200
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 22020 7410 22048 7890
rect 22192 7812 22244 7818
rect 22192 7754 22244 7760
rect 22204 7721 22232 7754
rect 22190 7712 22246 7721
rect 22190 7647 22246 7656
rect 22296 7478 22324 8191
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22296 6458 22324 6938
rect 22388 6662 22416 9590
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22834 9480 22890 9489
rect 22664 8294 22692 9454
rect 22834 9415 22890 9424
rect 22848 9042 22876 9415
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22848 8430 22876 8978
rect 22836 8424 22888 8430
rect 22742 8392 22798 8401
rect 22836 8366 22888 8372
rect 22742 8327 22798 8336
rect 22480 8266 22692 8294
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22008 6248 22060 6254
rect 22376 6248 22428 6254
rect 22008 6190 22060 6196
rect 22112 6196 22376 6202
rect 22112 6190 22428 6196
rect 22020 5778 22048 6190
rect 22112 6174 22416 6190
rect 22112 6118 22140 6174
rect 22100 6112 22152 6118
rect 22284 6112 22336 6118
rect 22100 6054 22152 6060
rect 22282 6080 22284 6089
rect 22336 6080 22338 6089
rect 22282 6015 22338 6024
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22020 5166 22048 5714
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 21822 3159 21824 3168
rect 21876 3159 21878 3168
rect 21916 3188 21968 3194
rect 21824 3130 21876 3136
rect 21916 3130 21968 3136
rect 22020 3058 22048 5102
rect 22204 4826 22232 5578
rect 22282 5536 22338 5545
rect 22282 5471 22338 5480
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 22204 3126 22232 4150
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22296 2990 22324 5471
rect 22374 4992 22430 5001
rect 22374 4927 22430 4936
rect 22388 4078 22416 4927
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22480 3670 22508 8266
rect 22756 8242 22784 8327
rect 22756 8214 22876 8242
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22572 7478 22600 7686
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22848 7002 22876 8214
rect 22836 6996 22888 7002
rect 22836 6938 22888 6944
rect 22742 6896 22798 6905
rect 22742 6831 22798 6840
rect 22756 6798 22784 6831
rect 22848 6798 22876 6938
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22650 5944 22706 5953
rect 22650 5879 22652 5888
rect 22704 5879 22706 5888
rect 22652 5850 22704 5856
rect 22756 5030 22784 6734
rect 22940 6458 22968 13398
rect 23032 8974 23060 14418
rect 23124 12374 23152 15642
rect 23216 15314 23244 18158
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23296 17264 23348 17270
rect 23348 17224 23520 17252
rect 23296 17206 23348 17212
rect 23296 17128 23348 17134
rect 23348 17088 23428 17116
rect 23296 17070 23348 17076
rect 23400 16454 23428 17088
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23308 15570 23336 16390
rect 23400 16028 23428 16390
rect 23492 16182 23520 17224
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23480 16040 23532 16046
rect 23400 16000 23480 16028
rect 23480 15982 23532 15988
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23480 15360 23532 15366
rect 23216 15286 23336 15314
rect 23480 15302 23532 15308
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23216 13190 23244 13466
rect 23204 13184 23256 13190
rect 23204 13126 23256 13132
rect 23308 12434 23336 15286
rect 23492 14958 23520 15302
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23216 12406 23336 12434
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23112 12164 23164 12170
rect 23112 12106 23164 12112
rect 23124 11354 23152 12106
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23216 8786 23244 12406
rect 23400 9178 23428 13330
rect 23492 13326 23520 14894
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23032 8758 23244 8786
rect 23032 7954 23060 8758
rect 23110 8664 23166 8673
rect 23110 8599 23166 8608
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23032 6458 23060 7890
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23124 6338 23152 8599
rect 23202 6488 23258 6497
rect 23202 6423 23258 6432
rect 22940 6310 23152 6338
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 22848 5710 22876 5850
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22468 3664 22520 3670
rect 22468 3606 22520 3612
rect 22480 3369 22508 3606
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 22466 3360 22522 3369
rect 22466 3295 22522 3304
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22296 2378 22324 2926
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22296 1902 22324 2314
rect 22284 1896 22336 1902
rect 22284 1838 22336 1844
rect 22572 800 22600 3130
rect 22664 2106 22692 3402
rect 22940 3126 22968 6310
rect 23216 4622 23244 6423
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 23032 3670 23060 3878
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 23124 3398 23152 3878
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 23216 800 23244 3334
rect 23308 2378 23336 8978
rect 23584 7546 23612 17614
rect 23676 15502 23704 18226
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23386 7440 23442 7449
rect 23386 7375 23442 7384
rect 23400 5234 23428 7375
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23492 6118 23520 6598
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 23492 2990 23520 4014
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23584 2514 23612 7482
rect 23676 6730 23704 15302
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23768 14550 23796 14962
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23768 14414 23796 14486
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23860 14362 23888 21966
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23952 21146 23980 21558
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23940 20936 23992 20942
rect 23938 20904 23940 20913
rect 23992 20904 23994 20913
rect 23938 20839 23994 20848
rect 24044 20788 24072 23190
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24136 21078 24164 21422
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 23952 20760 24072 20788
rect 23952 19446 23980 20760
rect 24032 19984 24084 19990
rect 24032 19926 24084 19932
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17270 23980 17478
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 24044 17134 24072 19926
rect 24136 19310 24164 21014
rect 24228 20992 24256 23310
rect 24412 22094 24440 27270
rect 24596 26926 24624 27950
rect 24780 27402 24808 28358
rect 24872 28150 24900 28358
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 24676 27396 24728 27402
rect 24676 27338 24728 27344
rect 24768 27396 24820 27402
rect 24768 27338 24820 27344
rect 24688 27282 24716 27338
rect 24688 27254 24808 27282
rect 24780 27062 24808 27254
rect 24676 27056 24728 27062
rect 24676 26998 24728 27004
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24492 26852 24544 26858
rect 24492 26794 24544 26800
rect 24504 26314 24532 26794
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24504 24750 24532 26250
rect 24596 25974 24624 26862
rect 24688 26586 24716 26998
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24676 26580 24728 26586
rect 24676 26522 24728 26528
rect 24780 26314 24808 26726
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24584 25968 24636 25974
rect 24584 25910 24636 25916
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24596 24993 24624 25162
rect 24582 24984 24638 24993
rect 24582 24919 24638 24928
rect 24492 24744 24544 24750
rect 24492 24686 24544 24692
rect 24780 24410 24808 25230
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24872 24342 24900 26862
rect 24952 26512 25004 26518
rect 24950 26480 24952 26489
rect 25004 26480 25006 26489
rect 24950 26415 25006 26424
rect 24964 25838 24992 26415
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 24952 25696 25004 25702
rect 24952 25638 25004 25644
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 24964 24018 24992 25638
rect 24872 23990 24992 24018
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24504 22778 24532 23054
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24412 22066 24532 22094
rect 24308 21004 24360 21010
rect 24228 20964 24308 20992
rect 24308 20946 24360 20952
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24228 20398 24256 20538
rect 24320 20398 24348 20946
rect 24400 20528 24452 20534
rect 24400 20470 24452 20476
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24228 18970 24256 19722
rect 24412 19334 24440 20470
rect 24320 19306 24440 19334
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24122 16280 24178 16289
rect 24122 16215 24124 16224
rect 24176 16215 24178 16224
rect 24124 16186 24176 16192
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 24044 15609 24072 16050
rect 24030 15600 24086 15609
rect 24030 15535 24086 15544
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 23860 14334 23980 14362
rect 23952 14074 23980 14334
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23768 11830 23796 14010
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23952 12918 23980 13126
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 23938 12472 23994 12481
rect 23938 12407 23994 12416
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23676 2378 23704 6190
rect 23768 4690 23796 11222
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23860 8498 23888 8774
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23952 5574 23980 12407
rect 24044 9110 24072 15302
rect 24214 14920 24270 14929
rect 24320 14890 24348 19306
rect 24504 19174 24532 22066
rect 24780 21146 24808 22986
rect 24872 21418 24900 23990
rect 24950 23896 25006 23905
rect 24950 23831 25006 23840
rect 24964 23662 24992 23831
rect 24952 23656 25004 23662
rect 24952 23598 25004 23604
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24964 22710 24992 23462
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 25056 22574 25084 28426
rect 25148 25945 25176 28494
rect 25134 25936 25190 25945
rect 25134 25871 25190 25880
rect 25148 22710 25176 25871
rect 25240 23730 25268 29106
rect 25504 27940 25556 27946
rect 25504 27882 25556 27888
rect 25410 27840 25466 27849
rect 25410 27775 25466 27784
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25332 26518 25360 27338
rect 25320 26512 25372 26518
rect 25320 26454 25372 26460
rect 25332 25702 25360 26454
rect 25320 25696 25372 25702
rect 25320 25638 25372 25644
rect 25424 24818 25452 27775
rect 25516 25838 25544 27882
rect 25504 25832 25556 25838
rect 25504 25774 25556 25780
rect 25504 25220 25556 25226
rect 25504 25162 25556 25168
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 25410 24712 25466 24721
rect 25410 24647 25466 24656
rect 25318 24440 25374 24449
rect 25318 24375 25374 24384
rect 25332 24206 25360 24375
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25424 24070 25452 24647
rect 25516 24410 25544 25162
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 25412 24064 25464 24070
rect 25412 24006 25464 24012
rect 25516 23882 25544 24210
rect 25332 23854 25544 23882
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 24964 20942 24992 21082
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 24964 20777 24992 20878
rect 24950 20768 25006 20777
rect 24950 20703 25006 20712
rect 25056 19922 25084 22510
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25148 21962 25176 22374
rect 25240 21962 25268 23462
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25148 21486 25176 21898
rect 25332 21842 25360 23854
rect 25608 23746 25636 30602
rect 26148 28960 26200 28966
rect 26148 28902 26200 28908
rect 26332 28960 26384 28966
rect 26332 28902 26384 28908
rect 26160 28626 26188 28902
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26344 28490 26372 28902
rect 26332 28484 26384 28490
rect 26332 28426 26384 28432
rect 25780 28144 25832 28150
rect 25780 28086 25832 28092
rect 25792 27849 25820 28086
rect 26528 28082 26556 37266
rect 27080 37126 27108 39200
rect 27724 37262 27752 39200
rect 29012 37262 29040 39200
rect 27528 37256 27580 37262
rect 27528 37198 27580 37204
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 26700 30320 26752 30326
rect 26700 30262 26752 30268
rect 26792 30320 26844 30326
rect 26792 30262 26844 30268
rect 26712 29646 26740 30262
rect 26804 29850 26832 30262
rect 26884 30048 26936 30054
rect 26884 29990 26936 29996
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26700 29640 26752 29646
rect 26700 29582 26752 29588
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 26516 28076 26568 28082
rect 26516 28018 26568 28024
rect 25870 27976 25926 27985
rect 25870 27911 25926 27920
rect 25778 27840 25834 27849
rect 25778 27775 25834 27784
rect 25780 27532 25832 27538
rect 25780 27474 25832 27480
rect 25792 26450 25820 27474
rect 25780 26444 25832 26450
rect 25780 26386 25832 26392
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25700 25430 25728 25842
rect 25792 25702 25820 26386
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 25688 25424 25740 25430
rect 25688 25366 25740 25372
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25700 24342 25728 24754
rect 25688 24336 25740 24342
rect 25688 24278 25740 24284
rect 25516 23718 25636 23746
rect 25688 23724 25740 23730
rect 25516 23322 25544 23718
rect 25688 23666 25740 23672
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25240 21814 25360 21842
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 21010 25176 21422
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25240 20534 25268 21814
rect 25424 20602 25452 22918
rect 25516 22642 25544 23258
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25516 21622 25544 21898
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 25516 20602 25544 20742
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25228 20528 25280 20534
rect 25228 20470 25280 20476
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24504 18766 24532 19110
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24504 16726 24532 17682
rect 24676 17604 24728 17610
rect 24780 17592 24808 18158
rect 24728 17564 24808 17592
rect 24676 17546 24728 17552
rect 24780 16998 24808 17564
rect 24858 17232 24914 17241
rect 24858 17167 24914 17176
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24492 16720 24544 16726
rect 24492 16662 24544 16668
rect 24872 16658 24900 17167
rect 25148 16946 25176 19994
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 25332 18442 25360 19926
rect 25608 18986 25636 23598
rect 25700 21049 25728 23666
rect 25792 23254 25820 25638
rect 25780 23248 25832 23254
rect 25780 23190 25832 23196
rect 25778 21584 25834 21593
rect 25778 21519 25834 21528
rect 25686 21040 25742 21049
rect 25686 20975 25742 20984
rect 25700 20806 25728 20975
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25792 20466 25820 21519
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25884 20233 25912 27911
rect 26252 27674 26280 28018
rect 26424 27872 26476 27878
rect 26424 27814 26476 27820
rect 26240 27668 26292 27674
rect 26240 27610 26292 27616
rect 26436 27402 26464 27814
rect 26700 27532 26752 27538
rect 26700 27474 26752 27480
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26148 26512 26200 26518
rect 26200 26460 26372 26466
rect 26148 26454 26372 26460
rect 26160 26450 26372 26454
rect 26160 26444 26384 26450
rect 26160 26438 26332 26444
rect 26332 26386 26384 26392
rect 26148 25968 26200 25974
rect 26148 25910 26200 25916
rect 26160 24834 26188 25910
rect 26160 24818 26372 24834
rect 26160 24812 26384 24818
rect 26160 24806 26332 24812
rect 26332 24754 26384 24760
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 25976 22098 26004 24686
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 26238 24576 26294 24585
rect 26068 23050 26096 24550
rect 26238 24511 26294 24520
rect 26252 23186 26280 24511
rect 26436 24342 26464 26930
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 26528 24410 26556 25094
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26620 24342 26648 27066
rect 26712 26450 26740 27474
rect 26896 27062 26924 29990
rect 27252 29028 27304 29034
rect 27252 28970 27304 28976
rect 26976 28484 27028 28490
rect 26976 28426 27028 28432
rect 26884 27056 26936 27062
rect 26884 26998 26936 27004
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 26700 26444 26752 26450
rect 26700 26386 26752 26392
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26712 24954 26740 25162
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26700 24744 26752 24750
rect 26700 24686 26752 24692
rect 26424 24336 26476 24342
rect 26608 24336 26660 24342
rect 26476 24284 26556 24290
rect 26424 24278 26556 24284
rect 26608 24278 26660 24284
rect 26436 24262 26556 24278
rect 26424 24200 26476 24206
rect 26424 24142 26476 24148
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 25964 21480 26016 21486
rect 25962 21448 25964 21457
rect 26016 21448 26018 21457
rect 25962 21383 26018 21392
rect 25870 20224 25926 20233
rect 25870 20159 25926 20168
rect 25884 20058 25912 20159
rect 25872 20052 25924 20058
rect 25872 19994 25924 20000
rect 25608 18958 25912 18986
rect 25686 18728 25742 18737
rect 25686 18663 25742 18672
rect 25780 18692 25832 18698
rect 25700 18630 25728 18663
rect 25780 18634 25832 18640
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25332 18414 25452 18442
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25056 16918 25176 16946
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24412 15162 24440 15438
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24214 14855 24270 14864
rect 24308 14884 24360 14890
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24136 10266 24164 14758
rect 24228 12782 24256 14855
rect 24308 14826 24360 14832
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24320 11558 24348 14826
rect 24412 12850 24440 15098
rect 24504 14414 24532 15370
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24492 13456 24544 13462
rect 24492 13398 24544 13404
rect 24504 13190 24532 13398
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24596 12434 24624 16526
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24688 15337 24716 16050
rect 24860 15904 24912 15910
rect 24860 15846 24912 15852
rect 24872 15609 24900 15846
rect 24858 15600 24914 15609
rect 24858 15535 24860 15544
rect 24912 15535 24914 15544
rect 24860 15506 24912 15512
rect 24674 15328 24730 15337
rect 24674 15263 24730 15272
rect 24964 14958 24992 16050
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 13938 24900 14418
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24768 13388 24820 13394
rect 24872 13376 24900 13874
rect 24820 13348 24900 13376
rect 24768 13330 24820 13336
rect 24964 13258 24992 14758
rect 25056 13258 25084 16918
rect 25332 16590 25360 18294
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25148 15502 25176 15642
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25148 15026 25176 15438
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25148 13734 25176 14554
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24596 12406 24716 12434
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 24412 10810 24440 10950
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24122 8528 24178 8537
rect 24122 8463 24178 8472
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24044 7002 24072 7278
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 24136 6882 24164 8463
rect 24412 7886 24440 8978
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24044 6854 24164 6882
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 23952 5098 23980 5510
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23860 2514 23888 2994
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 23296 2372 23348 2378
rect 23296 2314 23348 2320
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 23768 2106 23796 2246
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 23768 1630 23796 2042
rect 23952 1714 23980 3402
rect 24044 2854 24072 6854
rect 24228 6254 24256 7278
rect 24308 6656 24360 6662
rect 24306 6624 24308 6633
rect 24360 6624 24362 6633
rect 24306 6559 24362 6568
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24228 5778 24256 6190
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 24320 4690 24348 5102
rect 24412 5001 24440 7822
rect 24504 6390 24532 12242
rect 24582 12200 24638 12209
rect 24582 12135 24638 12144
rect 24596 11150 24624 12135
rect 24688 11150 24716 12406
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24582 10568 24638 10577
rect 24582 10503 24638 10512
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 24596 5930 24624 10503
rect 24688 9518 24716 11086
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24780 9654 24808 11018
rect 24964 10742 24992 12582
rect 24952 10736 25004 10742
rect 24952 10678 25004 10684
rect 25056 10606 25084 13194
rect 25148 11354 25176 13670
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24766 9480 24822 9489
rect 24766 9415 24822 9424
rect 24780 9382 24808 9415
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24674 9072 24730 9081
rect 24674 9007 24730 9016
rect 24504 5902 24624 5930
rect 24504 5302 24532 5902
rect 24582 5808 24638 5817
rect 24582 5743 24638 5752
rect 24492 5296 24544 5302
rect 24492 5238 24544 5244
rect 24398 4992 24454 5001
rect 24398 4927 24454 4936
rect 24308 4684 24360 4690
rect 24308 4626 24360 4632
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24228 4282 24256 4422
rect 24320 4282 24348 4626
rect 24504 4554 24532 5238
rect 24596 4758 24624 5743
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24492 4548 24544 4554
rect 24492 4490 24544 4496
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24228 3913 24256 4014
rect 24214 3904 24270 3913
rect 24214 3839 24270 3848
rect 24216 3052 24268 3058
rect 24320 3040 24348 4218
rect 24504 3777 24532 4218
rect 24582 4040 24638 4049
rect 24582 3975 24638 3984
rect 24490 3768 24546 3777
rect 24490 3703 24546 3712
rect 24504 3126 24532 3703
rect 24596 3534 24624 3975
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24492 3120 24544 3126
rect 24492 3062 24544 3068
rect 24268 3012 24348 3040
rect 24216 2994 24268 3000
rect 24124 2916 24176 2922
rect 24124 2858 24176 2864
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 24136 2378 24164 2858
rect 24688 2774 24716 9007
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24872 8650 24900 8842
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24780 8634 24900 8650
rect 24768 8628 24900 8634
rect 24820 8622 24900 8628
rect 24768 8570 24820 8576
rect 24872 8090 24900 8622
rect 24964 8430 24992 8774
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24780 7041 24808 8026
rect 24766 7032 24822 7041
rect 24766 6967 24822 6976
rect 24872 6882 24900 8026
rect 24780 6854 24900 6882
rect 24780 5710 24808 6854
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 4622 24808 5646
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24780 3670 24808 4558
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24688 2746 24808 2774
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24780 2106 24808 2746
rect 24872 2378 24900 4014
rect 24964 3126 24992 8230
rect 25056 4196 25084 10202
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 25148 8430 25176 9454
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25240 7478 25268 15846
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25332 12434 25360 15642
rect 25424 15638 25452 18414
rect 25792 17814 25820 18634
rect 25688 17808 25740 17814
rect 25688 17750 25740 17756
rect 25780 17808 25832 17814
rect 25780 17750 25832 17756
rect 25700 17610 25728 17750
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 25502 17368 25558 17377
rect 25502 17303 25558 17312
rect 25516 17270 25544 17303
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25516 16794 25544 17070
rect 25608 16794 25636 17546
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25700 16697 25728 17546
rect 25686 16688 25742 16697
rect 25686 16623 25742 16632
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25516 15910 25544 16390
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25412 15632 25464 15638
rect 25412 15574 25464 15580
rect 25504 13728 25556 13734
rect 25504 13670 25556 13676
rect 25332 12406 25452 12434
rect 25318 12336 25374 12345
rect 25318 12271 25374 12280
rect 25228 7472 25280 7478
rect 25228 7414 25280 7420
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6254 25176 6598
rect 25240 6458 25268 6734
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25228 5160 25280 5166
rect 25332 5148 25360 12271
rect 25280 5120 25360 5148
rect 25228 5102 25280 5108
rect 25136 4208 25188 4214
rect 25056 4168 25136 4196
rect 25136 4150 25188 4156
rect 25240 3233 25268 5102
rect 25424 4690 25452 12406
rect 25516 12306 25544 13670
rect 25596 12640 25648 12646
rect 25596 12582 25648 12588
rect 25608 12374 25636 12582
rect 25596 12368 25648 12374
rect 25596 12310 25648 12316
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25516 11762 25544 12106
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25700 11370 25728 16458
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25608 11342 25728 11370
rect 25502 11112 25558 11121
rect 25502 11047 25558 11056
rect 25516 8362 25544 11047
rect 25608 8838 25636 11342
rect 25792 11200 25820 15302
rect 25700 11172 25820 11200
rect 25700 9994 25728 11172
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 25884 9466 25912 18958
rect 25964 18964 26016 18970
rect 25964 18906 26016 18912
rect 25976 18426 26004 18906
rect 25964 18420 26016 18426
rect 25964 18362 26016 18368
rect 26068 17746 26096 22034
rect 26160 21146 26188 23054
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26252 21010 26280 22918
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26344 21962 26372 22374
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26160 19854 26188 19994
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 26160 19145 26188 19790
rect 26252 19446 26280 20198
rect 26240 19440 26292 19446
rect 26240 19382 26292 19388
rect 26344 19258 26372 20742
rect 26252 19230 26372 19258
rect 26146 19136 26202 19145
rect 26146 19071 26202 19080
rect 26056 17740 26108 17746
rect 26056 17682 26108 17688
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 15638 26188 15982
rect 26148 15632 26200 15638
rect 26148 15574 26200 15580
rect 26160 15094 26188 15574
rect 26252 15178 26280 19230
rect 26330 18864 26386 18873
rect 26330 18799 26386 18808
rect 26344 18358 26372 18799
rect 26332 18352 26384 18358
rect 26332 18294 26384 18300
rect 26436 18057 26464 24142
rect 26422 18048 26478 18057
rect 26422 17983 26478 17992
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 26436 16998 26464 17070
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26436 16794 26464 16934
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26528 16232 26556 24262
rect 26620 17814 26648 24278
rect 26712 23050 26740 24686
rect 26700 23044 26752 23050
rect 26700 22986 26752 22992
rect 26712 22953 26740 22986
rect 26698 22944 26754 22953
rect 26698 22879 26754 22888
rect 26804 19281 26832 26726
rect 26896 23662 26924 26998
rect 26988 24857 27016 28426
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27172 27985 27200 28018
rect 27158 27976 27214 27985
rect 27158 27911 27214 27920
rect 27264 27538 27292 28970
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27158 26888 27214 26897
rect 27158 26823 27160 26832
rect 27212 26823 27214 26832
rect 27160 26794 27212 26800
rect 27264 26518 27292 27474
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27356 27062 27384 27406
rect 27344 27056 27396 27062
rect 27344 26998 27396 27004
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 27356 26518 27384 26862
rect 27252 26512 27304 26518
rect 27252 26454 27304 26460
rect 27344 26512 27396 26518
rect 27344 26454 27396 26460
rect 27068 26444 27120 26450
rect 27068 26386 27120 26392
rect 27080 25514 27108 26386
rect 27160 26240 27212 26246
rect 27160 26182 27212 26188
rect 27172 25906 27200 26182
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27080 25486 27200 25514
rect 26974 24848 27030 24857
rect 26974 24783 27030 24792
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26882 23216 26938 23225
rect 26988 23202 27016 24783
rect 26938 23174 27016 23202
rect 26882 23151 26938 23160
rect 26896 21962 26924 23151
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 27080 21690 27108 23054
rect 27068 21684 27120 21690
rect 27068 21626 27120 21632
rect 27066 20496 27122 20505
rect 26884 20460 26936 20466
rect 27066 20431 27068 20440
rect 26884 20402 26936 20408
rect 27120 20431 27122 20440
rect 27068 20402 27120 20408
rect 26790 19272 26846 19281
rect 26790 19207 26846 19216
rect 26790 19136 26846 19145
rect 26790 19071 26846 19080
rect 26698 18728 26754 18737
rect 26698 18663 26700 18672
rect 26752 18663 26754 18672
rect 26700 18634 26752 18640
rect 26698 18048 26754 18057
rect 26698 17983 26754 17992
rect 26608 17808 26660 17814
rect 26608 17750 26660 17756
rect 26436 16204 26556 16232
rect 26332 15700 26384 15706
rect 26332 15642 26384 15648
rect 26344 15366 26372 15642
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26252 15150 26372 15178
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 25962 12336 26018 12345
rect 25962 12271 26018 12280
rect 25976 12170 26004 12271
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 26068 11830 26096 14758
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 25964 10736 26016 10742
rect 25964 10678 26016 10684
rect 25700 9438 25912 9466
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25594 6896 25650 6905
rect 25594 6831 25650 6840
rect 25608 6322 25636 6831
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 25700 4570 25728 9438
rect 25976 9364 26004 10678
rect 26054 10568 26110 10577
rect 26054 10503 26056 10512
rect 26108 10503 26110 10512
rect 26056 10474 26108 10480
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 26068 9761 26096 9930
rect 26054 9752 26110 9761
rect 26054 9687 26110 9696
rect 26160 9518 26188 14894
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26252 13802 26280 14418
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26252 11218 26280 13738
rect 26344 13462 26372 15150
rect 26332 13456 26384 13462
rect 26332 13398 26384 13404
rect 26436 12442 26464 16204
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26528 15026 26556 15438
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26516 13252 26568 13258
rect 26516 13194 26568 13200
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26344 11014 26372 12038
rect 26424 11620 26476 11626
rect 26424 11562 26476 11568
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26344 10130 26372 10406
rect 26332 10124 26384 10130
rect 26332 10066 26384 10072
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 26344 9382 26372 10066
rect 25884 9336 26004 9364
rect 26332 9376 26384 9382
rect 25780 8356 25832 8362
rect 25780 8298 25832 8304
rect 25792 5030 25820 8298
rect 25884 8294 25912 9336
rect 26332 9318 26384 9324
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 25608 4542 25728 4570
rect 25608 4078 25636 4542
rect 25688 4480 25740 4486
rect 25688 4422 25740 4428
rect 25780 4480 25832 4486
rect 25780 4422 25832 4428
rect 25700 4214 25728 4422
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25596 4072 25648 4078
rect 25596 4014 25648 4020
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 25226 3224 25282 3233
rect 25226 3159 25282 3168
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 23860 1686 23980 1714
rect 23756 1624 23808 1630
rect 23756 1566 23808 1572
rect 23860 800 23888 1686
rect 25148 870 25268 898
rect 25148 800 25176 870
rect 21376 734 21588 762
rect 22558 200 22614 800
rect 23202 200 23258 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 25240 762 25268 870
rect 25516 762 25544 3946
rect 25608 3602 25636 4014
rect 25792 3602 25820 4422
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 25884 3482 25912 7142
rect 25976 4826 26004 7822
rect 26068 5302 26096 9114
rect 26344 9042 26372 9318
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26436 8514 26464 11562
rect 26252 8486 26464 8514
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 8022 26188 8230
rect 26148 8016 26200 8022
rect 26148 7958 26200 7964
rect 26146 7848 26202 7857
rect 26252 7818 26280 8486
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 26146 7783 26148 7792
rect 26200 7783 26202 7792
rect 26240 7812 26292 7818
rect 26148 7754 26200 7760
rect 26240 7754 26292 7760
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26160 6322 26188 6802
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 26160 5574 26188 6122
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 25792 3454 25912 3482
rect 25792 800 25820 3454
rect 25976 2990 26004 4762
rect 26160 3466 26188 5306
rect 26252 4010 26280 7346
rect 26344 7154 26372 8298
rect 26528 7818 26556 13194
rect 26620 11393 26648 15438
rect 26712 13870 26740 17983
rect 26804 14618 26832 19071
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26896 13546 26924 20402
rect 27172 20346 27200 25486
rect 27264 25362 27292 26454
rect 27448 26314 27476 26930
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 27540 26042 27568 37198
rect 28908 37188 28960 37194
rect 28908 37130 28960 37136
rect 28920 36854 28948 37130
rect 29656 37126 29684 39200
rect 29736 37256 29788 37262
rect 30300 37244 30328 39200
rect 31588 37330 31616 39200
rect 31576 37324 31628 37330
rect 31576 37266 31628 37272
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 29736 37198 29788 37204
rect 30380 37198 30432 37204
rect 30748 37256 30800 37262
rect 30748 37198 30800 37204
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 28908 36848 28960 36854
rect 28908 36790 28960 36796
rect 27988 29232 28040 29238
rect 27988 29174 28040 29180
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27724 27334 27752 28018
rect 27896 27872 27948 27878
rect 27896 27814 27948 27820
rect 27908 27402 27936 27814
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27712 27328 27764 27334
rect 27712 27270 27764 27276
rect 27724 26382 27752 27270
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27252 25356 27304 25362
rect 27252 25298 27304 25304
rect 27620 25356 27672 25362
rect 27620 25298 27672 25304
rect 27434 24984 27490 24993
rect 27434 24919 27490 24928
rect 27448 24886 27476 24919
rect 27436 24880 27488 24886
rect 27436 24822 27488 24828
rect 27632 24614 27660 25298
rect 27804 25220 27856 25226
rect 27804 25162 27856 25168
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27436 24064 27488 24070
rect 27436 24006 27488 24012
rect 27448 23526 27476 24006
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27436 23520 27488 23526
rect 27540 23497 27568 23598
rect 27436 23462 27488 23468
rect 27526 23488 27582 23497
rect 27526 23423 27582 23432
rect 27816 23322 27844 25162
rect 27896 24948 27948 24954
rect 27896 24890 27948 24896
rect 27804 23316 27856 23322
rect 27804 23258 27856 23264
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27344 22976 27396 22982
rect 27724 22953 27752 23054
rect 27344 22918 27396 22924
rect 27710 22944 27766 22953
rect 27356 22710 27384 22918
rect 27710 22879 27766 22888
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27436 22568 27488 22574
rect 27436 22510 27488 22516
rect 27264 22166 27292 22510
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27264 22001 27292 22102
rect 27250 21992 27306 22001
rect 27250 21927 27306 21936
rect 27448 21350 27476 22510
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27436 21344 27488 21350
rect 27434 21312 27436 21321
rect 27488 21312 27490 21321
rect 27434 21247 27490 21256
rect 27540 21078 27568 21898
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27620 21548 27672 21554
rect 27620 21490 27672 21496
rect 27632 21146 27660 21490
rect 27710 21312 27766 21321
rect 27710 21247 27766 21256
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27528 21072 27580 21078
rect 27528 21014 27580 21020
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 27080 20318 27200 20346
rect 27080 19553 27108 20318
rect 27356 19689 27384 20470
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 27448 19922 27476 20266
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 27342 19680 27398 19689
rect 27342 19615 27398 19624
rect 27066 19544 27122 19553
rect 27066 19479 27122 19488
rect 27080 19378 27108 19479
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 27356 19310 27384 19382
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 26988 13802 27016 19110
rect 26976 13796 27028 13802
rect 26976 13738 27028 13744
rect 26896 13518 27016 13546
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26606 11384 26662 11393
rect 26606 11319 26662 11328
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26804 10742 26832 10950
rect 26792 10736 26844 10742
rect 26792 10678 26844 10684
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 26790 9888 26846 9897
rect 26516 7812 26568 7818
rect 26516 7754 26568 7760
rect 26712 7721 26740 9862
rect 26790 9823 26846 9832
rect 26698 7712 26754 7721
rect 26698 7647 26754 7656
rect 26698 7576 26754 7585
rect 26698 7511 26754 7520
rect 26712 7342 26740 7511
rect 26700 7336 26752 7342
rect 26700 7278 26752 7284
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 26620 7177 26648 7210
rect 26606 7168 26662 7177
rect 26344 7126 26464 7154
rect 26330 7032 26386 7041
rect 26330 6967 26332 6976
rect 26384 6967 26386 6976
rect 26332 6938 26384 6944
rect 26332 5636 26384 5642
rect 26332 5578 26384 5584
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26344 3126 26372 5578
rect 26436 5302 26464 7126
rect 26606 7103 26662 7112
rect 26804 6905 26832 9823
rect 26896 9042 26924 13398
rect 26988 13258 27016 13518
rect 26976 13252 27028 13258
rect 26976 13194 27028 13200
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26988 11898 27016 12378
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 26988 10198 27016 11834
rect 27080 11626 27108 19110
rect 27264 18902 27292 19246
rect 27448 19122 27476 19858
rect 27356 19094 27476 19122
rect 27252 18896 27304 18902
rect 27252 18838 27304 18844
rect 27356 18698 27384 19094
rect 27632 18986 27660 20334
rect 27448 18958 27660 18986
rect 27448 18902 27476 18958
rect 27436 18896 27488 18902
rect 27436 18838 27488 18844
rect 27528 18896 27580 18902
rect 27528 18838 27580 18844
rect 27344 18692 27396 18698
rect 27344 18634 27396 18640
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27264 17921 27292 18294
rect 27250 17912 27306 17921
rect 27250 17847 27306 17856
rect 27356 17814 27384 18634
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 27172 16454 27200 17682
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 16046 27292 16390
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27356 15162 27384 17070
rect 27448 15706 27476 18634
rect 27540 18086 27568 18838
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27632 17338 27660 18634
rect 27724 17746 27752 21247
rect 27712 17740 27764 17746
rect 27712 17682 27764 17688
rect 27620 17332 27672 17338
rect 27620 17274 27672 17280
rect 27816 17202 27844 21626
rect 27908 20398 27936 24890
rect 28000 24750 28028 29174
rect 28920 29170 28948 36790
rect 29012 32434 29040 37062
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 29104 30190 29132 30534
rect 29092 30184 29144 30190
rect 29092 30126 29144 30132
rect 28908 29164 28960 29170
rect 28908 29106 28960 29112
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28644 28150 28672 28358
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 28632 28144 28684 28150
rect 28632 28086 28684 28092
rect 29012 28014 29040 28154
rect 29104 28150 29132 30126
rect 29748 29510 29776 37198
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 30288 36848 30340 36854
rect 30288 36790 30340 36796
rect 30300 31754 30328 36790
rect 30208 31726 30328 31754
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 29092 28144 29144 28150
rect 29092 28086 29144 28092
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 29000 28008 29052 28014
rect 29000 27950 29052 27956
rect 28092 27334 28120 27950
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 28184 27441 28212 27474
rect 28170 27432 28226 27441
rect 28170 27367 28226 27376
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 28092 26926 28120 27270
rect 28080 26920 28132 26926
rect 28080 26862 28132 26868
rect 28092 25158 28120 26862
rect 28540 26376 28592 26382
rect 28538 26344 28540 26353
rect 28592 26344 28594 26353
rect 28538 26279 28594 26288
rect 28908 25968 28960 25974
rect 28908 25910 28960 25916
rect 28540 25900 28592 25906
rect 28540 25842 28592 25848
rect 28448 25696 28500 25702
rect 28448 25638 28500 25644
rect 28460 25158 28488 25638
rect 28552 25362 28580 25842
rect 28920 25702 28948 25910
rect 28816 25696 28868 25702
rect 28816 25638 28868 25644
rect 28908 25696 28960 25702
rect 28908 25638 28960 25644
rect 28540 25356 28592 25362
rect 28540 25298 28592 25304
rect 28828 25226 28856 25638
rect 28816 25220 28868 25226
rect 28816 25162 28868 25168
rect 28080 25152 28132 25158
rect 28080 25094 28132 25100
rect 28448 25152 28500 25158
rect 28448 25094 28500 25100
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 27988 24336 28040 24342
rect 27988 24278 28040 24284
rect 28000 24138 28028 24278
rect 28448 24268 28500 24274
rect 28448 24210 28500 24216
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 28460 23866 28488 24210
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28828 23662 28856 25162
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28172 23656 28224 23662
rect 28172 23598 28224 23604
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 28000 21010 28028 21830
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 28080 20868 28132 20874
rect 28080 20810 28132 20816
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27986 19952 28042 19961
rect 27986 19887 28042 19896
rect 28000 19854 28028 19887
rect 27988 19848 28040 19854
rect 27894 19816 27950 19825
rect 27988 19790 28040 19796
rect 27894 19751 27896 19760
rect 27948 19751 27950 19760
rect 27896 19722 27948 19728
rect 28092 19514 28120 20810
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27986 19000 28042 19009
rect 27986 18935 28042 18944
rect 28080 18964 28132 18970
rect 28000 18698 28028 18935
rect 28080 18906 28132 18912
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27908 18086 27936 18566
rect 27986 18456 28042 18465
rect 27986 18391 28042 18400
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27816 16658 27844 17138
rect 28000 17134 28028 18391
rect 28092 18222 28120 18906
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 27804 16652 27856 16658
rect 27724 16612 27804 16640
rect 27724 16250 27752 16612
rect 27804 16594 27856 16600
rect 27804 16516 27856 16522
rect 27804 16458 27856 16464
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27526 15736 27582 15745
rect 27436 15700 27488 15706
rect 27526 15671 27582 15680
rect 27436 15642 27488 15648
rect 27540 15552 27568 15671
rect 27620 15564 27672 15570
rect 27540 15524 27620 15552
rect 27620 15506 27672 15512
rect 27436 15496 27488 15502
rect 27724 15450 27752 16186
rect 27488 15444 27752 15450
rect 27436 15438 27752 15444
rect 27448 15422 27752 15438
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27252 15088 27304 15094
rect 27252 15030 27304 15036
rect 27264 14634 27292 15030
rect 27172 14606 27292 14634
rect 27172 14414 27200 14606
rect 27356 14550 27384 15098
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27436 14884 27488 14890
rect 27436 14826 27488 14832
rect 27344 14544 27396 14550
rect 27344 14486 27396 14492
rect 27252 14476 27304 14482
rect 27252 14418 27304 14424
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27160 13864 27212 13870
rect 27160 13806 27212 13812
rect 27172 13394 27200 13806
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27172 11694 27200 12242
rect 27160 11688 27212 11694
rect 27160 11630 27212 11636
rect 27068 11620 27120 11626
rect 27068 11562 27120 11568
rect 27172 10606 27200 11630
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 26976 10192 27028 10198
rect 26976 10134 27028 10140
rect 27172 10062 27200 10542
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 27172 9586 27200 9998
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26988 9382 27016 9522
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26884 8832 26936 8838
rect 26882 8800 26884 8809
rect 27068 8832 27120 8838
rect 26936 8800 26938 8809
rect 27068 8774 27120 8780
rect 26882 8735 26938 8744
rect 27080 8566 27108 8774
rect 27068 8560 27120 8566
rect 27068 8502 27120 8508
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 27066 8120 27122 8129
rect 27066 8055 27122 8064
rect 26976 7948 27028 7954
rect 26976 7890 27028 7896
rect 26988 7410 27016 7890
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 26790 6896 26846 6905
rect 26988 6866 27016 7346
rect 27080 7018 27108 8055
rect 27172 7954 27200 8366
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 27160 7540 27212 7546
rect 27264 7528 27292 14418
rect 27342 14376 27398 14385
rect 27342 14311 27344 14320
rect 27396 14311 27398 14320
rect 27344 14282 27396 14288
rect 27344 12640 27396 12646
rect 27344 12582 27396 12588
rect 27356 12306 27384 12582
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27344 11824 27396 11830
rect 27344 11766 27396 11772
rect 27356 8974 27384 11766
rect 27448 9994 27476 14826
rect 27540 14396 27568 14962
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27620 14408 27672 14414
rect 27540 14368 27620 14396
rect 27620 14350 27672 14356
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27434 9752 27490 9761
rect 27434 9687 27490 9696
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 27344 8560 27396 8566
rect 27342 8528 27344 8537
rect 27396 8528 27398 8537
rect 27342 8463 27398 8472
rect 27448 7721 27476 9687
rect 27540 8129 27568 13806
rect 27632 12209 27660 14214
rect 27724 14074 27752 14758
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27712 13456 27764 13462
rect 27712 13398 27764 13404
rect 27618 12200 27674 12209
rect 27618 12135 27674 12144
rect 27724 11830 27752 13398
rect 27712 11824 27764 11830
rect 27712 11766 27764 11772
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 27526 8120 27582 8129
rect 27526 8055 27582 8064
rect 27632 7886 27660 10134
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27724 9058 27752 9590
rect 27816 9178 27844 16458
rect 27896 16176 27948 16182
rect 27948 16124 28120 16130
rect 27896 16118 28120 16124
rect 27908 16102 28120 16118
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27908 15094 27936 15914
rect 27988 15904 28040 15910
rect 27988 15846 28040 15852
rect 27896 15088 27948 15094
rect 27896 15030 27948 15036
rect 28000 14090 28028 15846
rect 28092 15706 28120 16102
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 28080 15428 28132 15434
rect 28080 15370 28132 15376
rect 28092 15201 28120 15370
rect 28184 15314 28212 23598
rect 28920 23322 28948 23734
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28264 21480 28316 21486
rect 28262 21448 28264 21457
rect 28316 21448 28318 21457
rect 28262 21383 28318 21392
rect 28264 21004 28316 21010
rect 28264 20946 28316 20952
rect 28276 19990 28304 20946
rect 28368 20058 28396 23054
rect 28540 22976 28592 22982
rect 28540 22918 28592 22924
rect 28552 22710 28580 22918
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 28460 21962 28488 22034
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28908 21956 28960 21962
rect 28908 21898 28960 21904
rect 28814 21720 28870 21729
rect 28814 21655 28870 21664
rect 28632 21480 28684 21486
rect 28552 21440 28632 21468
rect 28552 21185 28580 21440
rect 28632 21422 28684 21428
rect 28722 21448 28778 21457
rect 28828 21434 28856 21655
rect 28920 21622 28948 21898
rect 28908 21616 28960 21622
rect 28908 21558 28960 21564
rect 29012 21434 29040 24686
rect 29196 24682 29224 28426
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29368 26784 29420 26790
rect 29368 26726 29420 26732
rect 29184 24676 29236 24682
rect 29184 24618 29236 24624
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 29104 23662 29132 24550
rect 29092 23656 29144 23662
rect 29092 23598 29144 23604
rect 29380 23118 29408 26726
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 29368 23112 29420 23118
rect 29368 23054 29420 23060
rect 28828 21406 29040 21434
rect 28722 21383 28778 21392
rect 28632 21344 28684 21350
rect 28630 21312 28632 21321
rect 28684 21312 28686 21321
rect 28630 21247 28686 21256
rect 28538 21176 28594 21185
rect 28538 21111 28594 21120
rect 28632 20868 28684 20874
rect 28632 20810 28684 20816
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28276 18193 28304 18702
rect 28262 18184 28318 18193
rect 28262 18119 28318 18128
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28276 17746 28304 18022
rect 28264 17740 28316 17746
rect 28264 17682 28316 17688
rect 28262 17640 28318 17649
rect 28262 17575 28318 17584
rect 28276 17270 28304 17575
rect 28264 17264 28316 17270
rect 28264 17206 28316 17212
rect 28264 16516 28316 16522
rect 28368 16504 28396 19246
rect 28460 18601 28488 19314
rect 28552 19174 28580 19314
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 28644 18737 28672 20810
rect 28736 19922 28764 21383
rect 29012 20482 29040 21406
rect 28920 20454 29040 20482
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28724 19916 28776 19922
rect 28724 19858 28776 19864
rect 28828 19718 28856 20334
rect 28816 19712 28868 19718
rect 28816 19654 28868 19660
rect 28724 19168 28776 19174
rect 28724 19110 28776 19116
rect 28736 19009 28764 19110
rect 28722 19000 28778 19009
rect 28722 18935 28778 18944
rect 28630 18728 28686 18737
rect 28540 18692 28592 18698
rect 28630 18663 28686 18672
rect 28540 18634 28592 18640
rect 28446 18592 28502 18601
rect 28446 18527 28502 18536
rect 28552 18290 28580 18634
rect 28724 18624 28776 18630
rect 28722 18592 28724 18601
rect 28776 18592 28778 18601
rect 28722 18527 28778 18536
rect 28828 18465 28856 19654
rect 28920 19378 28948 20454
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 29012 18902 29040 20334
rect 29000 18896 29052 18902
rect 28906 18864 28962 18873
rect 29000 18838 29052 18844
rect 28906 18799 28962 18808
rect 28814 18456 28870 18465
rect 28632 18420 28684 18426
rect 28920 18426 28948 18799
rect 28814 18391 28870 18400
rect 28908 18420 28960 18426
rect 28632 18362 28684 18368
rect 28908 18362 28960 18368
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28644 18086 28672 18362
rect 28816 18352 28868 18358
rect 28736 18312 28816 18340
rect 28632 18080 28684 18086
rect 28460 18006 28580 18034
rect 28632 18022 28684 18028
rect 28460 17921 28488 18006
rect 28552 17954 28580 18006
rect 28736 17954 28764 18312
rect 28816 18294 28868 18300
rect 28908 18216 28960 18222
rect 28828 18193 28908 18204
rect 28814 18184 28908 18193
rect 28870 18176 28908 18184
rect 28908 18158 28960 18164
rect 28814 18119 28870 18128
rect 28552 17926 28764 17954
rect 28446 17912 28502 17921
rect 28446 17847 28502 17856
rect 28906 17912 28962 17921
rect 28906 17847 28962 17856
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28316 16476 28396 16504
rect 28264 16458 28316 16464
rect 28276 15434 28304 16458
rect 28356 16040 28408 16046
rect 28356 15982 28408 15988
rect 28368 15881 28396 15982
rect 28354 15872 28410 15881
rect 28354 15807 28410 15816
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 28184 15286 28396 15314
rect 28078 15192 28134 15201
rect 28134 15162 28212 15178
rect 28134 15156 28224 15162
rect 28134 15150 28172 15156
rect 28078 15127 28134 15136
rect 28172 15098 28224 15104
rect 28080 15088 28132 15094
rect 28368 15042 28396 15286
rect 28080 15030 28132 15036
rect 27908 14062 28028 14090
rect 27908 13462 27936 14062
rect 27988 14000 28040 14006
rect 27988 13942 28040 13948
rect 27896 13456 27948 13462
rect 27896 13398 27948 13404
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 27908 9994 27936 13194
rect 28000 12986 28028 13942
rect 28092 13326 28120 15030
rect 28184 15014 28396 15042
rect 28460 15042 28488 17614
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28644 16114 28672 16526
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28460 15014 28580 15042
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 28078 11520 28134 11529
rect 28078 11455 28134 11464
rect 27986 11384 28042 11393
rect 27986 11319 28042 11328
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27724 9030 27844 9058
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27724 8809 27752 8842
rect 27710 8800 27766 8809
rect 27710 8735 27766 8744
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27816 7732 27844 9030
rect 27908 8090 27936 9930
rect 28000 8430 28028 11319
rect 28092 10606 28120 11455
rect 28184 11393 28212 15014
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 13954 28396 14894
rect 28448 14816 28500 14822
rect 28448 14758 28500 14764
rect 28460 14074 28488 14758
rect 28448 14068 28500 14074
rect 28448 14010 28500 14016
rect 28368 13926 28488 13954
rect 28460 13870 28488 13926
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28262 13696 28318 13705
rect 28262 13631 28318 13640
rect 28276 12986 28304 13631
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 28368 12434 28396 12815
rect 28552 12434 28580 15014
rect 28276 12406 28396 12434
rect 28460 12406 28580 12434
rect 28630 12472 28686 12481
rect 28630 12407 28632 12416
rect 28170 11384 28226 11393
rect 28170 11319 28226 11328
rect 28170 10840 28226 10849
rect 28170 10775 28226 10784
rect 28080 10600 28132 10606
rect 28080 10542 28132 10548
rect 28184 10418 28212 10775
rect 28092 10390 28212 10418
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 28092 8242 28120 10390
rect 28172 9036 28224 9042
rect 28172 8978 28224 8984
rect 28000 8214 28120 8242
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27908 7886 27936 8026
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27896 7744 27948 7750
rect 27434 7712 27490 7721
rect 27816 7704 27896 7732
rect 27896 7686 27948 7692
rect 27434 7647 27490 7656
rect 27212 7500 27292 7528
rect 27342 7576 27398 7585
rect 27342 7511 27344 7520
rect 27160 7482 27212 7488
rect 27396 7511 27398 7520
rect 27344 7482 27396 7488
rect 27172 7324 27200 7482
rect 27436 7472 27488 7478
rect 27356 7420 27436 7426
rect 27356 7414 27488 7420
rect 27356 7398 27476 7414
rect 27356 7324 27384 7398
rect 27172 7296 27384 7324
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27540 7177 27568 7278
rect 27526 7168 27582 7177
rect 27526 7103 27582 7112
rect 27080 6990 27292 7018
rect 26790 6831 26846 6840
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 27160 6860 27212 6866
rect 27264 6848 27292 6990
rect 27712 6860 27764 6866
rect 27264 6820 27712 6848
rect 27160 6802 27212 6808
rect 27712 6802 27764 6808
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26528 5574 26556 6598
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26424 5296 26476 5302
rect 26424 5238 26476 5244
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 26528 4554 26556 5034
rect 26516 4548 26568 4554
rect 26516 4490 26568 4496
rect 26422 3224 26478 3233
rect 26422 3159 26478 3168
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26436 3058 26464 3159
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26620 2774 26648 6394
rect 27172 6322 27200 6802
rect 27804 6792 27856 6798
rect 27540 6718 27660 6746
rect 27804 6734 27856 6740
rect 27540 6712 27568 6718
rect 27455 6684 27568 6712
rect 27455 6644 27483 6684
rect 27448 6616 27483 6644
rect 27448 6497 27476 6616
rect 27434 6488 27490 6497
rect 27434 6423 27490 6432
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27172 5778 27200 6258
rect 27448 5778 27476 6326
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27540 5953 27568 6190
rect 27526 5944 27582 5953
rect 27526 5879 27582 5888
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 26790 5672 26846 5681
rect 26700 5636 26752 5642
rect 26790 5607 26846 5616
rect 26700 5578 26752 5584
rect 26712 5030 26740 5578
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26804 4729 26832 5607
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 26790 4720 26846 4729
rect 26790 4655 26846 4664
rect 27172 4486 27200 5102
rect 27632 4690 27660 6718
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27160 4480 27212 4486
rect 27160 4422 27212 4428
rect 27172 4078 27200 4422
rect 27528 4208 27580 4214
rect 27528 4150 27580 4156
rect 27160 4072 27212 4078
rect 27540 4049 27568 4150
rect 27160 4014 27212 4020
rect 27526 4040 27582 4049
rect 27068 3120 27120 3126
rect 27068 3062 27120 3068
rect 26974 2952 27030 2961
rect 26974 2887 27030 2896
rect 26988 2854 27016 2887
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 26620 2746 26740 2774
rect 26712 2038 26740 2746
rect 26700 2032 26752 2038
rect 26700 1974 26752 1980
rect 27080 800 27108 3062
rect 27172 2990 27200 4014
rect 27526 3975 27582 3984
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27264 3670 27292 3878
rect 27252 3664 27304 3670
rect 27252 3606 27304 3612
rect 27434 3360 27490 3369
rect 27434 3295 27490 3304
rect 27448 2990 27476 3295
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27436 2984 27488 2990
rect 27436 2926 27488 2932
rect 27172 2854 27200 2926
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 27434 2408 27490 2417
rect 27434 2343 27436 2352
rect 27488 2343 27490 2352
rect 27436 2314 27488 2320
rect 27632 1970 27660 3878
rect 27724 3398 27752 5646
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27816 2774 27844 6734
rect 27894 3904 27950 3913
rect 28000 3890 28028 8214
rect 28080 8016 28132 8022
rect 28080 7958 28132 7964
rect 28092 7546 28120 7958
rect 28080 7540 28132 7546
rect 28080 7482 28132 7488
rect 28078 6488 28134 6497
rect 28078 6423 28134 6432
rect 28092 5642 28120 6423
rect 28080 5636 28132 5642
rect 28080 5578 28132 5584
rect 28184 5302 28212 8978
rect 28276 8537 28304 12406
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28262 8528 28318 8537
rect 28262 8463 28318 8472
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 28276 7546 28304 7754
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28264 6996 28316 7002
rect 28264 6938 28316 6944
rect 28276 6458 28304 6938
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28262 5808 28318 5817
rect 28262 5743 28318 5752
rect 28276 5642 28304 5743
rect 28264 5636 28316 5642
rect 28264 5578 28316 5584
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 28080 4548 28132 4554
rect 28080 4490 28132 4496
rect 27950 3862 28028 3890
rect 27894 3839 27950 3848
rect 27908 3534 27936 3839
rect 28092 3738 28120 4490
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 27988 3460 28040 3466
rect 27988 3402 28040 3408
rect 28000 2990 28028 3402
rect 27988 2984 28040 2990
rect 27988 2926 28040 2932
rect 27724 2746 27844 2774
rect 27620 1964 27672 1970
rect 27620 1906 27672 1912
rect 27724 800 27752 2746
rect 28368 2310 28396 12174
rect 28460 9722 28488 12406
rect 28684 12407 28686 12416
rect 28632 12378 28684 12384
rect 28630 11520 28686 11529
rect 28630 11455 28686 11464
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28644 9602 28672 11455
rect 28736 9738 28764 16594
rect 28816 16516 28868 16522
rect 28816 16458 28868 16464
rect 28828 13258 28856 16458
rect 28920 14618 28948 17847
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 29012 15026 29040 15438
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 28908 14612 28960 14618
rect 28908 14554 28960 14560
rect 28908 13796 28960 13802
rect 28908 13738 28960 13744
rect 28816 13252 28868 13258
rect 28816 13194 28868 13200
rect 28828 12850 28856 13194
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28920 12170 28948 13738
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 29012 10470 29040 14758
rect 29104 13938 29132 23054
rect 29276 22772 29328 22778
rect 29472 22760 29500 26930
rect 29328 22732 29500 22760
rect 29276 22714 29328 22720
rect 29184 20936 29236 20942
rect 29184 20878 29236 20884
rect 29196 18057 29224 20878
rect 29182 18048 29238 18057
rect 29182 17983 29238 17992
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29104 13802 29132 13874
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 29104 11150 29132 12582
rect 29288 12434 29316 22714
rect 29564 22710 29592 27950
rect 29736 27464 29788 27470
rect 29736 27406 29788 27412
rect 29748 27130 29776 27406
rect 29736 27124 29788 27130
rect 29736 27066 29788 27072
rect 29828 26308 29880 26314
rect 29828 26250 29880 26256
rect 29736 25968 29788 25974
rect 29736 25910 29788 25916
rect 29644 22772 29696 22778
rect 29644 22714 29696 22720
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29656 22166 29684 22714
rect 29644 22160 29696 22166
rect 29644 22102 29696 22108
rect 29644 21956 29696 21962
rect 29644 21898 29696 21904
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 29460 20596 29512 20602
rect 29460 20538 29512 20544
rect 29472 20398 29500 20538
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29564 19990 29592 21490
rect 29656 21418 29684 21898
rect 29644 21412 29696 21418
rect 29644 21354 29696 21360
rect 29552 19984 29604 19990
rect 29552 19926 29604 19932
rect 29368 19780 29420 19786
rect 29368 19722 29420 19728
rect 29380 17134 29408 19722
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29472 18193 29500 19314
rect 29656 19310 29684 21354
rect 29748 20602 29776 25910
rect 29840 25226 29868 26250
rect 30208 26058 30236 31726
rect 30484 31346 30512 37062
rect 30760 36718 30788 37198
rect 32232 36922 32260 39200
rect 33520 37126 33548 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 30748 36712 30800 36718
rect 30748 36654 30800 36660
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 30748 32224 30800 32230
rect 30748 32166 30800 32172
rect 30472 31340 30524 31346
rect 30472 31282 30524 31288
rect 30760 29238 30788 32166
rect 31116 30116 31168 30122
rect 31116 30058 31168 30064
rect 30748 29232 30800 29238
rect 30748 29174 30800 29180
rect 31024 29232 31076 29238
rect 31024 29174 31076 29180
rect 31036 28694 31064 29174
rect 31128 29034 31156 30058
rect 31116 29028 31168 29034
rect 31116 28970 31168 28976
rect 31024 28688 31076 28694
rect 31024 28630 31076 28636
rect 30472 28144 30524 28150
rect 30472 28086 30524 28092
rect 30484 27606 30512 28086
rect 30472 27600 30524 27606
rect 30472 27542 30524 27548
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30392 26994 30420 27406
rect 30472 27396 30524 27402
rect 30472 27338 30524 27344
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30484 26586 30512 27338
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30484 26450 30512 26522
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 30024 26030 30328 26058
rect 29920 25764 29972 25770
rect 29920 25706 29972 25712
rect 29932 25226 29960 25706
rect 29828 25220 29880 25226
rect 29828 25162 29880 25168
rect 29920 25220 29972 25226
rect 29920 25162 29972 25168
rect 29932 24886 29960 24917
rect 29920 24880 29972 24886
rect 30024 24834 30052 26030
rect 30104 25968 30156 25974
rect 30104 25910 30156 25916
rect 30116 25362 30144 25910
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 30208 25498 30236 25842
rect 30300 25838 30328 26030
rect 30288 25832 30340 25838
rect 30288 25774 30340 25780
rect 30196 25492 30248 25498
rect 30196 25434 30248 25440
rect 30104 25356 30156 25362
rect 30104 25298 30156 25304
rect 29972 24828 30052 24834
rect 29920 24822 30052 24828
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29932 24806 30052 24822
rect 29840 23730 29868 24754
rect 29828 23724 29880 23730
rect 29828 23666 29880 23672
rect 29828 23044 29880 23050
rect 29828 22986 29880 22992
rect 29840 22953 29868 22986
rect 29826 22944 29882 22953
rect 29826 22879 29882 22888
rect 29932 22778 29960 24806
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 30024 24274 30052 24686
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 30116 23497 30144 25298
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30288 24880 30340 24886
rect 30288 24822 30340 24828
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 30102 23488 30158 23497
rect 30102 23423 30158 23432
rect 30208 23338 30236 24686
rect 30300 23866 30328 24822
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 30576 23798 30604 24278
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30116 23310 30236 23338
rect 29920 22772 29972 22778
rect 29920 22714 29972 22720
rect 29828 22704 29880 22710
rect 29828 22646 29880 22652
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29734 19816 29790 19825
rect 29734 19751 29790 19760
rect 29748 19718 29776 19751
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29736 19440 29788 19446
rect 29736 19382 29788 19388
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29458 18184 29514 18193
rect 29458 18119 29514 18128
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29380 16998 29408 17070
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29460 16720 29512 16726
rect 29460 16662 29512 16668
rect 29368 14884 29420 14890
rect 29368 14826 29420 14832
rect 29380 14346 29408 14826
rect 29368 14340 29420 14346
rect 29368 14282 29420 14288
rect 29196 12406 29316 12434
rect 29196 11694 29224 12406
rect 29274 12200 29330 12209
rect 29274 12135 29330 12144
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29092 11008 29144 11014
rect 29092 10950 29144 10956
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 28736 9710 28948 9738
rect 28644 9574 28856 9602
rect 28632 9512 28684 9518
rect 28632 9454 28684 9460
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28460 1970 28488 8910
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28552 7206 28580 7822
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28644 7018 28672 9454
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28552 6990 28672 7018
rect 28552 4146 28580 6990
rect 28630 6896 28686 6905
rect 28630 6831 28686 6840
rect 28540 4140 28592 4146
rect 28540 4082 28592 4088
rect 28644 2990 28672 6831
rect 28736 3126 28764 8230
rect 28828 7206 28856 9574
rect 28920 9382 28948 9710
rect 28908 9376 28960 9382
rect 28908 9318 28960 9324
rect 28920 8022 28948 9318
rect 29012 8974 29040 10406
rect 29104 10305 29132 10950
rect 29196 10810 29224 11630
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29090 10296 29146 10305
rect 29090 10231 29146 10240
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 28908 8016 28960 8022
rect 28908 7958 28960 7964
rect 28906 7712 28962 7721
rect 28906 7647 28962 7656
rect 28920 7478 28948 7647
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 28816 7200 28868 7206
rect 28816 7142 28868 7148
rect 28920 6458 28948 7278
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 28724 3120 28776 3126
rect 28724 3062 28776 3068
rect 28632 2984 28684 2990
rect 28632 2926 28684 2932
rect 28448 1964 28500 1970
rect 28448 1906 28500 1912
rect 29012 800 29040 8774
rect 29104 7410 29132 9658
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 29196 6458 29224 8434
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29196 6254 29224 6394
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29184 5364 29236 5370
rect 29288 5352 29316 12135
rect 29380 11218 29408 14282
rect 29472 11665 29500 16662
rect 29656 16522 29684 18294
rect 29748 17746 29776 19382
rect 29840 18970 29868 22646
rect 29920 22500 29972 22506
rect 29920 22442 29972 22448
rect 29932 21418 29960 22442
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 29920 21412 29972 21418
rect 29920 21354 29972 21360
rect 29932 20262 29960 21354
rect 30024 20874 30052 21830
rect 30116 21622 30144 23310
rect 30104 21616 30156 21622
rect 30104 21558 30156 21564
rect 30300 21468 30328 23666
rect 30748 23588 30800 23594
rect 30748 23530 30800 23536
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 30392 22098 30420 22442
rect 30380 22092 30432 22098
rect 30380 22034 30432 22040
rect 30116 21440 30328 21468
rect 30012 20868 30064 20874
rect 30012 20810 30064 20816
rect 30012 20596 30064 20602
rect 30012 20538 30064 20544
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29920 19916 29972 19922
rect 29920 19858 29972 19864
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 29932 18698 29960 19858
rect 30024 19446 30052 20538
rect 30012 19440 30064 19446
rect 30012 19382 30064 19388
rect 30012 19304 30064 19310
rect 30012 19246 30064 19252
rect 30024 19174 30052 19246
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 29920 18692 29972 18698
rect 29920 18634 29972 18640
rect 30116 17762 30144 21440
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30194 21040 30250 21049
rect 30194 20975 30196 20984
rect 30248 20975 30250 20984
rect 30196 20946 30248 20952
rect 30392 20534 30420 21286
rect 30380 20528 30432 20534
rect 30380 20470 30432 20476
rect 30380 20392 30432 20398
rect 30380 20334 30432 20340
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 30208 20058 30236 20198
rect 30392 20058 30420 20334
rect 30196 20052 30248 20058
rect 30196 19994 30248 20000
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30194 19952 30250 19961
rect 30194 19887 30250 19896
rect 30208 19718 30236 19887
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30378 19680 30434 19689
rect 30378 19615 30434 19624
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 30196 18216 30248 18222
rect 30194 18184 30196 18193
rect 30248 18184 30250 18193
rect 30194 18119 30250 18128
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 29932 17734 30144 17762
rect 29644 16516 29696 16522
rect 29644 16458 29696 16464
rect 29552 16176 29604 16182
rect 29552 16118 29604 16124
rect 29564 13190 29592 16118
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29656 14958 29684 16050
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29748 15337 29776 15438
rect 29734 15328 29790 15337
rect 29734 15263 29790 15272
rect 29736 15020 29788 15026
rect 29736 14962 29788 14968
rect 29644 14952 29696 14958
rect 29644 14894 29696 14900
rect 29748 14550 29776 14962
rect 29828 14952 29880 14958
rect 29828 14894 29880 14900
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29840 14346 29868 14894
rect 29932 14890 29960 17734
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 30104 17604 30156 17610
rect 30104 17546 30156 17552
rect 30024 16522 30052 17546
rect 30116 17513 30144 17546
rect 30102 17504 30158 17513
rect 30102 17439 30158 17448
rect 30300 17338 30328 18362
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30104 17264 30156 17270
rect 30104 17206 30156 17212
rect 30012 16516 30064 16522
rect 30012 16458 30064 16464
rect 30116 16250 30144 17206
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30104 16244 30156 16250
rect 30104 16186 30156 16192
rect 30208 15314 30236 16730
rect 30286 15872 30342 15881
rect 30286 15807 30342 15816
rect 30300 15450 30328 15807
rect 30392 15552 30420 19615
rect 30484 19122 30512 23462
rect 30760 22574 30788 23530
rect 30944 23050 30972 25094
rect 31036 24274 31064 26386
rect 31024 24268 31076 24274
rect 31024 24210 31076 24216
rect 31024 23520 31076 23526
rect 31024 23462 31076 23468
rect 30932 23044 30984 23050
rect 30932 22986 30984 22992
rect 31036 22710 31064 23462
rect 31024 22704 31076 22710
rect 31024 22646 31076 22652
rect 30748 22568 30800 22574
rect 30748 22510 30800 22516
rect 30748 22432 30800 22438
rect 30748 22374 30800 22380
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30576 20482 30604 21490
rect 30576 20454 30696 20482
rect 30562 20360 30618 20369
rect 30562 20295 30564 20304
rect 30616 20295 30618 20304
rect 30564 20266 30616 20272
rect 30576 19854 30604 20266
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30668 19174 30696 20454
rect 30656 19168 30708 19174
rect 30484 19094 30604 19122
rect 30656 19110 30708 19116
rect 30470 17640 30526 17649
rect 30470 17575 30472 17584
rect 30524 17575 30526 17584
rect 30472 17546 30524 17552
rect 30470 17504 30526 17513
rect 30470 17439 30526 17448
rect 30484 15706 30512 17439
rect 30576 16114 30604 19094
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30668 17134 30696 18634
rect 30760 17218 30788 22374
rect 30944 21962 30972 22374
rect 30932 21956 30984 21962
rect 30932 21898 30984 21904
rect 31128 21078 31156 28970
rect 31772 27538 31800 34546
rect 33612 33862 33640 37198
rect 34440 37108 34468 39222
rect 34794 39200 34850 39800
rect 36082 39200 36138 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34808 37346 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34808 37318 35020 37346
rect 34992 37262 35020 37318
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 34980 37256 35032 37262
rect 34980 37198 35032 37204
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 34520 37062 34572 37068
rect 33600 33856 33652 33862
rect 33600 33798 33652 33804
rect 34612 33516 34664 33522
rect 34612 33458 34664 33464
rect 33324 32564 33376 32570
rect 33324 32506 33376 32512
rect 33140 32428 33192 32434
rect 33140 32370 33192 32376
rect 33152 28694 33180 32370
rect 33140 28688 33192 28694
rect 33140 28630 33192 28636
rect 32128 28552 32180 28558
rect 32128 28494 32180 28500
rect 31760 27532 31812 27538
rect 31760 27474 31812 27480
rect 31944 26920 31996 26926
rect 31944 26862 31996 26868
rect 31300 26784 31352 26790
rect 31300 26726 31352 26732
rect 31312 26382 31340 26726
rect 31392 26580 31444 26586
rect 31392 26522 31444 26528
rect 31300 26376 31352 26382
rect 31300 26318 31352 26324
rect 31300 24268 31352 24274
rect 31300 24210 31352 24216
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31220 22953 31248 23054
rect 31206 22944 31262 22953
rect 31206 22879 31262 22888
rect 30840 21072 30892 21078
rect 30840 21014 30892 21020
rect 31116 21072 31168 21078
rect 31116 21014 31168 21020
rect 30852 17377 30880 21014
rect 30932 21004 30984 21010
rect 30984 20964 31064 20992
rect 30932 20946 30984 20952
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 30944 19310 30972 20538
rect 31036 20330 31064 20964
rect 31024 20324 31076 20330
rect 31024 20266 31076 20272
rect 31024 19984 31076 19990
rect 31024 19926 31076 19932
rect 30932 19304 30984 19310
rect 30932 19246 30984 19252
rect 31036 18970 31064 19926
rect 31024 18964 31076 18970
rect 31024 18906 31076 18912
rect 31036 18698 31064 18906
rect 31128 18834 31156 21014
rect 31312 20602 31340 24210
rect 31404 22094 31432 26522
rect 31956 26382 31984 26862
rect 31944 26376 31996 26382
rect 31944 26318 31996 26324
rect 31576 26240 31628 26246
rect 31576 26182 31628 26188
rect 31588 25226 31616 26182
rect 31852 25696 31904 25702
rect 31852 25638 31904 25644
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31484 25220 31536 25226
rect 31484 25162 31536 25168
rect 31576 25220 31628 25226
rect 31576 25162 31628 25168
rect 31496 23798 31524 25162
rect 31772 24857 31800 25298
rect 31758 24848 31814 24857
rect 31758 24783 31814 24792
rect 31772 24342 31800 24783
rect 31760 24336 31812 24342
rect 31760 24278 31812 24284
rect 31484 23792 31536 23798
rect 31484 23734 31536 23740
rect 31864 23730 31892 25638
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 31852 23724 31904 23730
rect 31852 23666 31904 23672
rect 31864 23526 31892 23666
rect 31852 23520 31904 23526
rect 31852 23462 31904 23468
rect 31576 23316 31628 23322
rect 31576 23258 31628 23264
rect 31668 23316 31720 23322
rect 31668 23258 31720 23264
rect 31588 22658 31616 23258
rect 31680 22778 31708 23258
rect 32048 23050 32076 24686
rect 32036 23044 32088 23050
rect 32036 22986 32088 22992
rect 31668 22772 31720 22778
rect 31668 22714 31720 22720
rect 31588 22630 31708 22658
rect 31680 22574 31708 22630
rect 31484 22568 31536 22574
rect 31482 22536 31484 22545
rect 31668 22568 31720 22574
rect 31536 22536 31538 22545
rect 31668 22510 31720 22516
rect 31482 22471 31538 22480
rect 31404 22066 31524 22094
rect 31300 20596 31352 20602
rect 31300 20538 31352 20544
rect 31496 20210 31524 22066
rect 31760 22024 31812 22030
rect 31760 21966 31812 21972
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 31588 20505 31616 20538
rect 31574 20496 31630 20505
rect 31574 20431 31630 20440
rect 31496 20182 31708 20210
rect 31298 20088 31354 20097
rect 31298 20023 31354 20032
rect 31206 19816 31262 19825
rect 31312 19786 31340 20023
rect 31574 19816 31630 19825
rect 31206 19751 31208 19760
rect 31260 19751 31262 19760
rect 31300 19780 31352 19786
rect 31208 19722 31260 19728
rect 31574 19751 31630 19760
rect 31300 19722 31352 19728
rect 31220 19666 31248 19722
rect 31392 19712 31444 19718
rect 31220 19660 31392 19666
rect 31220 19654 31444 19660
rect 31220 19638 31432 19654
rect 31588 19514 31616 19751
rect 31576 19508 31628 19514
rect 31576 19450 31628 19456
rect 31680 19394 31708 20182
rect 31772 19553 31800 21966
rect 31852 21548 31904 21554
rect 31852 21490 31904 21496
rect 31758 19544 31814 19553
rect 31758 19479 31814 19488
rect 31496 19366 31708 19394
rect 31116 18828 31168 18834
rect 31116 18770 31168 18776
rect 31024 18692 31076 18698
rect 31024 18634 31076 18640
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30944 18426 30972 18566
rect 30932 18420 30984 18426
rect 30932 18362 30984 18368
rect 30944 17678 30972 18362
rect 31128 18222 31156 18770
rect 31496 18748 31524 19366
rect 31576 19236 31628 19242
rect 31576 19178 31628 19184
rect 31588 19145 31616 19178
rect 31574 19136 31630 19145
rect 31574 19071 31630 19080
rect 31668 18828 31720 18834
rect 31668 18770 31720 18776
rect 31404 18720 31524 18748
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 31300 17604 31352 17610
rect 31404 17592 31432 18720
rect 31576 18216 31628 18222
rect 31352 17564 31432 17592
rect 31496 18176 31576 18204
rect 31300 17546 31352 17552
rect 31116 17536 31168 17542
rect 31116 17478 31168 17484
rect 30838 17368 30894 17377
rect 30838 17303 30894 17312
rect 30760 17190 31064 17218
rect 31036 17134 31064 17190
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 30656 16992 30708 16998
rect 30656 16934 30708 16940
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30564 15972 30616 15978
rect 30564 15914 30616 15920
rect 30472 15700 30524 15706
rect 30472 15642 30524 15648
rect 30392 15524 30512 15552
rect 30300 15422 30420 15450
rect 30024 15286 30236 15314
rect 29920 14884 29972 14890
rect 29920 14826 29972 14832
rect 29828 14340 29880 14346
rect 29828 14282 29880 14288
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29642 12608 29698 12617
rect 29642 12543 29698 12552
rect 29458 11656 29514 11665
rect 29458 11591 29514 11600
rect 29656 11506 29684 12543
rect 29736 12096 29788 12102
rect 29736 12038 29788 12044
rect 29748 11626 29776 12038
rect 29736 11620 29788 11626
rect 29736 11562 29788 11568
rect 29472 11478 29684 11506
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 29472 11098 29500 11478
rect 29642 11384 29698 11393
rect 29642 11319 29698 11328
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 29380 11070 29500 11098
rect 29380 8498 29408 11070
rect 29458 10976 29514 10985
rect 29458 10911 29514 10920
rect 29472 10742 29500 10911
rect 29460 10736 29512 10742
rect 29460 10678 29512 10684
rect 29564 9586 29592 11154
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29472 9110 29500 9318
rect 29460 9104 29512 9110
rect 29460 9046 29512 9052
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 29368 7880 29420 7886
rect 29368 7822 29420 7828
rect 29380 7410 29408 7822
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 29380 6866 29408 7346
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 29380 6322 29408 6802
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 29380 5778 29408 6258
rect 29564 6089 29592 9522
rect 29656 9042 29684 11319
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 29550 6080 29606 6089
rect 29550 6015 29606 6024
rect 29368 5772 29420 5778
rect 29368 5714 29420 5720
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29656 5545 29684 5646
rect 29642 5536 29698 5545
rect 29642 5471 29698 5480
rect 29236 5324 29316 5352
rect 29184 5306 29236 5312
rect 29196 5234 29224 5306
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 29656 4690 29684 5102
rect 29644 4684 29696 4690
rect 29644 4626 29696 4632
rect 29656 4146 29684 4626
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29184 4072 29236 4078
rect 29182 4040 29184 4049
rect 29460 4072 29512 4078
rect 29236 4040 29238 4049
rect 29460 4014 29512 4020
rect 29182 3975 29238 3984
rect 29472 2650 29500 4014
rect 29748 3534 29776 10950
rect 29840 10130 29868 14282
rect 30024 13818 30052 15286
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30116 13954 30144 15098
rect 30196 14340 30248 14346
rect 30196 14282 30248 14288
rect 30208 14074 30236 14282
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30116 13926 30236 13954
rect 30024 13790 30144 13818
rect 30012 13252 30064 13258
rect 30012 13194 30064 13200
rect 29918 11792 29974 11801
rect 30024 11762 30052 13194
rect 29918 11727 29974 11736
rect 30012 11756 30064 11762
rect 29932 11150 29960 11727
rect 30012 11698 30064 11704
rect 30116 11642 30144 13790
rect 30208 12434 30236 13926
rect 30288 13184 30340 13190
rect 30288 13126 30340 13132
rect 30300 12850 30328 13126
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30208 12406 30328 12434
rect 30012 11620 30064 11626
rect 30116 11614 30236 11642
rect 30012 11562 30064 11568
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 29828 10124 29880 10130
rect 29828 10066 29880 10072
rect 29840 9926 29868 10066
rect 29828 9920 29880 9926
rect 29828 9862 29880 9868
rect 29932 9450 29960 10678
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 29826 8392 29882 8401
rect 29826 8327 29882 8336
rect 29840 7002 29868 8327
rect 30024 7834 30052 11562
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30116 10742 30144 11494
rect 30104 10736 30156 10742
rect 30104 10678 30156 10684
rect 29932 7806 30052 7834
rect 29828 6996 29880 7002
rect 29828 6938 29880 6944
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 29840 3890 29868 6394
rect 29932 4078 29960 7806
rect 30012 7744 30064 7750
rect 30012 7686 30064 7692
rect 30024 7002 30052 7686
rect 30012 6996 30064 7002
rect 30012 6938 30064 6944
rect 30208 6361 30236 11614
rect 30300 11218 30328 12406
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30286 10976 30342 10985
rect 30286 10911 30342 10920
rect 30300 10742 30328 10911
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30392 10690 30420 15422
rect 30484 12102 30512 15524
rect 30576 13938 30604 15914
rect 30668 15910 30696 16934
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30668 15094 30696 15302
rect 30656 15088 30708 15094
rect 30656 15030 30708 15036
rect 30656 14272 30708 14278
rect 30656 14214 30708 14220
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30564 13796 30616 13802
rect 30564 13738 30616 13744
rect 30576 12374 30604 13738
rect 30564 12368 30616 12374
rect 30564 12310 30616 12316
rect 30472 12096 30524 12102
rect 30472 12038 30524 12044
rect 30668 11830 30696 14214
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30470 11248 30526 11257
rect 30470 11183 30526 11192
rect 30564 11212 30616 11218
rect 30484 11150 30512 11183
rect 30564 11154 30616 11160
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 30392 10662 30512 10690
rect 30380 10600 30432 10606
rect 30380 10542 30432 10548
rect 30288 10532 30340 10538
rect 30288 10474 30340 10480
rect 30300 9654 30328 10474
rect 30288 9648 30340 9654
rect 30392 9625 30420 10542
rect 30288 9590 30340 9596
rect 30378 9616 30434 9625
rect 30378 9551 30434 9560
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 30300 9042 30328 9454
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 30288 9036 30340 9042
rect 30288 8978 30340 8984
rect 30392 8430 30420 9386
rect 30484 8838 30512 10662
rect 30576 9489 30604 11154
rect 30562 9480 30618 9489
rect 30562 9415 30618 9424
rect 30472 8832 30524 8838
rect 30472 8774 30524 8780
rect 30562 8528 30618 8537
rect 30562 8463 30618 8472
rect 30576 8430 30604 8463
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 30300 6730 30328 8230
rect 30470 8120 30526 8129
rect 30470 8055 30526 8064
rect 30484 7546 30512 8055
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30378 6760 30434 6769
rect 30288 6724 30340 6730
rect 30378 6695 30434 6704
rect 30288 6666 30340 6672
rect 30194 6352 30250 6361
rect 30194 6287 30250 6296
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30116 4729 30144 6054
rect 30286 5944 30342 5953
rect 30286 5879 30342 5888
rect 30300 5642 30328 5879
rect 30392 5817 30420 6695
rect 30562 6624 30618 6633
rect 30562 6559 30618 6568
rect 30378 5808 30434 5817
rect 30378 5743 30434 5752
rect 30288 5636 30340 5642
rect 30288 5578 30340 5584
rect 30470 5536 30526 5545
rect 30470 5471 30526 5480
rect 30194 5400 30250 5409
rect 30194 5335 30250 5344
rect 30208 5302 30236 5335
rect 30196 5296 30248 5302
rect 30196 5238 30248 5244
rect 30378 4856 30434 4865
rect 30378 4791 30434 4800
rect 30102 4720 30158 4729
rect 30102 4655 30158 4664
rect 30286 4312 30342 4321
rect 30286 4247 30288 4256
rect 30340 4247 30342 4256
rect 30288 4218 30340 4224
rect 29920 4072 29972 4078
rect 29920 4014 29972 4020
rect 29840 3862 30052 3890
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29644 3460 29696 3466
rect 29644 3402 29696 3408
rect 29656 2990 29684 3402
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 29920 2984 29972 2990
rect 29920 2926 29972 2932
rect 29656 2854 29684 2926
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29656 2514 29684 2790
rect 29932 2689 29960 2926
rect 29918 2680 29974 2689
rect 29918 2615 29974 2624
rect 29644 2508 29696 2514
rect 29644 2450 29696 2456
rect 30024 2378 30052 3862
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 30012 2372 30064 2378
rect 30012 2314 30064 2320
rect 29932 2106 29960 2314
rect 29920 2100 29972 2106
rect 29920 2042 29972 2048
rect 29644 1624 29696 1630
rect 29644 1566 29696 1572
rect 29656 800 29684 1566
rect 30300 800 30328 3334
rect 30392 2854 30420 4791
rect 30484 4078 30512 5471
rect 30576 4536 30604 6559
rect 30668 6186 30696 11630
rect 30760 11529 30788 17070
rect 31036 16726 31064 17070
rect 31024 16720 31076 16726
rect 31024 16662 31076 16668
rect 30932 16516 30984 16522
rect 30932 16458 30984 16464
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30852 13802 30880 16118
rect 30944 14056 30972 16458
rect 31128 16114 31156 17478
rect 31300 17264 31352 17270
rect 31300 17206 31352 17212
rect 31312 16250 31340 17206
rect 31392 16516 31444 16522
rect 31392 16458 31444 16464
rect 31300 16244 31352 16250
rect 31300 16186 31352 16192
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31022 15736 31078 15745
rect 31022 15671 31078 15680
rect 31036 15502 31064 15671
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 30944 14028 31064 14056
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30840 13796 30892 13802
rect 30840 13738 30892 13744
rect 30840 11552 30892 11558
rect 30746 11520 30802 11529
rect 30840 11494 30892 11500
rect 30746 11455 30802 11464
rect 30746 10840 30802 10849
rect 30746 10775 30802 10784
rect 30760 10742 30788 10775
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30748 10600 30800 10606
rect 30852 10588 30880 11494
rect 30944 11218 30972 13874
rect 31036 12442 31064 14028
rect 31024 12436 31076 12442
rect 31024 12378 31076 12384
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 31128 11098 31156 16050
rect 31404 15978 31432 16458
rect 31392 15972 31444 15978
rect 31392 15914 31444 15920
rect 31496 14346 31524 18176
rect 31576 18158 31628 18164
rect 31576 17604 31628 17610
rect 31576 17546 31628 17552
rect 31588 16266 31616 17546
rect 31680 16794 31708 18770
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 31772 16658 31800 19479
rect 31864 17610 31892 21490
rect 31944 21072 31996 21078
rect 31942 21040 31944 21049
rect 31996 21040 31998 21049
rect 31942 20975 31998 20984
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 31956 20058 31984 20810
rect 31944 20052 31996 20058
rect 31944 19994 31996 20000
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31852 17604 31904 17610
rect 31852 17546 31904 17552
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31588 16250 31800 16266
rect 31588 16244 31812 16250
rect 31588 16238 31760 16244
rect 31760 16186 31812 16192
rect 31668 16108 31720 16114
rect 31668 16050 31720 16056
rect 31576 15496 31628 15502
rect 31576 15438 31628 15444
rect 31484 14340 31536 14346
rect 31484 14282 31536 14288
rect 31588 12434 31616 15438
rect 31404 12406 31616 12434
rect 31404 11914 31432 12406
rect 31576 12368 31628 12374
rect 31576 12310 31628 12316
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31312 11886 31432 11914
rect 31036 11070 31156 11098
rect 31036 10849 31064 11070
rect 31116 11008 31168 11014
rect 31116 10950 31168 10956
rect 31022 10840 31078 10849
rect 31022 10775 31078 10784
rect 30852 10560 30972 10588
rect 30748 10542 30800 10548
rect 30760 9042 30788 10542
rect 30838 10432 30894 10441
rect 30838 10367 30894 10376
rect 30748 9036 30800 9042
rect 30748 8978 30800 8984
rect 30656 6180 30708 6186
rect 30656 6122 30708 6128
rect 30668 5953 30696 6122
rect 30654 5944 30710 5953
rect 30654 5879 30710 5888
rect 30760 5370 30788 8978
rect 30748 5364 30800 5370
rect 30748 5306 30800 5312
rect 30576 4508 30788 4536
rect 30564 4276 30616 4282
rect 30564 4218 30616 4224
rect 30472 4072 30524 4078
rect 30472 4014 30524 4020
rect 30576 3670 30604 4218
rect 30564 3664 30616 3670
rect 30564 3606 30616 3612
rect 30760 3602 30788 4508
rect 30852 4196 30880 10367
rect 30944 8362 30972 10560
rect 31022 10568 31078 10577
rect 31022 10503 31078 10512
rect 31036 9217 31064 10503
rect 31128 10130 31156 10950
rect 31220 10577 31248 11834
rect 31206 10568 31262 10577
rect 31206 10503 31262 10512
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 31220 10266 31248 10406
rect 31208 10260 31260 10266
rect 31208 10202 31260 10208
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31022 9208 31078 9217
rect 31022 9143 31078 9152
rect 31116 9104 31168 9110
rect 31116 9046 31168 9052
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 30932 8356 30984 8362
rect 30932 8298 30984 8304
rect 30932 8016 30984 8022
rect 30932 7958 30984 7964
rect 30944 5692 30972 7958
rect 31036 7721 31064 8366
rect 31022 7712 31078 7721
rect 31022 7647 31078 7656
rect 31128 5710 31156 9046
rect 31206 8256 31262 8265
rect 31206 8191 31262 8200
rect 31116 5704 31168 5710
rect 30944 5664 31064 5692
rect 30932 5092 30984 5098
rect 30932 5034 30984 5040
rect 30944 4321 30972 5034
rect 31036 4554 31064 5664
rect 31116 5646 31168 5652
rect 31024 4548 31076 4554
rect 31024 4490 31076 4496
rect 30930 4312 30986 4321
rect 30930 4247 30986 4256
rect 31220 4214 31248 8191
rect 31312 7206 31340 11886
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31312 6254 31340 7142
rect 31300 6248 31352 6254
rect 31300 6190 31352 6196
rect 31404 5574 31432 11698
rect 31588 11218 31616 12310
rect 31680 11898 31708 16050
rect 31864 15994 31892 16458
rect 31956 16046 31984 19790
rect 32048 18698 32076 22986
rect 32140 21876 32168 28494
rect 33336 27130 33364 32506
rect 33968 28008 34020 28014
rect 33968 27950 34020 27956
rect 33876 27600 33928 27606
rect 33876 27542 33928 27548
rect 33324 27124 33376 27130
rect 33324 27066 33376 27072
rect 33600 26988 33652 26994
rect 33600 26930 33652 26936
rect 33416 25152 33468 25158
rect 33416 25094 33468 25100
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 32220 24132 32272 24138
rect 32220 24074 32272 24080
rect 32232 23866 32260 24074
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 32220 22704 32272 22710
rect 32220 22646 32272 22652
rect 32232 22030 32260 22646
rect 32324 22438 32352 24210
rect 32876 23594 32904 24754
rect 32864 23588 32916 23594
rect 32864 23530 32916 23536
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32312 22432 32364 22438
rect 32312 22374 32364 22380
rect 32324 22166 32352 22374
rect 32312 22160 32364 22166
rect 32312 22102 32364 22108
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32140 21848 32260 21876
rect 32232 21554 32260 21848
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 32324 21298 32352 22102
rect 32494 21992 32550 22001
rect 32494 21927 32496 21936
rect 32548 21927 32550 21936
rect 32496 21898 32548 21904
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32416 21622 32444 21830
rect 32404 21616 32456 21622
rect 32404 21558 32456 21564
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32496 21344 32548 21350
rect 32324 21270 32444 21298
rect 32496 21286 32548 21292
rect 32220 20868 32272 20874
rect 32220 20810 32272 20816
rect 32128 20256 32180 20262
rect 32128 20198 32180 20204
rect 32140 20097 32168 20198
rect 32126 20088 32182 20097
rect 32126 20023 32182 20032
rect 32232 19854 32260 20810
rect 32416 20534 32444 21270
rect 32508 20874 32536 21286
rect 32496 20868 32548 20874
rect 32496 20810 32548 20816
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32324 19689 32352 19790
rect 32404 19712 32456 19718
rect 32310 19680 32366 19689
rect 32404 19654 32456 19660
rect 32310 19615 32366 19624
rect 32416 19446 32444 19654
rect 32404 19440 32456 19446
rect 32310 19408 32366 19417
rect 32404 19382 32456 19388
rect 32310 19343 32312 19352
rect 32364 19343 32366 19352
rect 32312 19314 32364 19320
rect 32404 19168 32456 19174
rect 32404 19110 32456 19116
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 32048 18222 32076 18634
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32036 18216 32088 18222
rect 32036 18158 32088 18164
rect 32220 17604 32272 17610
rect 32220 17546 32272 17552
rect 31772 15966 31892 15994
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 31772 15910 31800 15966
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31772 12102 31800 15846
rect 32232 15094 32260 17546
rect 32324 17338 32352 18566
rect 32416 17814 32444 19110
rect 32404 17808 32456 17814
rect 32404 17750 32456 17756
rect 32600 17626 32628 21490
rect 32692 18329 32720 23462
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32784 20942 32812 21966
rect 32772 20936 32824 20942
rect 32772 20878 32824 20884
rect 32784 19825 32812 20878
rect 32770 19816 32826 19825
rect 32770 19751 32826 19760
rect 32678 18320 32734 18329
rect 32678 18255 32734 18264
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32784 17882 32812 18022
rect 32772 17876 32824 17882
rect 32772 17818 32824 17824
rect 32876 17814 32904 23530
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 33060 23050 33088 23258
rect 33232 23248 33284 23254
rect 33232 23190 33284 23196
rect 33048 23044 33100 23050
rect 33048 22986 33100 22992
rect 33140 22432 33192 22438
rect 33140 22374 33192 22380
rect 33152 22234 33180 22374
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 32954 21856 33010 21865
rect 32954 21791 33010 21800
rect 32968 21554 32996 21791
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 33244 20942 33272 23190
rect 33428 21350 33456 25094
rect 33612 21554 33640 26930
rect 33692 25696 33744 25702
rect 33692 25638 33744 25644
rect 33704 25362 33732 25638
rect 33692 25356 33744 25362
rect 33692 25298 33744 25304
rect 33784 25220 33836 25226
rect 33784 25162 33836 25168
rect 33796 24818 33824 25162
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33888 23882 33916 27542
rect 33980 25158 34008 27950
rect 34520 27328 34572 27334
rect 34520 27270 34572 27276
rect 34532 25906 34560 27270
rect 34624 26586 34652 33458
rect 34704 26920 34756 26926
rect 34704 26862 34756 26868
rect 34612 26580 34664 26586
rect 34612 26522 34664 26528
rect 34716 26234 34744 26862
rect 34624 26206 34744 26234
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34428 25764 34480 25770
rect 34428 25706 34480 25712
rect 34440 25226 34468 25706
rect 34428 25220 34480 25226
rect 34428 25162 34480 25168
rect 33968 25152 34020 25158
rect 33968 25094 34020 25100
rect 34624 24274 34652 26206
rect 34612 24268 34664 24274
rect 34612 24210 34664 24216
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 33704 23854 33916 23882
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33048 20800 33100 20806
rect 33048 20742 33100 20748
rect 32954 20360 33010 20369
rect 32954 20295 32956 20304
rect 33008 20295 33010 20304
rect 32956 20266 33008 20272
rect 32954 20224 33010 20233
rect 32954 20159 33010 20168
rect 32968 19854 32996 20159
rect 33060 19961 33088 20742
rect 33612 20618 33640 21490
rect 33704 20754 33732 23854
rect 33876 23724 33928 23730
rect 33876 23666 33928 23672
rect 33784 23180 33836 23186
rect 33784 23122 33836 23128
rect 33796 22098 33824 23122
rect 33784 22092 33836 22098
rect 33784 22034 33836 22040
rect 33888 21894 33916 23666
rect 33968 22976 34020 22982
rect 33968 22918 34020 22924
rect 33876 21888 33928 21894
rect 33876 21830 33928 21836
rect 33888 20874 33916 21830
rect 33876 20868 33928 20874
rect 33876 20810 33928 20816
rect 33704 20726 33916 20754
rect 33612 20590 33824 20618
rect 33416 20528 33468 20534
rect 33416 20470 33468 20476
rect 33428 20058 33456 20470
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33416 20052 33468 20058
rect 33416 19994 33468 20000
rect 33046 19952 33102 19961
rect 33046 19887 33102 19896
rect 32956 19848 33008 19854
rect 32956 19790 33008 19796
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 33336 19514 33364 19654
rect 33324 19508 33376 19514
rect 33324 19450 33376 19456
rect 33508 19440 33560 19446
rect 33428 19388 33508 19394
rect 33428 19382 33560 19388
rect 33428 19366 33548 19382
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33232 19304 33284 19310
rect 33232 19246 33284 19252
rect 33152 18834 33180 19246
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33046 18320 33102 18329
rect 33046 18255 33048 18264
rect 33100 18255 33102 18264
rect 33048 18226 33100 18232
rect 32864 17808 32916 17814
rect 32864 17750 32916 17756
rect 32416 17598 32628 17626
rect 32312 17332 32364 17338
rect 32312 17274 32364 17280
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32324 16969 32352 17138
rect 32310 16960 32366 16969
rect 32310 16895 32366 16904
rect 32312 15428 32364 15434
rect 32312 15370 32364 15376
rect 32220 15088 32272 15094
rect 32220 15030 32272 15036
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 31668 11892 31720 11898
rect 31668 11834 31720 11840
rect 31576 11212 31628 11218
rect 31576 11154 31628 11160
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 31760 11076 31812 11082
rect 31760 11018 31812 11024
rect 31668 10600 31720 10606
rect 31668 10542 31720 10548
rect 31680 10441 31708 10542
rect 31666 10432 31722 10441
rect 31666 10367 31722 10376
rect 31484 10192 31536 10198
rect 31482 10160 31484 10169
rect 31536 10160 31538 10169
rect 31482 10095 31538 10104
rect 31576 9988 31628 9994
rect 31576 9930 31628 9936
rect 31588 9897 31616 9930
rect 31574 9888 31630 9897
rect 31574 9823 31630 9832
rect 31482 9616 31538 9625
rect 31482 9551 31538 9560
rect 31496 7562 31524 9551
rect 31772 9382 31800 11018
rect 31956 10198 31984 11086
rect 32034 10704 32090 10713
rect 32034 10639 32036 10648
rect 32088 10639 32090 10648
rect 32036 10610 32088 10616
rect 31944 10192 31996 10198
rect 31944 10134 31996 10140
rect 32048 10062 32076 10610
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31864 9194 31892 9454
rect 31772 9166 31892 9194
rect 31942 9208 31998 9217
rect 31772 9042 31800 9166
rect 31942 9143 31998 9152
rect 31760 9036 31812 9042
rect 31760 8978 31812 8984
rect 31852 9036 31904 9042
rect 31852 8978 31904 8984
rect 31864 8945 31892 8978
rect 31850 8936 31906 8945
rect 31850 8871 31906 8880
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31680 8430 31708 8774
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 31668 8288 31720 8294
rect 31666 8256 31668 8265
rect 31720 8256 31722 8265
rect 31956 8242 31984 9143
rect 32034 8664 32090 8673
rect 32034 8599 32090 8608
rect 32048 8566 32076 8599
rect 32036 8560 32088 8566
rect 32036 8502 32088 8508
rect 31666 8191 31722 8200
rect 31864 8214 31984 8242
rect 31680 8044 31800 8072
rect 31680 7954 31708 8044
rect 31668 7948 31720 7954
rect 31668 7890 31720 7896
rect 31576 7744 31628 7750
rect 31574 7712 31576 7721
rect 31668 7744 31720 7750
rect 31628 7712 31630 7721
rect 31668 7686 31720 7692
rect 31574 7647 31630 7656
rect 31496 7546 31616 7562
rect 31496 7540 31628 7546
rect 31496 7534 31576 7540
rect 31576 7482 31628 7488
rect 31482 7168 31538 7177
rect 31482 7103 31538 7112
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 31404 5166 31432 5510
rect 31496 5409 31524 7103
rect 31574 7032 31630 7041
rect 31574 6967 31630 6976
rect 31588 6662 31616 6967
rect 31680 6798 31708 7686
rect 31772 7290 31800 8044
rect 31864 7410 31892 8214
rect 31944 8084 31996 8090
rect 31944 8026 31996 8032
rect 32036 8084 32088 8090
rect 32036 8026 32088 8032
rect 31852 7404 31904 7410
rect 31852 7346 31904 7352
rect 31772 7262 31892 7290
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31576 6656 31628 6662
rect 31576 6598 31628 6604
rect 31864 6202 31892 7262
rect 31956 7041 31984 8026
rect 32048 7478 32076 8026
rect 32036 7472 32088 7478
rect 32036 7414 32088 7420
rect 32036 7200 32088 7206
rect 32036 7142 32088 7148
rect 31942 7032 31998 7041
rect 31942 6967 31998 6976
rect 31956 6322 31984 6967
rect 32048 6390 32076 7142
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 31944 6316 31996 6322
rect 31944 6258 31996 6264
rect 31864 6174 31984 6202
rect 31576 6112 31628 6118
rect 31576 6054 31628 6060
rect 31760 6112 31812 6118
rect 31760 6054 31812 6060
rect 31588 5681 31616 6054
rect 31772 5846 31800 6054
rect 31760 5840 31812 5846
rect 31760 5782 31812 5788
rect 31574 5672 31630 5681
rect 31574 5607 31630 5616
rect 31758 5672 31814 5681
rect 31758 5607 31814 5616
rect 31576 5568 31628 5574
rect 31576 5510 31628 5516
rect 31482 5400 31538 5409
rect 31588 5370 31616 5510
rect 31482 5335 31538 5344
rect 31576 5364 31628 5370
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31208 4208 31260 4214
rect 30852 4168 30972 4196
rect 30944 3602 30972 4168
rect 31208 4150 31260 4156
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 30748 3596 30800 3602
rect 30748 3538 30800 3544
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30760 3398 30788 3538
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 31312 3194 31340 3878
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31496 2990 31524 5335
rect 31576 5306 31628 5312
rect 31574 5264 31630 5273
rect 31574 5199 31630 5208
rect 31588 4282 31616 5199
rect 31772 5030 31800 5607
rect 31850 5400 31906 5409
rect 31850 5335 31906 5344
rect 31864 5302 31892 5335
rect 31956 5302 31984 6174
rect 32140 5896 32168 12038
rect 32324 11694 32352 15370
rect 32416 12714 32444 17598
rect 32680 16720 32732 16726
rect 32680 16662 32732 16668
rect 32588 16516 32640 16522
rect 32588 16458 32640 16464
rect 32600 15706 32628 16458
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32404 12708 32456 12714
rect 32404 12650 32456 12656
rect 32600 11898 32628 15302
rect 32692 12102 32720 16662
rect 32772 15632 32824 15638
rect 32772 15574 32824 15580
rect 32680 12096 32732 12102
rect 32680 12038 32732 12044
rect 32588 11892 32640 11898
rect 32588 11834 32640 11840
rect 32680 11824 32732 11830
rect 32680 11766 32732 11772
rect 32312 11688 32364 11694
rect 32312 11630 32364 11636
rect 32218 10296 32274 10305
rect 32218 10231 32220 10240
rect 32272 10231 32274 10240
rect 32220 10202 32272 10208
rect 32220 9376 32272 9382
rect 32220 9318 32272 9324
rect 32232 7206 32260 9318
rect 32324 7800 32352 11630
rect 32588 11076 32640 11082
rect 32588 11018 32640 11024
rect 32600 10810 32628 11018
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32416 8634 32444 10746
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32508 8022 32536 10202
rect 32588 9988 32640 9994
rect 32588 9930 32640 9936
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32324 7772 32444 7800
rect 32416 7698 32444 7772
rect 32416 7670 32536 7698
rect 32220 7200 32272 7206
rect 32220 7142 32272 7148
rect 32404 6860 32456 6866
rect 32404 6802 32456 6808
rect 32310 6624 32366 6633
rect 32310 6559 32366 6568
rect 32324 6474 32352 6559
rect 32232 6446 32352 6474
rect 32232 6254 32260 6446
rect 32312 6384 32364 6390
rect 32416 6361 32444 6802
rect 32312 6326 32364 6332
rect 32402 6352 32458 6361
rect 32220 6248 32272 6254
rect 32220 6190 32272 6196
rect 32324 5914 32352 6326
rect 32402 6287 32458 6296
rect 32508 6254 32536 7670
rect 32600 7478 32628 9930
rect 32692 8809 32720 11766
rect 32784 11014 32812 15574
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32770 9208 32826 9217
rect 32770 9143 32826 9152
rect 32784 8974 32812 9143
rect 32772 8968 32824 8974
rect 32772 8910 32824 8916
rect 32678 8800 32734 8809
rect 32678 8735 32734 8744
rect 32770 8664 32826 8673
rect 32770 8599 32826 8608
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32588 7472 32640 7478
rect 32588 7414 32640 7420
rect 32496 6248 32548 6254
rect 32496 6190 32548 6196
rect 32312 5908 32364 5914
rect 32140 5868 32260 5896
rect 32126 5808 32182 5817
rect 32126 5743 32182 5752
rect 32140 5370 32168 5743
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 31852 5296 31904 5302
rect 31852 5238 31904 5244
rect 31944 5296 31996 5302
rect 31944 5238 31996 5244
rect 32232 5166 32260 5868
rect 32312 5850 32364 5856
rect 32496 5568 32548 5574
rect 32496 5510 32548 5516
rect 32310 5264 32366 5273
rect 32310 5199 32366 5208
rect 32220 5160 32272 5166
rect 32218 5128 32220 5137
rect 32272 5128 32274 5137
rect 32324 5098 32352 5199
rect 32508 5166 32536 5510
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32588 5160 32640 5166
rect 32588 5102 32640 5108
rect 32218 5063 32274 5072
rect 32312 5092 32364 5098
rect 32312 5034 32364 5040
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 32600 4842 32628 5102
rect 32232 4814 32628 4842
rect 31852 4548 31904 4554
rect 31852 4490 31904 4496
rect 31864 4282 31892 4490
rect 31576 4276 31628 4282
rect 31576 4218 31628 4224
rect 31852 4276 31904 4282
rect 31852 4218 31904 4224
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 31576 2848 31628 2854
rect 31576 2790 31628 2796
rect 31298 2544 31354 2553
rect 31298 2479 31354 2488
rect 31312 2378 31340 2479
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 31588 800 31616 2790
rect 32232 800 32260 4814
rect 32312 4684 32364 4690
rect 32312 4626 32364 4632
rect 32324 4214 32352 4626
rect 32692 4570 32720 8434
rect 32508 4554 32720 4570
rect 32496 4548 32720 4554
rect 32548 4542 32720 4548
rect 32496 4490 32548 4496
rect 32588 4480 32640 4486
rect 32588 4422 32640 4428
rect 32600 4282 32628 4422
rect 32588 4276 32640 4282
rect 32588 4218 32640 4224
rect 32680 4276 32732 4282
rect 32680 4218 32732 4224
rect 32312 4208 32364 4214
rect 32312 4150 32364 4156
rect 32324 2990 32352 4150
rect 32586 3768 32642 3777
rect 32586 3703 32642 3712
rect 32600 3602 32628 3703
rect 32588 3596 32640 3602
rect 32588 3538 32640 3544
rect 32600 3097 32628 3538
rect 32692 3126 32720 4218
rect 32680 3120 32732 3126
rect 32586 3088 32642 3097
rect 32680 3062 32732 3068
rect 32586 3023 32642 3032
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 32324 2514 32352 2926
rect 32312 2508 32364 2514
rect 32312 2450 32364 2456
rect 32784 2106 32812 8599
rect 32876 8129 32904 17750
rect 33152 17626 33180 18770
rect 33244 18154 33272 19246
rect 33232 18148 33284 18154
rect 33232 18090 33284 18096
rect 33244 17746 33272 18090
rect 33232 17740 33284 17746
rect 33232 17682 33284 17688
rect 33324 17672 33376 17678
rect 33152 17598 33272 17626
rect 33324 17614 33376 17620
rect 33048 17536 33100 17542
rect 33048 17478 33100 17484
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 33060 17338 33088 17478
rect 33048 17332 33100 17338
rect 33048 17274 33100 17280
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 32968 13025 32996 17138
rect 33152 15978 33180 17478
rect 33140 15972 33192 15978
rect 33140 15914 33192 15920
rect 33244 15586 33272 17598
rect 33152 15570 33272 15586
rect 33140 15564 33272 15570
rect 33192 15558 33272 15564
rect 33140 15506 33192 15512
rect 33048 14408 33100 14414
rect 33048 14350 33100 14356
rect 32954 13016 33010 13025
rect 32954 12951 33010 12960
rect 33060 9586 33088 14350
rect 33336 12889 33364 17614
rect 33428 15162 33456 19366
rect 33508 19236 33560 19242
rect 33508 19178 33560 19184
rect 33520 18290 33548 19178
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 33508 16516 33560 16522
rect 33508 16458 33560 16464
rect 33520 16046 33548 16458
rect 33508 16040 33560 16046
rect 33508 15982 33560 15988
rect 33416 15156 33468 15162
rect 33416 15098 33468 15104
rect 33322 12880 33378 12889
rect 33140 12844 33192 12850
rect 33322 12815 33378 12824
rect 33140 12786 33192 12792
rect 33152 10674 33180 12786
rect 33508 12164 33560 12170
rect 33508 12106 33560 12112
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 33152 9586 33180 10610
rect 33416 10464 33468 10470
rect 33416 10406 33468 10412
rect 33324 10056 33376 10062
rect 33324 9998 33376 10004
rect 33336 9897 33364 9998
rect 33322 9888 33378 9897
rect 33322 9823 33378 9832
rect 33048 9580 33100 9586
rect 33048 9522 33100 9528
rect 33140 9580 33192 9586
rect 33140 9522 33192 9528
rect 33060 9466 33088 9522
rect 33324 9512 33376 9518
rect 33060 9438 33180 9466
rect 33324 9454 33376 9460
rect 33152 9382 33180 9438
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 33230 9072 33286 9081
rect 33230 9007 33286 9016
rect 33244 8974 33272 9007
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 33140 8900 33192 8906
rect 33140 8842 33192 8848
rect 32956 8628 33008 8634
rect 32956 8570 33008 8576
rect 32862 8120 32918 8129
rect 32862 8055 32918 8064
rect 32968 7313 32996 8570
rect 33152 8090 33180 8842
rect 33230 8800 33286 8809
rect 33230 8735 33286 8744
rect 33244 8498 33272 8735
rect 33232 8492 33284 8498
rect 33232 8434 33284 8440
rect 33140 8084 33192 8090
rect 33140 8026 33192 8032
rect 33244 7886 33272 8434
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 33138 7712 33194 7721
rect 33138 7647 33194 7656
rect 33152 7410 33180 7647
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 32954 7304 33010 7313
rect 32864 7268 32916 7274
rect 32954 7239 33010 7248
rect 32864 7210 32916 7216
rect 32876 6730 32904 7210
rect 32954 7032 33010 7041
rect 32954 6967 33010 6976
rect 32968 6798 32996 6967
rect 32956 6792 33008 6798
rect 32956 6734 33008 6740
rect 32864 6724 32916 6730
rect 32864 6666 32916 6672
rect 33152 5846 33180 7346
rect 33336 7206 33364 9454
rect 33324 7200 33376 7206
rect 33324 7142 33376 7148
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 33140 5840 33192 5846
rect 33140 5782 33192 5788
rect 33060 5370 33088 5782
rect 33048 5364 33100 5370
rect 33048 5306 33100 5312
rect 32862 4992 32918 5001
rect 32862 4927 32918 4936
rect 32876 4690 32904 4927
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 33428 4214 33456 10406
rect 33520 8974 33548 12106
rect 33704 11665 33732 20402
rect 33796 16561 33824 20590
rect 33782 16552 33838 16561
rect 33782 16487 33838 16496
rect 33888 13326 33916 20726
rect 33980 18426 34008 22918
rect 34072 20534 34100 24006
rect 34808 23866 34836 37198
rect 36096 37126 36124 39200
rect 36174 38176 36230 38185
rect 36174 38111 36230 38120
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35452 35894 35480 37062
rect 36188 36922 36216 38111
rect 36268 37256 36320 37262
rect 36268 37198 36320 37204
rect 36176 36916 36228 36922
rect 36176 36858 36228 36864
rect 35532 36780 35584 36786
rect 35532 36722 35584 36728
rect 35544 36582 35572 36722
rect 35532 36576 35584 36582
rect 35532 36518 35584 36524
rect 35360 35866 35480 35894
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30190 35388 35866
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 35348 30184 35400 30190
rect 35348 30126 35400 30132
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35348 26852 35400 26858
rect 35348 26794 35400 26800
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 24818 35388 26794
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34532 22098 34560 23598
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35360 22642 35388 23054
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34520 22092 34572 22098
rect 34520 22034 34572 22040
rect 34336 21344 34388 21350
rect 34336 21286 34388 21292
rect 34348 21010 34376 21286
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34060 20528 34112 20534
rect 34060 20470 34112 20476
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 34164 19938 34192 20402
rect 34164 19910 34284 19938
rect 34624 19922 34652 22510
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34152 19848 34204 19854
rect 34152 19790 34204 19796
rect 34060 19440 34112 19446
rect 34060 19382 34112 19388
rect 34072 18698 34100 19382
rect 34060 18692 34112 18698
rect 34060 18634 34112 18640
rect 33968 18420 34020 18426
rect 33968 18362 34020 18368
rect 33968 17672 34020 17678
rect 33968 17614 34020 17620
rect 33980 16697 34008 17614
rect 33966 16688 34022 16697
rect 33966 16623 34022 16632
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 34072 16250 34100 16390
rect 34060 16244 34112 16250
rect 34060 16186 34112 16192
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 34164 12782 34192 19790
rect 34256 13161 34284 19910
rect 34612 19916 34664 19922
rect 34612 19858 34664 19864
rect 34796 19848 34848 19854
rect 34796 19790 34848 19796
rect 34428 19780 34480 19786
rect 34428 19722 34480 19728
rect 34440 18970 34468 19722
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34532 17814 34560 19314
rect 34716 18766 34744 19654
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34520 17808 34572 17814
rect 34520 17750 34572 17756
rect 34808 17270 34836 19790
rect 35360 19718 35388 22578
rect 35452 21078 35480 31282
rect 35544 29034 35572 36518
rect 35532 29028 35584 29034
rect 35532 28970 35584 28976
rect 35440 21072 35492 21078
rect 35440 21014 35492 21020
rect 35900 20868 35952 20874
rect 35900 20810 35952 20816
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34888 18896 34940 18902
rect 34888 18838 34940 18844
rect 34900 18426 34928 18838
rect 35912 18834 35940 20810
rect 36280 19514 36308 37198
rect 36740 36922 36768 39200
rect 36818 38856 36874 38865
rect 36818 38791 36874 38800
rect 36728 36916 36780 36922
rect 36728 36858 36780 36864
rect 36832 36786 36860 38791
rect 38028 37330 38056 39200
rect 38016 37324 38068 37330
rect 38016 37266 38068 37272
rect 37096 37120 37148 37126
rect 37096 37062 37148 37068
rect 36820 36780 36872 36786
rect 36820 36722 36872 36728
rect 36820 36576 36872 36582
rect 36820 36518 36872 36524
rect 36832 36310 36860 36518
rect 36820 36304 36872 36310
rect 36820 36246 36872 36252
rect 36544 36168 36596 36174
rect 36544 36110 36596 36116
rect 36360 22024 36412 22030
rect 36360 21966 36412 21972
rect 36372 21554 36400 21966
rect 36556 21894 36584 36110
rect 37108 36106 37136 37062
rect 38290 36816 38346 36825
rect 38290 36751 38346 36760
rect 37372 36644 37424 36650
rect 37372 36586 37424 36592
rect 37188 36168 37240 36174
rect 37188 36110 37240 36116
rect 37096 36100 37148 36106
rect 37096 36042 37148 36048
rect 36728 35692 36780 35698
rect 36728 35634 36780 35640
rect 36740 33658 36768 35634
rect 37200 35290 37228 36110
rect 37188 35284 37240 35290
rect 37188 35226 37240 35232
rect 37384 35086 37412 36586
rect 37648 36576 37700 36582
rect 37648 36518 37700 36524
rect 37556 36100 37608 36106
rect 37556 36042 37608 36048
rect 37372 35080 37424 35086
rect 37372 35022 37424 35028
rect 37464 34944 37516 34950
rect 37464 34886 37516 34892
rect 37188 34536 37240 34542
rect 37188 34478 37240 34484
rect 37200 34105 37228 34478
rect 37186 34096 37242 34105
rect 37186 34031 37242 34040
rect 36728 33652 36780 33658
rect 36728 33594 36780 33600
rect 37476 32609 37504 34886
rect 37462 32600 37518 32609
rect 37462 32535 37518 32544
rect 37464 32360 37516 32366
rect 37464 32302 37516 32308
rect 37476 32065 37504 32302
rect 37462 32056 37518 32065
rect 37462 31991 37518 32000
rect 37188 29096 37240 29102
rect 37188 29038 37240 29044
rect 37200 28665 37228 29038
rect 37186 28656 37242 28665
rect 37186 28591 37242 28600
rect 37280 26784 37332 26790
rect 37280 26726 37332 26732
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 34888 18420 34940 18426
rect 34888 18362 34940 18368
rect 35624 18284 35676 18290
rect 35624 18226 35676 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35636 17338 35664 18226
rect 35624 17332 35676 17338
rect 35624 17274 35676 17280
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 34532 15434 34560 15982
rect 34520 15428 34572 15434
rect 34520 15370 34572 15376
rect 34242 13152 34298 13161
rect 34242 13087 34298 13096
rect 34520 12980 34572 12986
rect 34520 12922 34572 12928
rect 34532 12889 34560 12922
rect 34518 12880 34574 12889
rect 34518 12815 34574 12824
rect 34152 12776 34204 12782
rect 34152 12718 34204 12724
rect 33690 11656 33746 11665
rect 33690 11591 33746 11600
rect 34060 11076 34112 11082
rect 34060 11018 34112 11024
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 33612 10169 33640 10202
rect 33598 10160 33654 10169
rect 33598 10095 33654 10104
rect 33692 10056 33744 10062
rect 33612 10016 33692 10044
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33612 8820 33640 10016
rect 33692 9998 33744 10004
rect 33784 9920 33836 9926
rect 33784 9862 33836 9868
rect 33692 9444 33744 9450
rect 33692 9386 33744 9392
rect 33520 8792 33640 8820
rect 33520 7886 33548 8792
rect 33704 8673 33732 9386
rect 33690 8664 33746 8673
rect 33690 8599 33746 8608
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33598 7848 33654 7857
rect 33598 7783 33600 7792
rect 33652 7783 33654 7792
rect 33600 7754 33652 7760
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 33520 7188 33548 7346
rect 33692 7336 33744 7342
rect 33692 7278 33744 7284
rect 33520 7160 33640 7188
rect 33506 6896 33562 6905
rect 33506 6831 33562 6840
rect 33520 6322 33548 6831
rect 33508 6316 33560 6322
rect 33508 6258 33560 6264
rect 33612 4486 33640 7160
rect 33704 7002 33732 7278
rect 33692 6996 33744 7002
rect 33692 6938 33744 6944
rect 33796 6798 33824 9862
rect 33876 9376 33928 9382
rect 33876 9318 33928 9324
rect 33888 8974 33916 9318
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33876 8356 33928 8362
rect 33876 8298 33928 8304
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 33784 6656 33836 6662
rect 33784 6598 33836 6604
rect 33690 6352 33746 6361
rect 33796 6322 33824 6598
rect 33690 6287 33746 6296
rect 33784 6316 33836 6322
rect 33704 4622 33732 6287
rect 33784 6258 33836 6264
rect 33784 5840 33836 5846
rect 33784 5782 33836 5788
rect 33796 4826 33824 5782
rect 33888 5409 33916 8298
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33874 5400 33930 5409
rect 33874 5335 33930 5344
rect 33784 4820 33836 4826
rect 33784 4762 33836 4768
rect 33980 4706 34008 8026
rect 34072 7750 34100 11018
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34152 10056 34204 10062
rect 34152 9998 34204 10004
rect 34164 9722 34192 9998
rect 34242 9888 34298 9897
rect 34242 9823 34298 9832
rect 34152 9716 34204 9722
rect 34152 9658 34204 9664
rect 34256 9586 34284 9823
rect 34532 9654 34560 10134
rect 34612 9920 34664 9926
rect 34612 9862 34664 9868
rect 34520 9648 34572 9654
rect 34520 9590 34572 9596
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 34060 7744 34112 7750
rect 34060 7686 34112 7692
rect 34058 7576 34114 7585
rect 34058 7511 34060 7520
rect 34112 7511 34114 7520
rect 34060 7482 34112 7488
rect 34164 7206 34192 9522
rect 34256 9042 34284 9522
rect 34336 9376 34388 9382
rect 34336 9318 34388 9324
rect 34348 9178 34376 9318
rect 34336 9172 34388 9178
rect 34336 9114 34388 9120
rect 34244 9036 34296 9042
rect 34244 8978 34296 8984
rect 34440 8401 34468 9522
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34532 8498 34560 8910
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34426 8392 34482 8401
rect 34426 8327 34482 8336
rect 34520 8356 34572 8362
rect 34520 8298 34572 8304
rect 34244 8288 34296 8294
rect 34244 8230 34296 8236
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34256 8022 34284 8230
rect 34440 8090 34468 8230
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34244 8016 34296 8022
rect 34244 7958 34296 7964
rect 34244 7880 34296 7886
rect 34244 7822 34296 7828
rect 34152 7200 34204 7206
rect 34256 7177 34284 7822
rect 34152 7142 34204 7148
rect 34242 7168 34298 7177
rect 34242 7103 34298 7112
rect 34060 6996 34112 7002
rect 34060 6938 34112 6944
rect 34072 6662 34100 6938
rect 34428 6928 34480 6934
rect 34428 6870 34480 6876
rect 34336 6792 34388 6798
rect 34336 6734 34388 6740
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 34244 6656 34296 6662
rect 34244 6598 34296 6604
rect 34152 6248 34204 6254
rect 34152 6190 34204 6196
rect 34058 5128 34114 5137
rect 34058 5063 34114 5072
rect 33796 4678 34008 4706
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 33416 4208 33468 4214
rect 33416 4150 33468 4156
rect 33508 3936 33560 3942
rect 33336 3896 33508 3924
rect 33336 3482 33364 3896
rect 33508 3878 33560 3884
rect 33152 3466 33364 3482
rect 33140 3460 33364 3466
rect 33192 3454 33364 3460
rect 33140 3402 33192 3408
rect 33612 2990 33640 4422
rect 33796 3942 33824 4678
rect 33876 4548 33928 4554
rect 33876 4490 33928 4496
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 33520 870 33640 898
rect 33520 800 33548 870
rect 25240 734 25544 762
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 29642 200 29698 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 33612 762 33640 870
rect 33888 762 33916 4490
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 33980 3466 34008 3878
rect 34072 3466 34100 5063
rect 34164 4146 34192 6190
rect 34256 4865 34284 6598
rect 34348 5681 34376 6734
rect 34440 6390 34468 6870
rect 34428 6384 34480 6390
rect 34428 6326 34480 6332
rect 34532 5794 34560 8298
rect 34440 5766 34560 5794
rect 34334 5672 34390 5681
rect 34334 5607 34390 5616
rect 34334 5536 34390 5545
rect 34334 5471 34390 5480
rect 34242 4856 34298 4865
rect 34242 4791 34298 4800
rect 34348 4690 34376 5471
rect 34336 4684 34388 4690
rect 34336 4626 34388 4632
rect 34244 4616 34296 4622
rect 34244 4558 34296 4564
rect 34152 4140 34204 4146
rect 34152 4082 34204 4088
rect 33968 3460 34020 3466
rect 33968 3402 34020 3408
rect 34060 3460 34112 3466
rect 34060 3402 34112 3408
rect 34152 2916 34204 2922
rect 34152 2858 34204 2864
rect 34060 2848 34112 2854
rect 34060 2790 34112 2796
rect 34072 2038 34100 2790
rect 34060 2032 34112 2038
rect 34060 1974 34112 1980
rect 34164 800 34192 2858
rect 34256 2650 34284 4558
rect 34440 4264 34468 5766
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34348 4236 34468 4264
rect 34348 3602 34376 4236
rect 34532 4162 34560 5646
rect 34440 4134 34560 4162
rect 34440 4078 34468 4134
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34336 3596 34388 3602
rect 34336 3538 34388 3544
rect 34426 3360 34482 3369
rect 34426 3295 34482 3304
rect 34440 3126 34468 3295
rect 34624 3126 34652 9862
rect 34716 8090 34744 16730
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35716 15428 35768 15434
rect 35716 15370 35768 15376
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34808 12442 34836 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 12436 34848 12442
rect 34796 12378 34848 12384
rect 35348 11824 35400 11830
rect 35348 11766 35400 11772
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9376 34848 9382
rect 34796 9318 34848 9324
rect 34808 8922 34836 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34980 9104 35032 9110
rect 34980 9046 35032 9052
rect 34808 8894 34928 8922
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34716 6866 34744 7414
rect 34704 6860 34756 6866
rect 34704 6802 34756 6808
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34716 5846 34744 6598
rect 34808 6361 34836 8774
rect 34900 8362 34928 8894
rect 34992 8634 35020 9046
rect 35256 8900 35308 8906
rect 35256 8842 35308 8848
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 35268 8362 35296 8842
rect 34888 8356 34940 8362
rect 34888 8298 34940 8304
rect 35256 8356 35308 8362
rect 35256 8298 35308 8304
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35268 7478 35296 7686
rect 35256 7472 35308 7478
rect 35256 7414 35308 7420
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34794 6352 34850 6361
rect 34794 6287 34850 6296
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34704 5840 34756 5846
rect 34704 5782 34756 5788
rect 35072 5840 35124 5846
rect 35072 5782 35124 5788
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 34716 4434 34744 5510
rect 35084 5302 35112 5782
rect 35360 5642 35388 11766
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35440 10056 35492 10062
rect 35440 9998 35492 10004
rect 35452 8498 35480 9998
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35440 8356 35492 8362
rect 35440 8298 35492 8304
rect 35452 6662 35480 8298
rect 35440 6656 35492 6662
rect 35440 6598 35492 6604
rect 35440 6248 35492 6254
rect 35440 6190 35492 6196
rect 35452 5778 35480 6190
rect 35440 5772 35492 5778
rect 35440 5714 35492 5720
rect 35544 5658 35572 10406
rect 35636 10033 35664 10610
rect 35622 10024 35678 10033
rect 35622 9959 35678 9968
rect 35728 8974 35756 15370
rect 35992 13184 36044 13190
rect 35992 13126 36044 13132
rect 35898 12200 35954 12209
rect 35898 12135 35954 12144
rect 35912 11150 35940 12135
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 35900 10464 35952 10470
rect 35900 10406 35952 10412
rect 35808 9988 35860 9994
rect 35808 9930 35860 9936
rect 35820 9586 35848 9930
rect 35808 9580 35860 9586
rect 35808 9522 35860 9528
rect 35716 8968 35768 8974
rect 35716 8910 35768 8916
rect 35624 8424 35676 8430
rect 35624 8366 35676 8372
rect 35636 8090 35664 8366
rect 35624 8084 35676 8090
rect 35624 8026 35676 8032
rect 35728 7954 35756 8910
rect 35808 8900 35860 8906
rect 35808 8842 35860 8848
rect 35716 7948 35768 7954
rect 35716 7890 35768 7896
rect 35716 7744 35768 7750
rect 35716 7686 35768 7692
rect 35624 7540 35676 7546
rect 35624 7482 35676 7488
rect 35636 7206 35664 7482
rect 35728 7449 35756 7686
rect 35714 7440 35770 7449
rect 35714 7375 35770 7384
rect 35716 7336 35768 7342
rect 35716 7278 35768 7284
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35636 6798 35664 7142
rect 35728 6866 35756 7278
rect 35716 6860 35768 6866
rect 35716 6802 35768 6808
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35624 6656 35676 6662
rect 35624 6598 35676 6604
rect 35716 6656 35768 6662
rect 35716 6598 35768 6604
rect 35636 6118 35664 6598
rect 35728 6497 35756 6598
rect 35714 6488 35770 6497
rect 35714 6423 35770 6432
rect 35820 6361 35848 8842
rect 35806 6352 35862 6361
rect 35806 6287 35862 6296
rect 35716 6248 35768 6254
rect 35716 6190 35768 6196
rect 35624 6112 35676 6118
rect 35624 6054 35676 6060
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 35452 5630 35572 5658
rect 35624 5704 35676 5710
rect 35624 5646 35676 5652
rect 35072 5296 35124 5302
rect 35072 5238 35124 5244
rect 34888 5160 34940 5166
rect 34886 5128 34888 5137
rect 34940 5128 34942 5137
rect 34886 5063 34942 5072
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34716 4406 34836 4434
rect 34704 4072 34756 4078
rect 34704 4014 34756 4020
rect 34428 3120 34480 3126
rect 34428 3062 34480 3068
rect 34612 3120 34664 3126
rect 34612 3062 34664 3068
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 34716 2378 34744 4014
rect 34808 3126 34836 4406
rect 35452 4078 35480 5630
rect 35532 5568 35584 5574
rect 35532 5510 35584 5516
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 35348 4004 35400 4010
rect 35348 3946 35400 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35256 3596 35308 3602
rect 35256 3538 35308 3544
rect 35268 3505 35296 3538
rect 35254 3496 35310 3505
rect 35360 3466 35388 3946
rect 35254 3431 35310 3440
rect 35348 3460 35400 3466
rect 35348 3402 35400 3408
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34808 2961 34836 3062
rect 34794 2952 34850 2961
rect 34794 2887 34850 2896
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 34704 2372 34756 2378
rect 34704 2314 34756 2320
rect 34808 800 34836 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35544 2514 35572 5510
rect 35636 5030 35664 5646
rect 35624 5024 35676 5030
rect 35624 4966 35676 4972
rect 35624 4072 35676 4078
rect 35622 4040 35624 4049
rect 35676 4040 35678 4049
rect 35622 3975 35678 3984
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 35728 1465 35756 6190
rect 35808 4480 35860 4486
rect 35808 4422 35860 4428
rect 35820 2825 35848 4422
rect 35912 4146 35940 10406
rect 36004 4146 36032 13126
rect 36176 12096 36228 12102
rect 36176 12038 36228 12044
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 36096 11121 36124 11698
rect 36082 11112 36138 11121
rect 36082 11047 36138 11056
rect 36084 11008 36136 11014
rect 36084 10950 36136 10956
rect 36096 7954 36124 10950
rect 36188 8498 36216 12038
rect 36268 11212 36320 11218
rect 36268 11154 36320 11160
rect 36280 10130 36308 11154
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 36280 8566 36308 10066
rect 36268 8560 36320 8566
rect 36268 8502 36320 8508
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36084 7948 36136 7954
rect 36136 7908 36216 7936
rect 36084 7890 36136 7896
rect 36188 7290 36216 7908
rect 36096 7262 36216 7290
rect 36096 6934 36124 7262
rect 36280 7002 36308 8298
rect 36268 6996 36320 7002
rect 36268 6938 36320 6944
rect 36084 6928 36136 6934
rect 36084 6870 36136 6876
rect 36096 6322 36124 6870
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 36266 6760 36322 6769
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 36188 5817 36216 6734
rect 36266 6695 36322 6704
rect 36174 5808 36230 5817
rect 36174 5743 36230 5752
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 36280 4010 36308 6695
rect 36268 4004 36320 4010
rect 36268 3946 36320 3952
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 35806 2816 35862 2825
rect 35806 2751 35862 2760
rect 35714 1456 35770 1465
rect 35714 1391 35770 1400
rect 36096 800 36124 3878
rect 36372 3058 36400 21490
rect 37292 21146 37320 26726
rect 37568 26234 37596 36042
rect 37476 26206 37596 26234
rect 37476 24410 37504 26206
rect 37660 25430 37688 36518
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38304 35834 38332 36751
rect 38672 36378 38700 39200
rect 39316 37126 39344 39200
rect 39304 37120 39356 37126
rect 39304 37062 39356 37068
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 38292 35828 38344 35834
rect 38292 35770 38344 35776
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38200 31952 38252 31958
rect 38200 31894 38252 31900
rect 38016 31816 38068 31822
rect 38016 31758 38068 31764
rect 38028 31482 38056 31758
rect 38016 31476 38068 31482
rect 38016 31418 38068 31424
rect 38212 31385 38240 31894
rect 38198 31376 38254 31385
rect 38198 31311 38254 31320
rect 38108 30252 38160 30258
rect 38108 30194 38160 30200
rect 38120 30025 38148 30194
rect 38292 30116 38344 30122
rect 38292 30058 38344 30064
rect 38106 30016 38162 30025
rect 38106 29951 38162 29960
rect 38016 29640 38068 29646
rect 38016 29582 38068 29588
rect 37740 29096 37792 29102
rect 37740 29038 37792 29044
rect 37752 28626 37780 29038
rect 37740 28620 37792 28626
rect 37740 28562 37792 28568
rect 38028 26042 38056 29582
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38212 29345 38240 29446
rect 38198 29336 38254 29345
rect 38198 29271 38254 29280
rect 38304 28098 38332 30058
rect 38212 28070 38332 28098
rect 38016 26036 38068 26042
rect 38016 25978 38068 25984
rect 38212 25974 38240 28070
rect 38292 27464 38344 27470
rect 38292 27406 38344 27412
rect 38304 27305 38332 27406
rect 38290 27296 38346 27305
rect 38290 27231 38346 27240
rect 38292 26988 38344 26994
rect 38292 26930 38344 26936
rect 38304 26625 38332 26930
rect 38290 26616 38346 26625
rect 38290 26551 38346 26560
rect 38200 25968 38252 25974
rect 38200 25910 38252 25916
rect 37648 25424 37700 25430
rect 37648 25366 37700 25372
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 38198 25256 38254 25265
rect 37464 24404 37516 24410
rect 37464 24346 37516 24352
rect 37740 24268 37792 24274
rect 37740 24210 37792 24216
rect 37280 21140 37332 21146
rect 37280 21082 37332 21088
rect 37648 19712 37700 19718
rect 37648 19654 37700 19660
rect 37464 19304 37516 19310
rect 37464 19246 37516 19252
rect 37476 18358 37504 19246
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37280 18148 37332 18154
rect 37280 18090 37332 18096
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 37200 16114 37228 17478
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 36634 15600 36690 15609
rect 36634 15535 36690 15544
rect 36648 12434 36676 15535
rect 37292 15473 37320 18090
rect 37278 15464 37334 15473
rect 37278 15399 37334 15408
rect 37476 14278 37504 18294
rect 37556 16720 37608 16726
rect 37556 16662 37608 16668
rect 37568 14414 37596 16662
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37464 14272 37516 14278
rect 37464 14214 37516 14220
rect 37568 13530 37596 14350
rect 37556 13524 37608 13530
rect 37556 13466 37608 13472
rect 36648 12406 36768 12434
rect 36544 11076 36596 11082
rect 36544 11018 36596 11024
rect 36452 9580 36504 9586
rect 36452 9522 36504 9528
rect 36464 9178 36492 9522
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36556 9058 36584 11018
rect 36740 10674 36768 12406
rect 37372 12232 37424 12238
rect 37372 12174 37424 12180
rect 37004 12164 37056 12170
rect 37004 12106 37056 12112
rect 36728 10668 36780 10674
rect 36728 10610 36780 10616
rect 36636 9920 36688 9926
rect 36636 9862 36688 9868
rect 36648 9722 36676 9862
rect 36636 9716 36688 9722
rect 36636 9658 36688 9664
rect 36464 9030 36584 9058
rect 36464 6769 36492 9030
rect 36544 8968 36596 8974
rect 36544 8910 36596 8916
rect 36450 6760 36506 6769
rect 36450 6695 36506 6704
rect 36452 6656 36504 6662
rect 36452 6598 36504 6604
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36464 2378 36492 6598
rect 36556 6458 36584 8910
rect 36636 7200 36688 7206
rect 36636 7142 36688 7148
rect 36648 6730 36676 7142
rect 36740 6798 36768 10610
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 36820 9580 36872 9586
rect 36820 9522 36872 9528
rect 36832 8945 36860 9522
rect 36818 8936 36874 8945
rect 36818 8871 36874 8880
rect 36820 7880 36872 7886
rect 36820 7822 36872 7828
rect 36832 7546 36860 7822
rect 36820 7540 36872 7546
rect 36820 7482 36872 7488
rect 36728 6792 36780 6798
rect 36728 6734 36780 6740
rect 36636 6724 36688 6730
rect 36636 6666 36688 6672
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 36726 5536 36782 5545
rect 36726 5471 36782 5480
rect 36634 4720 36690 4729
rect 36634 4655 36690 4664
rect 36648 3466 36676 4655
rect 36740 4622 36768 5471
rect 36820 5024 36872 5030
rect 36820 4966 36872 4972
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 36832 4185 36860 4966
rect 36818 4176 36874 4185
rect 36818 4111 36874 4120
rect 36636 3460 36688 3466
rect 36636 3402 36688 3408
rect 36924 2774 36952 9998
rect 37016 9178 37044 12106
rect 37280 11756 37332 11762
rect 37280 11698 37332 11704
rect 37096 9716 37148 9722
rect 37096 9658 37148 9664
rect 37004 9172 37056 9178
rect 37004 9114 37056 9120
rect 37004 8288 37056 8294
rect 37004 8230 37056 8236
rect 37016 7546 37044 8230
rect 37004 7540 37056 7546
rect 37004 7482 37056 7488
rect 37004 7404 37056 7410
rect 37004 7346 37056 7352
rect 36740 2746 36952 2774
rect 36452 2372 36504 2378
rect 36452 2314 36504 2320
rect 36636 2304 36688 2310
rect 36636 2246 36688 2252
rect 36648 2106 36676 2246
rect 36636 2100 36688 2106
rect 36636 2042 36688 2048
rect 36740 800 36768 2746
rect 37016 1630 37044 7346
rect 37108 4146 37136 9658
rect 37292 9194 37320 11698
rect 37384 11150 37412 12174
rect 37464 11280 37516 11286
rect 37462 11248 37464 11257
rect 37516 11248 37518 11257
rect 37462 11183 37518 11192
rect 37372 11144 37424 11150
rect 37372 11086 37424 11092
rect 37370 10976 37426 10985
rect 37370 10911 37426 10920
rect 37384 10062 37412 10911
rect 37556 10260 37608 10266
rect 37556 10202 37608 10208
rect 37372 10056 37424 10062
rect 37372 9998 37424 10004
rect 37372 9444 37424 9450
rect 37372 9386 37424 9392
rect 37200 9166 37320 9194
rect 37200 8838 37228 9166
rect 37280 9104 37332 9110
rect 37280 9046 37332 9052
rect 37188 8832 37240 8838
rect 37188 8774 37240 8780
rect 37292 5710 37320 9046
rect 37384 5710 37412 9386
rect 37464 9376 37516 9382
rect 37464 9318 37516 9324
rect 37476 6798 37504 9318
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 37464 5568 37516 5574
rect 37464 5510 37516 5516
rect 37096 4140 37148 4146
rect 37096 4082 37148 4088
rect 37476 4026 37504 5510
rect 37568 4146 37596 10202
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37476 3998 37596 4026
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37476 2514 37504 2790
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 37004 1624 37056 1630
rect 37004 1566 37056 1572
rect 33612 734 33916 762
rect 34150 200 34206 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 36726 200 36782 800
rect 37568 785 37596 3998
rect 37660 2514 37688 19654
rect 37752 3058 37780 24210
rect 38028 23866 38056 25230
rect 38198 25191 38254 25200
rect 38660 25220 38712 25226
rect 38212 25158 38240 25191
rect 38660 25162 38712 25168
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38108 24064 38160 24070
rect 38108 24006 38160 24012
rect 38016 23860 38068 23866
rect 38016 23802 38068 23808
rect 37924 23724 37976 23730
rect 37924 23666 37976 23672
rect 37936 22778 37964 23666
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 37924 22772 37976 22778
rect 37924 22714 37976 22720
rect 37936 21146 37964 22714
rect 38028 22642 38056 22918
rect 38120 22710 38148 24006
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 38108 22704 38160 22710
rect 38108 22646 38160 22652
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38016 21956 38068 21962
rect 38016 21898 38068 21904
rect 37924 21140 37976 21146
rect 37924 21082 37976 21088
rect 38028 19514 38056 21898
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38304 20505 38332 20878
rect 38290 20496 38346 20505
rect 38290 20431 38346 20440
rect 38106 19816 38162 19825
rect 38106 19751 38108 19760
rect 38160 19751 38162 19760
rect 38108 19722 38160 19728
rect 38016 19508 38068 19514
rect 38016 19450 38068 19456
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 38304 19145 38332 19314
rect 38290 19136 38346 19145
rect 38290 19071 38346 19080
rect 38568 18828 38620 18834
rect 38568 18770 38620 18776
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 37924 18080 37976 18086
rect 37924 18022 37976 18028
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 37844 8974 37872 14758
rect 37936 14414 37964 18022
rect 38120 17785 38148 18226
rect 38106 17776 38162 17785
rect 38106 17711 38162 17720
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 38304 17105 38332 17138
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 38120 16658 38148 16934
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 38016 15496 38068 15502
rect 38016 15438 38068 15444
rect 38028 14618 38056 15438
rect 38120 15026 38148 16594
rect 38474 16416 38530 16425
rect 38474 16351 38530 16360
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38212 15065 38240 15302
rect 38198 15056 38254 15065
rect 38108 15020 38160 15026
rect 38198 14991 38254 15000
rect 38108 14962 38160 14968
rect 38016 14612 38068 14618
rect 38016 14554 38068 14560
rect 37924 14408 37976 14414
rect 37924 14350 37976 14356
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 37936 10266 37964 14214
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38304 13025 38332 13262
rect 38290 13016 38346 13025
rect 38290 12951 38346 12960
rect 38108 12844 38160 12850
rect 38108 12786 38160 12792
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 37924 10260 37976 10266
rect 37924 10202 37976 10208
rect 38028 10146 38056 12582
rect 38120 12345 38148 12786
rect 38198 12744 38254 12753
rect 38198 12679 38254 12688
rect 38212 12646 38240 12679
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38106 12336 38162 12345
rect 38106 12271 38162 12280
rect 38108 11552 38160 11558
rect 38108 11494 38160 11500
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38120 11218 38148 11494
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 38120 10985 38148 11018
rect 38106 10976 38162 10985
rect 38106 10911 38162 10920
rect 38108 10668 38160 10674
rect 38108 10610 38160 10616
rect 38120 10305 38148 10610
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 37936 10118 38056 10146
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37844 7698 37872 8774
rect 37936 7886 37964 10118
rect 38108 9920 38160 9926
rect 38108 9862 38160 9868
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 38028 8498 38056 9318
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 37924 7880 37976 7886
rect 37924 7822 37976 7828
rect 38120 7818 38148 9862
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38200 8356 38252 8362
rect 38200 8298 38252 8304
rect 38212 8265 38240 8298
rect 38198 8256 38254 8265
rect 38198 8191 38254 8200
rect 38108 7812 38160 7818
rect 38108 7754 38160 7760
rect 37844 7670 37964 7698
rect 37936 7410 37964 7670
rect 37924 7404 37976 7410
rect 37924 7346 37976 7352
rect 38120 7290 38148 7754
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38212 7585 38240 7686
rect 38198 7576 38254 7585
rect 38198 7511 38254 7520
rect 38304 7410 38332 11494
rect 38384 10056 38436 10062
rect 38384 9998 38436 10004
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 37936 7262 38148 7290
rect 37936 3534 37964 7262
rect 38108 7200 38160 7206
rect 38108 7142 38160 7148
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 38028 800 38056 5510
rect 38120 5234 38148 7142
rect 38292 6656 38344 6662
rect 38292 6598 38344 6604
rect 38198 6216 38254 6225
rect 38198 6151 38254 6160
rect 38212 6118 38240 6151
rect 38200 6112 38252 6118
rect 38200 6054 38252 6060
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 38200 3732 38252 3738
rect 38200 3674 38252 3680
rect 38212 3641 38240 3674
rect 38198 3632 38254 3641
rect 38198 3567 38254 3576
rect 38304 3505 38332 6598
rect 38396 5545 38424 9998
rect 38382 5536 38438 5545
rect 38382 5471 38438 5480
rect 38488 3602 38516 16351
rect 38580 5166 38608 18770
rect 38672 11286 38700 25162
rect 38752 19916 38804 19922
rect 38752 19858 38804 19864
rect 38660 11280 38712 11286
rect 38660 11222 38712 11228
rect 38660 11144 38712 11150
rect 38660 11086 38712 11092
rect 38568 5160 38620 5166
rect 38568 5102 38620 5108
rect 38672 4554 38700 11086
rect 38764 10742 38792 19858
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38752 10736 38804 10742
rect 38752 10678 38804 10684
rect 38856 4622 38884 18702
rect 39028 12096 39080 12102
rect 39028 12038 39080 12044
rect 38936 11620 38988 11626
rect 38936 11562 38988 11568
rect 38844 4616 38896 4622
rect 38844 4558 38896 4564
rect 38660 4548 38712 4554
rect 38660 4490 38712 4496
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 38476 3596 38528 3602
rect 38476 3538 38528 3544
rect 38290 3496 38346 3505
rect 38290 3431 38346 3440
rect 38672 800 38700 4014
rect 38948 3369 38976 11562
rect 38934 3360 38990 3369
rect 38934 3295 38990 3304
rect 39040 1834 39068 12038
rect 39304 4684 39356 4690
rect 39304 4626 39356 4632
rect 39028 1828 39080 1834
rect 39028 1770 39080 1776
rect 39316 800 39344 4626
rect 37554 776 37610 785
rect 37554 711 37610 720
rect 38014 200 38070 800
rect 38658 200 38714 800
rect 39302 200 39358 800
<< via2 >>
rect 2870 38800 2926 38856
rect 3146 38120 3202 38176
rect 1582 36760 1638 36816
rect 1674 36116 1676 36136
rect 1676 36116 1728 36136
rect 1728 36116 1730 36136
rect 1674 36080 1730 36116
rect 1766 35436 1768 35456
rect 1768 35436 1820 35456
rect 1820 35436 1822 35456
rect 1766 35400 1822 35436
rect 1766 34040 1822 34096
rect 1766 33380 1822 33416
rect 1766 33360 1768 33380
rect 1768 33360 1820 33380
rect 1820 33360 1822 33380
rect 1582 32000 1638 32056
rect 846 26968 902 27024
rect 1766 31320 1822 31376
rect 1766 30676 1768 30696
rect 1768 30676 1820 30696
rect 1820 30676 1822 30696
rect 1766 30640 1822 30676
rect 1766 29280 1822 29336
rect 1766 28600 1822 28656
rect 1766 27276 1768 27296
rect 1768 27276 1820 27296
rect 1820 27276 1822 27296
rect 1766 27240 1822 27276
rect 1766 26560 1822 26616
rect 1766 25200 1822 25256
rect 1766 24520 1822 24576
rect 1766 23840 1822 23896
rect 1766 22480 1822 22536
rect 1766 21836 1768 21856
rect 1768 21836 1820 21856
rect 1820 21836 1822 21856
rect 1766 21800 1822 21836
rect 1766 20440 1822 20496
rect 1582 19796 1584 19816
rect 1584 19796 1636 19816
rect 1636 19796 1638 19816
rect 1582 19760 1638 19796
rect 1766 19116 1768 19136
rect 1768 19116 1820 19136
rect 1820 19116 1822 19136
rect 1766 19080 1822 19116
rect 1766 17720 1822 17776
rect 1582 17076 1584 17096
rect 1584 17076 1636 17096
rect 1636 17076 1638 17096
rect 1582 17040 1638 17076
rect 1766 15680 1822 15736
rect 1674 15000 1730 15056
rect 1766 14320 1822 14376
rect 1858 13776 1914 13832
rect 1582 12960 1638 13016
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 2594 23432 2650 23488
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 2318 18536 2374 18592
rect 1398 8200 1454 8256
rect 1674 12280 1730 12336
rect 1766 10956 1768 10976
rect 1768 10956 1820 10976
rect 1820 10956 1822 10976
rect 1766 10920 1822 10956
rect 1766 10240 1822 10296
rect 1766 9560 1822 9616
rect 1766 7520 1822 7576
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 1858 5888 1914 5944
rect 1674 5480 1730 5536
rect 2226 7112 2282 7168
rect 1766 3440 1822 3496
rect 1674 2760 1730 2816
rect 1490 1400 1546 1456
rect 1950 3576 2006 3632
rect 2134 5480 2190 5536
rect 2226 3440 2282 3496
rect 2318 2624 2374 2680
rect 2594 6740 2596 6760
rect 2596 6740 2648 6760
rect 2648 6740 2650 6760
rect 2594 6704 2650 6740
rect 3054 8744 3110 8800
rect 2870 4800 2926 4856
rect 3330 7928 3386 7984
rect 3054 4664 3110 4720
rect 3514 7384 3570 7440
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4986 15544 5042 15600
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4066 12416 4122 12472
rect 3882 12280 3938 12336
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 5078 13640 5134 13696
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4066 10104 4122 10160
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4250 8608 4306 8664
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4710 8744 4766 8800
rect 4618 7520 4674 7576
rect 4986 8200 5042 8256
rect 3606 4120 3662 4176
rect 4526 7248 4582 7304
rect 3882 6568 3938 6624
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4250 6316 4306 6352
rect 4250 6296 4252 6316
rect 4252 6296 4304 6316
rect 4304 6296 4306 6316
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4250 5752 4306 5808
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4526 4256 4582 4312
rect 3974 4020 3976 4040
rect 3976 4020 4028 4040
rect 4028 4020 4030 4040
rect 3974 3984 4030 4020
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3974 3168 4030 3224
rect 5078 6996 5134 7032
rect 5078 6976 5080 6996
rect 5080 6976 5132 6996
rect 5132 6976 5134 6996
rect 5078 6840 5134 6896
rect 4802 2896 4858 2952
rect 5354 11464 5410 11520
rect 5538 9424 5594 9480
rect 5538 9016 5594 9072
rect 5354 8084 5410 8120
rect 5354 8064 5356 8084
rect 5356 8064 5408 8084
rect 5408 8064 5410 8084
rect 5354 7828 5356 7848
rect 5356 7828 5408 7848
rect 5408 7828 5410 7848
rect 5354 7792 5410 7828
rect 6550 18708 6552 18728
rect 6552 18708 6604 18728
rect 6604 18708 6606 18728
rect 6550 18672 6606 18708
rect 6182 11600 6238 11656
rect 5906 10784 5962 10840
rect 5814 10004 5816 10024
rect 5816 10004 5868 10024
rect 5868 10004 5870 10024
rect 5814 9968 5870 10004
rect 5906 9596 5908 9616
rect 5908 9596 5960 9616
rect 5960 9596 5962 9616
rect 5906 9560 5962 9596
rect 5078 3304 5134 3360
rect 4986 2896 5042 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4158 2488 4214 2544
rect 5630 5092 5686 5128
rect 5630 5072 5632 5092
rect 5632 5072 5684 5092
rect 5684 5072 5686 5092
rect 5722 4936 5778 4992
rect 6366 10920 6422 10976
rect 6274 9832 6330 9888
rect 6182 9152 6238 9208
rect 6090 8336 6146 8392
rect 6458 9696 6514 9752
rect 6366 9560 6422 9616
rect 6642 11056 6698 11112
rect 8482 27240 8538 27296
rect 6734 9968 6790 10024
rect 6918 10648 6974 10704
rect 6734 9152 6790 9208
rect 6366 8492 6422 8528
rect 6366 8472 6368 8492
rect 6368 8472 6420 8492
rect 6420 8472 6422 8492
rect 6274 7112 6330 7168
rect 5998 2896 6054 2952
rect 6366 5636 6422 5672
rect 6366 5616 6368 5636
rect 6368 5616 6420 5636
rect 6420 5616 6422 5636
rect 6366 3984 6422 4040
rect 7194 11756 7250 11792
rect 7194 11736 7196 11756
rect 7196 11736 7248 11756
rect 7248 11736 7250 11756
rect 7010 7656 7066 7712
rect 6826 6180 6882 6216
rect 6826 6160 6828 6180
rect 6828 6160 6880 6180
rect 6880 6160 6882 6180
rect 7010 5480 7066 5536
rect 7010 5208 7066 5264
rect 6642 4256 6698 4312
rect 8022 15136 8078 15192
rect 7930 11328 7986 11384
rect 7746 10920 7802 10976
rect 7470 10104 7526 10160
rect 7378 8472 7434 8528
rect 7378 6024 7434 6080
rect 7654 9988 7710 10024
rect 7654 9968 7656 9988
rect 7656 9968 7708 9988
rect 7708 9968 7710 9988
rect 7930 9560 7986 9616
rect 7746 8200 7802 8256
rect 7930 8336 7986 8392
rect 7838 8064 7894 8120
rect 7838 7792 7894 7848
rect 7838 6976 7894 7032
rect 7838 6840 7894 6896
rect 7562 5480 7618 5536
rect 7562 3460 7618 3496
rect 7562 3440 7564 3460
rect 7564 3440 7616 3460
rect 7616 3440 7618 3460
rect 7194 2760 7250 2816
rect 7746 6432 7802 6488
rect 7838 4936 7894 4992
rect 7838 3304 7894 3360
rect 7654 2760 7710 2816
rect 8482 11872 8538 11928
rect 8206 10648 8262 10704
rect 8390 9832 8446 9888
rect 8022 7384 8078 7440
rect 8206 6840 8262 6896
rect 8390 9424 8446 9480
rect 8390 9152 8446 9208
rect 8574 7656 8630 7712
rect 8298 5772 8354 5808
rect 8298 5752 8300 5772
rect 8300 5752 8352 5772
rect 8352 5752 8354 5772
rect 8114 5072 8170 5128
rect 8850 13912 8906 13968
rect 9494 17992 9550 18048
rect 9126 13268 9128 13288
rect 9128 13268 9180 13288
rect 9180 13268 9182 13288
rect 9126 13232 9182 13268
rect 9678 16632 9734 16688
rect 9770 14900 9772 14920
rect 9772 14900 9824 14920
rect 9824 14900 9826 14920
rect 9770 14864 9826 14900
rect 10322 21664 10378 21720
rect 11242 26424 11298 26480
rect 10598 17620 10600 17640
rect 10600 17620 10652 17640
rect 10652 17620 10654 17640
rect 10598 17584 10654 17620
rect 10230 16360 10286 16416
rect 10138 15988 10140 16008
rect 10140 15988 10192 16008
rect 10192 15988 10194 16008
rect 10138 15952 10194 15988
rect 9954 15000 10010 15056
rect 9126 12844 9182 12880
rect 9126 12824 9128 12844
rect 9128 12824 9180 12844
rect 9180 12824 9182 12844
rect 8850 7520 8906 7576
rect 8758 6840 8814 6896
rect 8758 6024 8814 6080
rect 8666 3440 8722 3496
rect 9310 11872 9366 11928
rect 9678 12300 9734 12336
rect 9678 12280 9680 12300
rect 9680 12280 9732 12300
rect 9732 12280 9734 12300
rect 9678 12144 9734 12200
rect 9494 11736 9550 11792
rect 9678 10648 9734 10704
rect 9310 8336 9366 8392
rect 9310 6860 9366 6896
rect 9310 6840 9312 6860
rect 9312 6840 9364 6860
rect 9364 6840 9366 6860
rect 9494 6452 9550 6488
rect 9494 6432 9496 6452
rect 9496 6432 9548 6452
rect 9548 6432 9550 6452
rect 9126 5244 9128 5264
rect 9128 5244 9180 5264
rect 9180 5244 9182 5264
rect 8942 4140 8998 4176
rect 8942 4120 8944 4140
rect 8944 4120 8996 4140
rect 8996 4120 8998 4140
rect 9126 5208 9182 5244
rect 9402 5108 9404 5128
rect 9404 5108 9456 5128
rect 9456 5108 9458 5128
rect 9402 5072 9458 5108
rect 9402 3188 9458 3224
rect 9402 3168 9404 3188
rect 9404 3168 9456 3188
rect 9456 3168 9458 3188
rect 9770 10376 9826 10432
rect 10230 12280 10286 12336
rect 10138 11620 10194 11656
rect 10138 11600 10140 11620
rect 10140 11600 10192 11620
rect 10192 11600 10194 11620
rect 10046 11056 10102 11112
rect 9862 9696 9918 9752
rect 9862 8608 9918 8664
rect 9678 7112 9734 7168
rect 10230 10920 10286 10976
rect 10230 8880 10286 8936
rect 9954 8200 10010 8256
rect 9770 5772 9826 5808
rect 9770 5752 9772 5772
rect 9772 5752 9824 5772
rect 9824 5752 9826 5772
rect 10506 12416 10562 12472
rect 10598 11600 10654 11656
rect 10506 10512 10562 10568
rect 10506 9560 10562 9616
rect 10598 9288 10654 9344
rect 10598 6724 10654 6760
rect 10598 6704 10600 6724
rect 10600 6704 10652 6724
rect 10652 6704 10654 6724
rect 10690 6296 10746 6352
rect 11058 13368 11114 13424
rect 11058 12008 11114 12064
rect 11058 11328 11114 11384
rect 10966 8880 11022 8936
rect 10874 8744 10930 8800
rect 11702 24792 11758 24848
rect 12806 26424 12862 26480
rect 11702 21392 11758 21448
rect 12346 19916 12402 19952
rect 12346 19896 12348 19916
rect 12348 19896 12400 19916
rect 12400 19896 12402 19916
rect 11426 16088 11482 16144
rect 11334 15408 11390 15464
rect 11794 16496 11850 16552
rect 11518 12552 11574 12608
rect 11334 10784 11390 10840
rect 11150 8472 11206 8528
rect 11334 6432 11390 6488
rect 11702 12688 11758 12744
rect 11702 12280 11758 12336
rect 11702 11872 11758 11928
rect 11978 12164 12034 12200
rect 11978 12144 11980 12164
rect 11980 12144 12032 12164
rect 12032 12144 12034 12164
rect 11978 9988 12034 10024
rect 11978 9968 11980 9988
rect 11980 9968 12032 9988
rect 12032 9968 12034 9988
rect 11518 8744 11574 8800
rect 11426 5616 11482 5672
rect 10966 4392 11022 4448
rect 10782 4020 10784 4040
rect 10784 4020 10836 4040
rect 10836 4020 10838 4040
rect 10782 3984 10838 4020
rect 10782 2896 10838 2952
rect 10966 2760 11022 2816
rect 11610 7112 11666 7168
rect 11886 6996 11942 7032
rect 11886 6976 11888 6996
rect 11888 6976 11940 6996
rect 11940 6976 11942 6996
rect 12530 21548 12586 21584
rect 12530 21528 12532 21548
rect 12532 21528 12584 21548
rect 12584 21528 12586 21548
rect 12898 26016 12954 26072
rect 13082 25744 13138 25800
rect 13726 22616 13782 22672
rect 13358 21528 13414 21584
rect 13358 20712 13414 20768
rect 12714 19896 12770 19952
rect 12806 18128 12862 18184
rect 12438 12824 12494 12880
rect 12622 11636 12624 11656
rect 12624 11636 12676 11656
rect 12676 11636 12678 11656
rect 12622 11600 12678 11636
rect 12622 10684 12624 10704
rect 12624 10684 12676 10704
rect 12676 10684 12678 10704
rect 12622 10648 12678 10684
rect 12438 9832 12494 9888
rect 12438 8628 12494 8664
rect 12438 8608 12440 8628
rect 12440 8608 12492 8628
rect 12492 8608 12494 8628
rect 12438 6996 12494 7032
rect 12438 6976 12440 6996
rect 12440 6976 12492 6996
rect 12492 6976 12494 6996
rect 12622 6840 12678 6896
rect 13266 17856 13322 17912
rect 12990 16108 13046 16144
rect 12990 16088 12992 16108
rect 12992 16088 13044 16108
rect 13044 16088 13046 16108
rect 12898 14864 12954 14920
rect 12898 14456 12954 14512
rect 12898 14184 12954 14240
rect 13634 20848 13690 20904
rect 13634 19488 13690 19544
rect 13634 16496 13690 16552
rect 13266 14184 13322 14240
rect 12898 12552 12954 12608
rect 13082 12824 13138 12880
rect 13634 13504 13690 13560
rect 13358 12280 13414 12336
rect 13450 10648 13506 10704
rect 13174 8780 13176 8800
rect 13176 8780 13228 8800
rect 13228 8780 13230 8800
rect 13174 8744 13230 8780
rect 13082 6840 13138 6896
rect 13634 12300 13690 12336
rect 13634 12280 13636 12300
rect 13636 12280 13688 12300
rect 13688 12280 13690 12300
rect 13910 11328 13966 11384
rect 14554 25336 14610 25392
rect 14370 17040 14426 17096
rect 14462 16632 14518 16688
rect 14094 11192 14150 11248
rect 14462 14456 14518 14512
rect 13818 10512 13874 10568
rect 14002 10376 14058 10432
rect 13542 6976 13598 7032
rect 13818 7112 13874 7168
rect 13726 5344 13782 5400
rect 13726 4800 13782 4856
rect 14094 9832 14150 9888
rect 14002 4936 14058 4992
rect 13910 4528 13966 4584
rect 14094 4120 14150 4176
rect 15014 24404 15070 24440
rect 15014 24384 15016 24404
rect 15016 24384 15068 24404
rect 15068 24384 15070 24404
rect 15842 26988 15898 27024
rect 15842 26968 15844 26988
rect 15844 26968 15896 26988
rect 15896 26968 15898 26988
rect 15474 19780 15530 19816
rect 15474 19760 15476 19780
rect 15476 19760 15528 19780
rect 15528 19760 15530 19780
rect 15290 16632 15346 16688
rect 15382 16360 15438 16416
rect 14830 13232 14886 13288
rect 14830 12416 14886 12472
rect 14738 11872 14794 11928
rect 14554 8744 14610 8800
rect 14830 10920 14886 10976
rect 14830 9288 14886 9344
rect 14738 7248 14794 7304
rect 14646 4256 14702 4312
rect 18234 29688 18290 29744
rect 16486 23024 16542 23080
rect 16394 21684 16450 21720
rect 16394 21664 16396 21684
rect 16396 21664 16448 21684
rect 16448 21664 16450 21684
rect 15658 16904 15714 16960
rect 15106 5344 15162 5400
rect 15106 4936 15162 4992
rect 15106 4256 15162 4312
rect 15566 13232 15622 13288
rect 15290 8336 15346 8392
rect 15474 11348 15530 11384
rect 15474 11328 15476 11348
rect 15476 11328 15528 11348
rect 15528 11328 15530 11348
rect 15474 11212 15530 11248
rect 15474 11192 15476 11212
rect 15476 11192 15528 11212
rect 15528 11192 15530 11212
rect 15842 19932 15844 19952
rect 15844 19932 15896 19952
rect 15896 19932 15898 19952
rect 15842 19896 15898 19932
rect 15842 16632 15898 16688
rect 15842 9152 15898 9208
rect 15750 8744 15806 8800
rect 15934 8608 15990 8664
rect 16210 15308 16212 15328
rect 16212 15308 16264 15328
rect 16264 15308 16266 15328
rect 16210 15272 16266 15308
rect 16486 17876 16542 17912
rect 16486 17856 16488 17876
rect 16488 17856 16540 17876
rect 16540 17856 16542 17876
rect 16302 13640 16358 13696
rect 16118 9424 16174 9480
rect 16026 7248 16082 7304
rect 16394 12824 16450 12880
rect 16486 11872 16542 11928
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 17682 26036 17738 26072
rect 17682 26016 17684 26036
rect 17684 26016 17736 26036
rect 17736 26016 17738 26036
rect 17314 24384 17370 24440
rect 17682 20868 17738 20904
rect 17682 20848 17684 20868
rect 17684 20848 17736 20868
rect 17736 20848 17738 20868
rect 18510 24928 18566 24984
rect 18418 24656 18474 24712
rect 18418 23432 18474 23488
rect 17314 19352 17370 19408
rect 16854 15952 16910 16008
rect 17038 14728 17094 14784
rect 16946 13640 17002 13696
rect 17406 13640 17462 13696
rect 16762 11192 16818 11248
rect 16946 11056 17002 11112
rect 16670 9968 16726 10024
rect 16946 8880 17002 8936
rect 16302 8064 16358 8120
rect 16118 5480 16174 5536
rect 16578 5752 16634 5808
rect 16302 5344 16358 5400
rect 16026 3304 16082 3360
rect 16302 4020 16304 4040
rect 16304 4020 16356 4040
rect 16356 4020 16358 4040
rect 16302 3984 16358 4020
rect 17130 12008 17186 12064
rect 17130 8900 17186 8936
rect 17130 8880 17132 8900
rect 17132 8880 17184 8900
rect 17184 8880 17186 8900
rect 16946 7384 17002 7440
rect 17406 9016 17462 9072
rect 18050 19488 18106 19544
rect 17590 9968 17646 10024
rect 17406 7540 17462 7576
rect 17406 7520 17408 7540
rect 17408 7520 17460 7540
rect 17460 7520 17462 7540
rect 17590 6976 17646 7032
rect 17406 6840 17462 6896
rect 18326 18164 18328 18184
rect 18328 18164 18380 18184
rect 18380 18164 18382 18184
rect 18326 18128 18382 18164
rect 18786 26424 18842 26480
rect 18970 25880 19026 25936
rect 18694 16768 18750 16824
rect 18602 16652 18658 16688
rect 18602 16632 18604 16652
rect 18604 16632 18656 16652
rect 18656 16632 18658 16652
rect 18418 15272 18474 15328
rect 19154 25744 19210 25800
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19614 24520 19670 24576
rect 19890 24384 19946 24440
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19890 23160 19946 23216
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20166 26460 20168 26480
rect 20168 26460 20220 26480
rect 20220 26460 20222 26480
rect 20166 26424 20222 26460
rect 19522 22208 19578 22264
rect 19338 21936 19394 21992
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20074 22072 20130 22128
rect 19062 20440 19118 20496
rect 18142 11192 18198 11248
rect 18050 9696 18106 9752
rect 17866 8064 17922 8120
rect 17682 5752 17738 5808
rect 18878 15272 18934 15328
rect 19062 15000 19118 15056
rect 18786 13232 18842 13288
rect 18234 8200 18290 8256
rect 18602 9696 18658 9752
rect 18418 9424 18474 9480
rect 18510 8916 18512 8936
rect 18512 8916 18564 8936
rect 18564 8916 18566 8936
rect 18510 8880 18566 8916
rect 18234 6160 18290 6216
rect 17314 4936 17370 4992
rect 17590 4936 17646 4992
rect 17406 4548 17462 4584
rect 17406 4528 17408 4548
rect 17408 4528 17460 4548
rect 17460 4528 17462 4548
rect 17498 3884 17500 3904
rect 17500 3884 17552 3904
rect 17552 3884 17554 3904
rect 17498 3848 17554 3884
rect 16670 2644 16726 2680
rect 16670 2624 16672 2644
rect 16672 2624 16724 2644
rect 16724 2624 16726 2644
rect 18510 7520 18566 7576
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20258 25236 20260 25256
rect 20260 25236 20312 25256
rect 20312 25236 20314 25256
rect 20258 25200 20314 25236
rect 20626 25336 20682 25392
rect 20442 24248 20498 24304
rect 20442 23840 20498 23896
rect 20350 23296 20406 23352
rect 20258 22072 20314 22128
rect 20166 21936 20222 21992
rect 20258 20848 20314 20904
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19890 18300 19892 18320
rect 19892 18300 19944 18320
rect 19944 18300 19946 18320
rect 19890 18264 19946 18300
rect 19430 18028 19432 18048
rect 19432 18028 19484 18048
rect 19484 18028 19486 18048
rect 19430 17992 19486 18028
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19430 16088 19486 16144
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19430 14728 19486 14784
rect 20166 18264 20222 18320
rect 20718 23432 20774 23488
rect 20534 20848 20590 20904
rect 20258 16496 20314 16552
rect 20258 16088 20314 16144
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19338 13948 19340 13968
rect 19340 13948 19392 13968
rect 19392 13948 19394 13968
rect 19338 13912 19394 13948
rect 19154 12708 19210 12744
rect 19154 12688 19156 12708
rect 19156 12688 19208 12708
rect 19208 12688 19210 12708
rect 19338 12688 19394 12744
rect 19614 13776 19670 13832
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19430 12436 19486 12472
rect 19430 12416 19432 12436
rect 19432 12416 19484 12436
rect 19484 12416 19486 12436
rect 20350 15680 20406 15736
rect 20074 12552 20130 12608
rect 20074 12416 20130 12472
rect 19890 12280 19946 12336
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19246 9460 19248 9480
rect 19248 9460 19300 9480
rect 19300 9460 19302 9480
rect 19246 9424 19302 9460
rect 19890 9424 19946 9480
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19154 8336 19210 8392
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 18970 7112 19026 7168
rect 18878 6976 18934 7032
rect 19154 6432 19210 6488
rect 18878 4528 18934 4584
rect 19062 3304 19118 3360
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20350 12552 20406 12608
rect 20534 16904 20590 16960
rect 21178 27784 21234 27840
rect 20902 21392 20958 21448
rect 20994 21120 21050 21176
rect 20902 20304 20958 20360
rect 20994 19896 21050 19952
rect 20718 18128 20774 18184
rect 20902 15680 20958 15736
rect 20626 14048 20682 14104
rect 20718 13948 20720 13968
rect 20720 13948 20772 13968
rect 20772 13948 20774 13968
rect 20718 13912 20774 13948
rect 20810 13776 20866 13832
rect 20718 13524 20774 13560
rect 20718 13504 20720 13524
rect 20720 13504 20772 13524
rect 20772 13504 20774 13524
rect 21086 15680 21142 15736
rect 21086 15408 21142 15464
rect 20994 13640 21050 13696
rect 20902 13232 20958 13288
rect 20534 13132 20536 13152
rect 20536 13132 20588 13152
rect 20588 13132 20590 13152
rect 20534 13096 20590 13132
rect 20718 13096 20774 13152
rect 20534 12688 20590 12744
rect 20442 12416 20498 12472
rect 20258 12144 20314 12200
rect 20534 12144 20590 12200
rect 20442 10920 20498 10976
rect 20350 10648 20406 10704
rect 20166 7404 20222 7440
rect 20166 7384 20168 7404
rect 20168 7384 20220 7404
rect 20220 7384 20222 7404
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20442 9832 20498 9888
rect 20626 11600 20682 11656
rect 20718 10648 20774 10704
rect 20534 6976 20590 7032
rect 20442 6840 20498 6896
rect 20258 6432 20314 6488
rect 19430 4392 19486 4448
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 21546 20984 21602 21040
rect 21454 17876 21510 17912
rect 21454 17856 21456 17876
rect 21456 17856 21508 17876
rect 21508 17856 21510 17876
rect 20994 11192 21050 11248
rect 20994 9596 20996 9616
rect 20996 9596 21048 9616
rect 21048 9596 21050 9616
rect 20994 9560 21050 9596
rect 21178 8064 21234 8120
rect 21178 7792 21234 7848
rect 21086 7248 21142 7304
rect 22374 27920 22430 27976
rect 22190 27648 22246 27704
rect 22006 20712 22062 20768
rect 22282 21664 22338 21720
rect 22374 19780 22430 19816
rect 22374 19760 22376 19780
rect 22376 19760 22428 19780
rect 22428 19760 22430 19780
rect 22098 19388 22100 19408
rect 22100 19388 22152 19408
rect 22152 19388 22154 19408
rect 22098 19352 22154 19388
rect 21638 12416 21694 12472
rect 21546 12280 21602 12336
rect 21454 10648 21510 10704
rect 22558 21392 22614 21448
rect 22374 12552 22430 12608
rect 22742 21972 22744 21992
rect 22744 21972 22796 21992
rect 22796 21972 22798 21992
rect 22742 21936 22798 21972
rect 23478 26832 23534 26888
rect 23202 23704 23258 23760
rect 23202 23604 23204 23624
rect 23204 23604 23256 23624
rect 23256 23604 23258 23624
rect 23202 23568 23258 23604
rect 22834 21120 22890 21176
rect 23018 19624 23074 19680
rect 23294 21120 23350 21176
rect 24858 30096 24914 30152
rect 24122 27376 24178 27432
rect 24214 26288 24270 26344
rect 23846 23568 23902 23624
rect 24214 23724 24270 23760
rect 24214 23704 24216 23724
rect 24216 23704 24268 23724
rect 24268 23704 24270 23724
rect 23570 21564 23572 21584
rect 23572 21564 23624 21584
rect 23624 21564 23626 21584
rect 23570 21528 23626 21564
rect 23478 20848 23534 20904
rect 22742 16904 22798 16960
rect 22558 11736 22614 11792
rect 23018 18028 23020 18048
rect 23020 18028 23072 18048
rect 23072 18028 23074 18048
rect 23018 17992 23074 18028
rect 23110 15816 23166 15872
rect 21454 6296 21510 6352
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21454 4120 21510 4176
rect 21270 3168 21326 3224
rect 1858 720 1914 776
rect 21822 6024 21878 6080
rect 21730 3712 21786 3768
rect 21822 3188 21878 3224
rect 22282 8200 22338 8256
rect 22190 7656 22246 7712
rect 22834 9424 22890 9480
rect 22742 8336 22798 8392
rect 22282 6060 22284 6080
rect 22284 6060 22336 6080
rect 22336 6060 22338 6080
rect 22282 6024 22338 6060
rect 21822 3168 21824 3188
rect 21824 3168 21876 3188
rect 21876 3168 21878 3188
rect 22282 5480 22338 5536
rect 22374 4936 22430 4992
rect 22742 6840 22798 6896
rect 22650 5908 22706 5944
rect 22650 5888 22652 5908
rect 22652 5888 22704 5908
rect 22704 5888 22706 5908
rect 23110 8608 23166 8664
rect 23202 6432 23258 6488
rect 22466 3304 22522 3360
rect 23386 7384 23442 7440
rect 23938 20884 23940 20904
rect 23940 20884 23992 20904
rect 23992 20884 23994 20904
rect 23938 20848 23994 20884
rect 24582 24928 24638 24984
rect 24950 26460 24952 26480
rect 24952 26460 25004 26480
rect 25004 26460 25006 26480
rect 24950 26424 25006 26460
rect 24122 16244 24178 16280
rect 24122 16224 24124 16244
rect 24124 16224 24176 16244
rect 24176 16224 24178 16244
rect 24030 15544 24086 15600
rect 23938 12416 23994 12472
rect 24214 14864 24270 14920
rect 24950 23840 25006 23896
rect 25134 25880 25190 25936
rect 25410 27784 25466 27840
rect 25410 24656 25466 24712
rect 25318 24384 25374 24440
rect 24950 20712 25006 20768
rect 25870 27920 25926 27976
rect 25778 27784 25834 27840
rect 24858 17176 24914 17232
rect 25778 21528 25834 21584
rect 25686 20984 25742 21040
rect 26238 24520 26294 24576
rect 25962 21428 25964 21448
rect 25964 21428 26016 21448
rect 26016 21428 26018 21448
rect 25962 21392 26018 21428
rect 25870 20168 25926 20224
rect 25686 18672 25742 18728
rect 24858 15564 24914 15600
rect 24858 15544 24860 15564
rect 24860 15544 24912 15564
rect 24912 15544 24914 15564
rect 24674 15272 24730 15328
rect 24122 8472 24178 8528
rect 24306 6604 24308 6624
rect 24308 6604 24360 6624
rect 24360 6604 24362 6624
rect 24306 6568 24362 6604
rect 24582 12144 24638 12200
rect 24582 10512 24638 10568
rect 24766 9424 24822 9480
rect 24674 9016 24730 9072
rect 24582 5752 24638 5808
rect 24398 4936 24454 4992
rect 24214 3848 24270 3904
rect 24582 3984 24638 4040
rect 24490 3712 24546 3768
rect 24766 6976 24822 7032
rect 25502 17312 25558 17368
rect 25686 16632 25742 16688
rect 25318 12280 25374 12336
rect 25502 11056 25558 11112
rect 26146 19080 26202 19136
rect 26330 18808 26386 18864
rect 26422 17992 26478 18048
rect 26698 22888 26754 22944
rect 27158 27920 27214 27976
rect 27158 26852 27214 26888
rect 27158 26832 27160 26852
rect 27160 26832 27212 26852
rect 27212 26832 27214 26852
rect 26974 24792 27030 24848
rect 26882 23160 26938 23216
rect 27066 20460 27122 20496
rect 27066 20440 27068 20460
rect 27068 20440 27120 20460
rect 27120 20440 27122 20460
rect 26790 19216 26846 19272
rect 26790 19080 26846 19136
rect 26698 18692 26754 18728
rect 26698 18672 26700 18692
rect 26700 18672 26752 18692
rect 26752 18672 26754 18692
rect 26698 17992 26754 18048
rect 25962 12280 26018 12336
rect 25594 6840 25650 6896
rect 26054 10532 26110 10568
rect 26054 10512 26056 10532
rect 26056 10512 26108 10532
rect 26108 10512 26110 10532
rect 26054 9696 26110 9752
rect 25226 3168 25282 3224
rect 26146 7812 26202 7848
rect 26146 7792 26148 7812
rect 26148 7792 26200 7812
rect 26200 7792 26202 7812
rect 27434 24928 27490 24984
rect 27526 23432 27582 23488
rect 27710 22888 27766 22944
rect 27250 21936 27306 21992
rect 27434 21292 27436 21312
rect 27436 21292 27488 21312
rect 27488 21292 27490 21312
rect 27434 21256 27490 21292
rect 27710 21256 27766 21312
rect 27342 19624 27398 19680
rect 27066 19488 27122 19544
rect 26606 11328 26662 11384
rect 26790 9832 26846 9888
rect 26698 7656 26754 7712
rect 26698 7520 26754 7576
rect 26330 6996 26386 7032
rect 26330 6976 26332 6996
rect 26332 6976 26384 6996
rect 26384 6976 26386 6996
rect 26606 7112 26662 7168
rect 27250 17856 27306 17912
rect 28170 27376 28226 27432
rect 28538 26324 28540 26344
rect 28540 26324 28592 26344
rect 28592 26324 28594 26344
rect 28538 26288 28594 26324
rect 27986 19896 28042 19952
rect 27894 19780 27950 19816
rect 27894 19760 27896 19780
rect 27896 19760 27948 19780
rect 27948 19760 27950 19780
rect 27986 18944 28042 19000
rect 27986 18400 28042 18456
rect 27526 15680 27582 15736
rect 26882 8780 26884 8800
rect 26884 8780 26936 8800
rect 26936 8780 26938 8800
rect 26882 8744 26938 8780
rect 27066 8064 27122 8120
rect 26790 6840 26846 6896
rect 27342 14340 27398 14376
rect 27342 14320 27344 14340
rect 27344 14320 27396 14340
rect 27396 14320 27398 14340
rect 27434 9696 27490 9752
rect 27342 8508 27344 8528
rect 27344 8508 27396 8528
rect 27396 8508 27398 8528
rect 27342 8472 27398 8508
rect 27618 12144 27674 12200
rect 27526 8064 27582 8120
rect 28262 21428 28264 21448
rect 28264 21428 28316 21448
rect 28316 21428 28318 21448
rect 28262 21392 28318 21428
rect 28814 21664 28870 21720
rect 28722 21392 28778 21448
rect 28630 21292 28632 21312
rect 28632 21292 28684 21312
rect 28684 21292 28686 21312
rect 28630 21256 28686 21292
rect 28538 21120 28594 21176
rect 28262 18128 28318 18184
rect 28262 17584 28318 17640
rect 28722 18944 28778 19000
rect 28630 18672 28686 18728
rect 28446 18536 28502 18592
rect 28722 18572 28724 18592
rect 28724 18572 28776 18592
rect 28776 18572 28778 18592
rect 28722 18536 28778 18572
rect 28906 18808 28962 18864
rect 28814 18400 28870 18456
rect 28814 18128 28870 18184
rect 28446 17856 28502 17912
rect 28906 17856 28962 17912
rect 28354 15816 28410 15872
rect 28078 15136 28134 15192
rect 28078 11464 28134 11520
rect 27986 11328 28042 11384
rect 27710 8744 27766 8800
rect 28262 13640 28318 13696
rect 28354 12824 28410 12880
rect 28630 12436 28686 12472
rect 28630 12416 28632 12436
rect 28632 12416 28684 12436
rect 28684 12416 28686 12436
rect 28170 11328 28226 11384
rect 28170 10784 28226 10840
rect 27434 7656 27490 7712
rect 27342 7540 27398 7576
rect 27342 7520 27344 7540
rect 27344 7520 27396 7540
rect 27396 7520 27398 7540
rect 27526 7112 27582 7168
rect 26422 3168 26478 3224
rect 27434 6432 27490 6488
rect 27526 5888 27582 5944
rect 26790 5616 26846 5672
rect 26790 4664 26846 4720
rect 26974 2896 27030 2952
rect 27526 3984 27582 4040
rect 27434 3304 27490 3360
rect 27434 2372 27490 2408
rect 27434 2352 27436 2372
rect 27436 2352 27488 2372
rect 27488 2352 27490 2372
rect 27894 3848 27950 3904
rect 28078 6432 28134 6488
rect 28262 8472 28318 8528
rect 28262 5752 28318 5808
rect 28630 11464 28686 11520
rect 29182 17992 29238 18048
rect 29826 22888 29882 22944
rect 30102 23432 30158 23488
rect 29734 19760 29790 19816
rect 29458 18128 29514 18184
rect 29274 12144 29330 12200
rect 28630 6840 28686 6896
rect 29090 10240 29146 10296
rect 28906 7656 28962 7712
rect 30194 21004 30250 21040
rect 30194 20984 30196 21004
rect 30196 20984 30248 21004
rect 30248 20984 30250 21004
rect 30194 19896 30250 19952
rect 30378 19624 30434 19680
rect 30194 18164 30196 18184
rect 30196 18164 30248 18184
rect 30248 18164 30250 18184
rect 30194 18128 30250 18164
rect 29734 15272 29790 15328
rect 30102 17448 30158 17504
rect 30286 15816 30342 15872
rect 30562 20324 30618 20360
rect 30562 20304 30564 20324
rect 30564 20304 30616 20324
rect 30616 20304 30618 20324
rect 30470 17604 30526 17640
rect 30470 17584 30472 17604
rect 30472 17584 30524 17604
rect 30524 17584 30526 17604
rect 30470 17448 30526 17504
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 31206 22888 31262 22944
rect 31758 24792 31814 24848
rect 31482 22516 31484 22536
rect 31484 22516 31536 22536
rect 31536 22516 31538 22536
rect 31482 22480 31538 22516
rect 31574 20440 31630 20496
rect 31298 20032 31354 20088
rect 31206 19780 31262 19816
rect 31206 19760 31208 19780
rect 31208 19760 31260 19780
rect 31260 19760 31262 19780
rect 31574 19760 31630 19816
rect 31758 19488 31814 19544
rect 31574 19080 31630 19136
rect 30838 17312 30894 17368
rect 29642 12552 29698 12608
rect 29458 11600 29514 11656
rect 29642 11328 29698 11384
rect 29458 10920 29514 10976
rect 29550 6024 29606 6080
rect 29642 5480 29698 5536
rect 29182 4020 29184 4040
rect 29184 4020 29236 4040
rect 29236 4020 29238 4040
rect 29182 3984 29238 4020
rect 29918 11736 29974 11792
rect 29826 8336 29882 8392
rect 30286 10920 30342 10976
rect 30470 11192 30526 11248
rect 30378 9560 30434 9616
rect 30562 9424 30618 9480
rect 30562 8472 30618 8528
rect 30470 8064 30526 8120
rect 30378 6704 30434 6760
rect 30194 6296 30250 6352
rect 30286 5888 30342 5944
rect 30562 6568 30618 6624
rect 30378 5752 30434 5808
rect 30470 5480 30526 5536
rect 30194 5344 30250 5400
rect 30378 4800 30434 4856
rect 30102 4664 30158 4720
rect 30286 4276 30342 4312
rect 30286 4256 30288 4276
rect 30288 4256 30340 4276
rect 30340 4256 30342 4276
rect 29918 2624 29974 2680
rect 31022 15680 31078 15736
rect 30746 11464 30802 11520
rect 30746 10784 30802 10840
rect 31942 21020 31944 21040
rect 31944 21020 31996 21040
rect 31996 21020 31998 21040
rect 31942 20984 31998 21020
rect 31022 10784 31078 10840
rect 30838 10376 30894 10432
rect 30654 5888 30710 5944
rect 31022 10512 31078 10568
rect 31206 10512 31262 10568
rect 31022 9152 31078 9208
rect 31022 7656 31078 7712
rect 31206 8200 31262 8256
rect 30930 4256 30986 4312
rect 32494 21956 32550 21992
rect 32494 21936 32496 21956
rect 32496 21936 32548 21956
rect 32548 21936 32550 21956
rect 32126 20032 32182 20088
rect 32310 19624 32366 19680
rect 32310 19372 32366 19408
rect 32310 19352 32312 19372
rect 32312 19352 32364 19372
rect 32364 19352 32366 19372
rect 32770 19760 32826 19816
rect 32678 18264 32734 18320
rect 32954 21800 33010 21856
rect 32954 20324 33010 20360
rect 32954 20304 32956 20324
rect 32956 20304 33008 20324
rect 33008 20304 33010 20324
rect 32954 20168 33010 20224
rect 33046 19896 33102 19952
rect 33046 18284 33102 18320
rect 33046 18264 33048 18284
rect 33048 18264 33100 18284
rect 33100 18264 33102 18284
rect 32310 16904 32366 16960
rect 31666 10376 31722 10432
rect 31482 10140 31484 10160
rect 31484 10140 31536 10160
rect 31536 10140 31538 10160
rect 31482 10104 31538 10140
rect 31574 9832 31630 9888
rect 31482 9560 31538 9616
rect 32034 10668 32090 10704
rect 32034 10648 32036 10668
rect 32036 10648 32088 10668
rect 32088 10648 32090 10668
rect 31942 9152 31998 9208
rect 31850 8880 31906 8936
rect 31666 8236 31668 8256
rect 31668 8236 31720 8256
rect 31720 8236 31722 8256
rect 32034 8608 32090 8664
rect 31666 8200 31722 8236
rect 31574 7692 31576 7712
rect 31576 7692 31628 7712
rect 31628 7692 31630 7712
rect 31574 7656 31630 7692
rect 31482 7112 31538 7168
rect 31574 6976 31630 7032
rect 31942 6976 31998 7032
rect 31574 5616 31630 5672
rect 31758 5616 31814 5672
rect 31482 5344 31538 5400
rect 31574 5208 31630 5264
rect 31850 5344 31906 5400
rect 32218 10260 32274 10296
rect 32218 10240 32220 10260
rect 32220 10240 32272 10260
rect 32272 10240 32274 10260
rect 32310 6568 32366 6624
rect 32402 6296 32458 6352
rect 32770 9152 32826 9208
rect 32678 8744 32734 8800
rect 32770 8608 32826 8664
rect 32126 5752 32182 5808
rect 32310 5208 32366 5264
rect 32218 5108 32220 5128
rect 32220 5108 32272 5128
rect 32272 5108 32274 5128
rect 32218 5072 32274 5108
rect 31298 2488 31354 2544
rect 32586 3712 32642 3768
rect 32586 3032 32642 3088
rect 32954 12960 33010 13016
rect 33322 12824 33378 12880
rect 33322 9832 33378 9888
rect 33230 9016 33286 9072
rect 32862 8064 32918 8120
rect 33230 8744 33286 8800
rect 33138 7656 33194 7712
rect 32954 7248 33010 7304
rect 32954 6976 33010 7032
rect 32862 4936 32918 4992
rect 33782 16496 33838 16552
rect 36174 38120 36230 38176
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 33966 16632 34022 16688
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 36818 38800 36874 38856
rect 38290 36760 38346 36816
rect 37186 34040 37242 34096
rect 37462 32544 37518 32600
rect 37462 32000 37518 32056
rect 37186 28600 37242 28656
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34242 13096 34298 13152
rect 34518 12824 34574 12880
rect 33690 11600 33746 11656
rect 33598 10104 33654 10160
rect 33690 8608 33746 8664
rect 33598 7812 33654 7848
rect 33598 7792 33600 7812
rect 33600 7792 33652 7812
rect 33652 7792 33654 7812
rect 33506 6840 33562 6896
rect 33690 6296 33746 6352
rect 33874 5344 33930 5400
rect 34242 9832 34298 9888
rect 34058 7540 34114 7576
rect 34058 7520 34060 7540
rect 34060 7520 34112 7540
rect 34112 7520 34114 7540
rect 34426 8336 34482 8392
rect 34242 7112 34298 7168
rect 34058 5072 34114 5128
rect 34334 5616 34390 5672
rect 34334 5480 34390 5536
rect 34242 4800 34298 4856
rect 34426 3304 34482 3360
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34794 6296 34850 6352
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35622 9968 35678 10024
rect 35898 12144 35954 12200
rect 35714 7384 35770 7440
rect 35714 6432 35770 6488
rect 35806 6296 35862 6352
rect 34886 5108 34888 5128
rect 34888 5108 34940 5128
rect 34940 5108 34942 5128
rect 34886 5072 34942 5108
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35254 3440 35310 3496
rect 34794 2896 34850 2952
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35622 4020 35624 4040
rect 35624 4020 35676 4040
rect 35676 4020 35678 4040
rect 35622 3984 35678 4020
rect 36082 11056 36138 11112
rect 36266 6704 36322 6760
rect 36174 5752 36230 5808
rect 35806 2760 35862 2816
rect 35714 1400 35770 1456
rect 38198 36080 38254 36136
rect 38198 34720 38254 34776
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38198 31320 38254 31376
rect 38106 29960 38162 30016
rect 38198 29280 38254 29336
rect 38290 27240 38346 27296
rect 38290 26560 38346 26616
rect 36634 15544 36690 15600
rect 37278 15408 37334 15464
rect 36450 6704 36506 6760
rect 36818 8880 36874 8936
rect 36726 5480 36782 5536
rect 36634 4664 36690 4720
rect 36818 4120 36874 4176
rect 37462 11228 37464 11248
rect 37464 11228 37516 11248
rect 37516 11228 37518 11248
rect 37462 11192 37518 11228
rect 37370 10920 37426 10976
rect 38198 25200 38254 25256
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38290 23840 38346 23896
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38290 21800 38346 21856
rect 38290 20440 38346 20496
rect 38106 19780 38162 19816
rect 38106 19760 38108 19780
rect 38108 19760 38160 19780
rect 38160 19760 38162 19780
rect 38290 19080 38346 19136
rect 38106 17720 38162 17776
rect 38290 17040 38346 17096
rect 38474 16360 38530 16416
rect 38198 15680 38254 15736
rect 38198 15000 38254 15056
rect 38198 14320 38254 14376
rect 38290 12960 38346 13016
rect 38198 12688 38254 12744
rect 38106 12280 38162 12336
rect 38106 10920 38162 10976
rect 38106 10240 38162 10296
rect 38198 8880 38254 8936
rect 38198 8200 38254 8256
rect 38198 7520 38254 7576
rect 38198 6160 38254 6216
rect 38198 3576 38254 3632
rect 38382 5480 38438 5536
rect 38290 3440 38346 3496
rect 38934 3304 38990 3360
rect 37554 720 37610 776
<< metal3 >>
rect 200 38858 800 38888
rect 2865 38858 2931 38861
rect 200 38856 2931 38858
rect 200 38800 2870 38856
rect 2926 38800 2931 38856
rect 200 38798 2931 38800
rect 200 38768 800 38798
rect 2865 38795 2931 38798
rect 36813 38858 36879 38861
rect 39200 38858 39800 38888
rect 36813 38856 39800 38858
rect 36813 38800 36818 38856
rect 36874 38800 39800 38856
rect 36813 38798 39800 38800
rect 36813 38795 36879 38798
rect 39200 38768 39800 38798
rect 200 38178 800 38208
rect 3141 38178 3207 38181
rect 200 38176 3207 38178
rect 200 38120 3146 38176
rect 3202 38120 3207 38176
rect 200 38118 3207 38120
rect 200 38088 800 38118
rect 3141 38115 3207 38118
rect 36169 38178 36235 38181
rect 39200 38178 39800 38208
rect 36169 38176 39800 38178
rect 36169 38120 36174 38176
rect 36230 38120 39800 38176
rect 36169 38118 39800 38120
rect 36169 38115 36235 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 1577 36818 1643 36821
rect 200 36816 1643 36818
rect 200 36760 1582 36816
rect 1638 36760 1643 36816
rect 200 36758 1643 36760
rect 200 36728 800 36758
rect 1577 36755 1643 36758
rect 38285 36818 38351 36821
rect 39200 36818 39800 36848
rect 38285 36816 39800 36818
rect 38285 36760 38290 36816
rect 38346 36760 39800 36816
rect 38285 36758 39800 36760
rect 38285 36755 38351 36758
rect 39200 36728 39800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 36048 800 36078
rect 1669 36075 1735 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35458 800 35488
rect 1761 35458 1827 35461
rect 200 35456 1827 35458
rect 200 35400 1766 35456
rect 1822 35400 1827 35456
rect 200 35398 1827 35400
rect 200 35368 800 35398
rect 1761 35395 1827 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 37181 34098 37247 34101
rect 39200 34098 39800 34128
rect 37181 34096 39800 34098
rect 37181 34040 37186 34096
rect 37242 34040 39800 34096
rect 37181 34038 39800 34040
rect 37181 34035 37247 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 24158 32540 24164 32604
rect 24228 32602 24234 32604
rect 37457 32602 37523 32605
rect 24228 32600 37523 32602
rect 24228 32544 37462 32600
rect 37518 32544 37523 32600
rect 24228 32542 37523 32544
rect 24228 32540 24234 32542
rect 37457 32539 37523 32542
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31968 800 31998
rect 1577 31995 1643 31998
rect 37457 32058 37523 32061
rect 39200 32058 39800 32088
rect 37457 32056 39800 32058
rect 37457 32000 37462 32056
rect 37518 32000 39800 32056
rect 37457 31998 39800 32000
rect 37457 31995 37523 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1761 31378 1827 31381
rect 200 31376 1827 31378
rect 200 31320 1766 31376
rect 1822 31320 1827 31376
rect 200 31318 1827 31320
rect 200 31288 800 31318
rect 1761 31315 1827 31318
rect 38193 31378 38259 31381
rect 39200 31378 39800 31408
rect 38193 31376 39800 31378
rect 38193 31320 38198 31376
rect 38254 31320 39800 31376
rect 38193 31318 39800 31320
rect 38193 31315 38259 31318
rect 39200 31288 39800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4838 30092 4844 30156
rect 4908 30154 4914 30156
rect 24853 30154 24919 30157
rect 4908 30152 24919 30154
rect 4908 30096 24858 30152
rect 24914 30096 24919 30152
rect 4908 30094 24919 30096
rect 4908 30092 4914 30094
rect 24853 30091 24919 30094
rect 38101 30018 38167 30021
rect 39200 30018 39800 30048
rect 38101 30016 39800 30018
rect 38101 29960 38106 30016
rect 38162 29960 39800 30016
rect 38101 29958 39800 29960
rect 38101 29955 38167 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 9070 29684 9076 29748
rect 9140 29746 9146 29748
rect 18229 29746 18295 29749
rect 9140 29744 18295 29746
rect 9140 29688 18234 29744
rect 18290 29688 18295 29744
rect 9140 29686 18295 29688
rect 9140 29684 9146 29686
rect 18229 29683 18295 29686
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 38193 29338 38259 29341
rect 39200 29338 39800 29368
rect 38193 29336 39800 29338
rect 38193 29280 38198 29336
rect 38254 29280 39800 29336
rect 38193 29278 39800 29280
rect 38193 29275 38259 29278
rect 39200 29248 39800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 37181 28658 37247 28661
rect 39200 28658 39800 28688
rect 37181 28656 39800 28658
rect 37181 28600 37186 28656
rect 37242 28600 39800 28656
rect 37181 28598 39800 28600
rect 37181 28595 37247 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 22369 27978 22435 27981
rect 25865 27978 25931 27981
rect 27153 27978 27219 27981
rect 22369 27976 27219 27978
rect 22369 27920 22374 27976
rect 22430 27920 25870 27976
rect 25926 27920 27158 27976
rect 27214 27920 27219 27976
rect 22369 27918 27219 27920
rect 22369 27915 22435 27918
rect 25865 27915 25931 27918
rect 27153 27915 27219 27918
rect 21173 27842 21239 27845
rect 25405 27842 25471 27845
rect 25773 27842 25839 27845
rect 21173 27840 25839 27842
rect 21173 27784 21178 27840
rect 21234 27784 25410 27840
rect 25466 27784 25778 27840
rect 25834 27784 25839 27840
rect 21173 27782 25839 27784
rect 21173 27779 21239 27782
rect 25405 27779 25471 27782
rect 25773 27779 25839 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 22185 27706 22251 27709
rect 23422 27706 23428 27708
rect 22185 27704 23428 27706
rect 22185 27648 22190 27704
rect 22246 27648 23428 27704
rect 22185 27646 23428 27648
rect 22185 27643 22251 27646
rect 23422 27644 23428 27646
rect 23492 27644 23498 27708
rect 24117 27434 24183 27437
rect 28165 27434 28231 27437
rect 24117 27432 28231 27434
rect 24117 27376 24122 27432
rect 24178 27376 28170 27432
rect 28226 27376 28231 27432
rect 24117 27374 28231 27376
rect 24117 27371 24183 27374
rect 28165 27371 28231 27374
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 8477 27300 8543 27301
rect 8477 27298 8524 27300
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 8432 27296 8524 27298
rect 8432 27240 8482 27296
rect 8432 27238 8524 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 8477 27236 8524 27238
rect 8588 27236 8594 27300
rect 38285 27298 38351 27301
rect 39200 27298 39800 27328
rect 38285 27296 39800 27298
rect 38285 27240 38290 27296
rect 38346 27240 39800 27296
rect 38285 27238 39800 27240
rect 8477 27235 8543 27236
rect 38285 27235 38351 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 841 27026 907 27029
rect 15837 27026 15903 27029
rect 841 27024 15903 27026
rect 841 26968 846 27024
rect 902 26968 15842 27024
rect 15898 26968 15903 27024
rect 841 26966 15903 26968
rect 841 26963 907 26966
rect 15837 26963 15903 26966
rect 23473 26890 23539 26893
rect 27153 26890 27219 26893
rect 23473 26888 27219 26890
rect 23473 26832 23478 26888
rect 23534 26832 27158 26888
rect 27214 26832 27219 26888
rect 23473 26830 27219 26832
rect 23473 26827 23539 26830
rect 27153 26827 27219 26830
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1761 26618 1827 26621
rect 200 26616 1827 26618
rect 200 26560 1766 26616
rect 1822 26560 1827 26616
rect 200 26558 1827 26560
rect 200 26528 800 26558
rect 1761 26555 1827 26558
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 11237 26482 11303 26485
rect 12801 26482 12867 26485
rect 18781 26482 18847 26485
rect 11237 26480 18847 26482
rect 11237 26424 11242 26480
rect 11298 26424 12806 26480
rect 12862 26424 18786 26480
rect 18842 26424 18847 26480
rect 11237 26422 18847 26424
rect 11237 26419 11303 26422
rect 12801 26419 12867 26422
rect 18781 26419 18847 26422
rect 20161 26482 20227 26485
rect 24945 26482 25011 26485
rect 20161 26480 25011 26482
rect 20161 26424 20166 26480
rect 20222 26424 24950 26480
rect 25006 26424 25011 26480
rect 20161 26422 25011 26424
rect 20161 26419 20227 26422
rect 24945 26419 25011 26422
rect 24209 26346 24275 26349
rect 28533 26346 28599 26349
rect 24209 26344 28599 26346
rect 24209 26288 24214 26344
rect 24270 26288 28538 26344
rect 28594 26288 28599 26344
rect 24209 26286 28599 26288
rect 24209 26283 24275 26286
rect 28533 26283 28599 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 12893 26074 12959 26077
rect 17677 26074 17743 26077
rect 12893 26072 17743 26074
rect 12893 26016 12898 26072
rect 12954 26016 17682 26072
rect 17738 26016 17743 26072
rect 12893 26014 17743 26016
rect 12893 26011 12959 26014
rect 17677 26011 17743 26014
rect 18965 25938 19031 25941
rect 25129 25938 25195 25941
rect 18965 25936 25195 25938
rect 18965 25880 18970 25936
rect 19026 25880 25134 25936
rect 25190 25880 25195 25936
rect 18965 25878 25195 25880
rect 18965 25875 19031 25878
rect 25129 25875 25195 25878
rect 13077 25802 13143 25805
rect 19149 25802 19215 25805
rect 13077 25800 19215 25802
rect 13077 25744 13082 25800
rect 13138 25744 19154 25800
rect 19210 25744 19215 25800
rect 13077 25742 19215 25744
rect 13077 25739 13143 25742
rect 19149 25739 19215 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 14549 25394 14615 25397
rect 20294 25394 20300 25396
rect 14549 25392 20300 25394
rect 14549 25336 14554 25392
rect 14610 25336 20300 25392
rect 14549 25334 20300 25336
rect 14549 25331 14615 25334
rect 20294 25332 20300 25334
rect 20364 25394 20370 25396
rect 20621 25394 20687 25397
rect 20364 25392 20687 25394
rect 20364 25336 20626 25392
rect 20682 25336 20687 25392
rect 20364 25334 20687 25336
rect 20364 25332 20370 25334
rect 20621 25331 20687 25334
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 20253 25258 20319 25261
rect 20478 25258 20484 25260
rect 20253 25256 20484 25258
rect 20253 25200 20258 25256
rect 20314 25200 20484 25256
rect 20253 25198 20484 25200
rect 20253 25195 20319 25198
rect 20478 25196 20484 25198
rect 20548 25196 20554 25260
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 17534 24924 17540 24988
rect 17604 24986 17610 24988
rect 18505 24986 18571 24989
rect 17604 24984 18571 24986
rect 17604 24928 18510 24984
rect 18566 24928 18571 24984
rect 17604 24926 18571 24928
rect 17604 24924 17610 24926
rect 18505 24923 18571 24926
rect 24577 24986 24643 24989
rect 27429 24986 27495 24989
rect 24577 24984 27495 24986
rect 24577 24928 24582 24984
rect 24638 24928 27434 24984
rect 27490 24928 27495 24984
rect 24577 24926 27495 24928
rect 24577 24923 24643 24926
rect 27429 24923 27495 24926
rect 11697 24850 11763 24853
rect 12014 24850 12020 24852
rect 11697 24848 12020 24850
rect 11697 24792 11702 24848
rect 11758 24792 12020 24848
rect 11697 24790 12020 24792
rect 11697 24787 11763 24790
rect 12014 24788 12020 24790
rect 12084 24788 12090 24852
rect 26969 24850 27035 24853
rect 31753 24850 31819 24853
rect 26969 24848 31819 24850
rect 26969 24792 26974 24848
rect 27030 24792 31758 24848
rect 31814 24792 31819 24848
rect 26969 24790 31819 24792
rect 26969 24787 27035 24790
rect 31753 24787 31819 24790
rect 18413 24716 18479 24717
rect 18413 24714 18460 24716
rect 18368 24712 18460 24714
rect 18524 24714 18530 24716
rect 25405 24714 25471 24717
rect 18524 24712 25471 24714
rect 18368 24656 18418 24712
rect 18524 24656 25410 24712
rect 25466 24656 25471 24712
rect 18368 24654 18460 24656
rect 18413 24652 18460 24654
rect 18524 24654 25471 24656
rect 18524 24652 18530 24654
rect 18413 24651 18479 24652
rect 25405 24651 25471 24654
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 19609 24578 19675 24581
rect 26233 24578 26299 24581
rect 19609 24576 26299 24578
rect 19609 24520 19614 24576
rect 19670 24520 26238 24576
rect 26294 24520 26299 24576
rect 19609 24518 26299 24520
rect 19609 24515 19675 24518
rect 26233 24515 26299 24518
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 15009 24442 15075 24445
rect 17309 24442 17375 24445
rect 15009 24440 17375 24442
rect 15009 24384 15014 24440
rect 15070 24384 17314 24440
rect 17370 24384 17375 24440
rect 15009 24382 17375 24384
rect 15009 24379 15075 24382
rect 17309 24379 17375 24382
rect 19885 24442 19951 24445
rect 25313 24442 25379 24445
rect 19885 24440 25379 24442
rect 19885 24384 19890 24440
rect 19946 24384 25318 24440
rect 25374 24384 25379 24440
rect 19885 24382 25379 24384
rect 19885 24379 19951 24382
rect 25313 24379 25379 24382
rect 20437 24306 20503 24309
rect 20302 24304 20503 24306
rect 20302 24248 20442 24304
rect 20498 24248 20503 24304
rect 20302 24246 20503 24248
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 1894 23428 1900 23492
rect 1964 23490 1970 23492
rect 2589 23490 2655 23493
rect 1964 23488 2655 23490
rect 1964 23432 2594 23488
rect 2650 23432 2655 23488
rect 1964 23430 2655 23432
rect 1964 23428 1970 23430
rect 2589 23427 2655 23430
rect 18270 23428 18276 23492
rect 18340 23490 18346 23492
rect 18413 23490 18479 23493
rect 18340 23488 18479 23490
rect 18340 23432 18418 23488
rect 18474 23432 18479 23488
rect 18340 23430 18479 23432
rect 18340 23428 18346 23430
rect 18413 23427 18479 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 20302 23357 20362 24246
rect 20437 24243 20503 24246
rect 20437 23898 20503 23901
rect 24945 23898 25011 23901
rect 20437 23896 25011 23898
rect 20437 23840 20442 23896
rect 20498 23840 24950 23896
rect 25006 23840 25011 23896
rect 20437 23838 25011 23840
rect 20437 23835 20503 23838
rect 24945 23835 25011 23838
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 22870 23700 22876 23764
rect 22940 23762 22946 23764
rect 23197 23762 23263 23765
rect 24209 23762 24275 23765
rect 22940 23760 24275 23762
rect 22940 23704 23202 23760
rect 23258 23704 24214 23760
rect 24270 23704 24275 23760
rect 22940 23702 24275 23704
rect 22940 23700 22946 23702
rect 23197 23699 23263 23702
rect 24209 23699 24275 23702
rect 23197 23626 23263 23629
rect 23606 23626 23612 23628
rect 23197 23624 23612 23626
rect 23197 23568 23202 23624
rect 23258 23568 23612 23624
rect 23197 23566 23612 23568
rect 23197 23563 23263 23566
rect 23606 23564 23612 23566
rect 23676 23626 23682 23628
rect 23841 23626 23907 23629
rect 23676 23624 23907 23626
rect 23676 23568 23846 23624
rect 23902 23568 23907 23624
rect 23676 23566 23907 23568
rect 23676 23564 23682 23566
rect 23841 23563 23907 23566
rect 20713 23490 20779 23493
rect 27521 23490 27587 23493
rect 30097 23492 30163 23493
rect 20713 23488 27587 23490
rect 20713 23432 20718 23488
rect 20774 23432 27526 23488
rect 27582 23432 27587 23488
rect 20713 23430 27587 23432
rect 20713 23427 20779 23430
rect 27521 23427 27587 23430
rect 30046 23428 30052 23492
rect 30116 23490 30163 23492
rect 30116 23488 30208 23490
rect 30158 23432 30208 23488
rect 30116 23430 30208 23432
rect 30116 23428 30163 23430
rect 30097 23427 30163 23428
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 20302 23352 20411 23357
rect 20302 23296 20350 23352
rect 20406 23296 20411 23352
rect 20302 23294 20411 23296
rect 20345 23291 20411 23294
rect 19885 23218 19951 23221
rect 26877 23218 26943 23221
rect 19885 23216 26943 23218
rect 19885 23160 19890 23216
rect 19946 23160 26882 23216
rect 26938 23160 26943 23216
rect 19885 23158 26943 23160
rect 19885 23155 19951 23158
rect 26877 23155 26943 23158
rect 16481 23082 16547 23085
rect 36854 23082 36860 23084
rect 16481 23080 36860 23082
rect 16481 23024 16486 23080
rect 16542 23024 36860 23080
rect 16481 23022 36860 23024
rect 16481 23019 16547 23022
rect 36854 23020 36860 23022
rect 36924 23020 36930 23084
rect 26693 22946 26759 22949
rect 26918 22946 26924 22948
rect 26693 22944 26924 22946
rect 26693 22888 26698 22944
rect 26754 22888 26924 22944
rect 26693 22886 26924 22888
rect 26693 22883 26759 22886
rect 26918 22884 26924 22886
rect 26988 22884 26994 22948
rect 27705 22946 27771 22949
rect 28206 22946 28212 22948
rect 27705 22944 28212 22946
rect 27705 22888 27710 22944
rect 27766 22888 28212 22944
rect 27705 22886 28212 22888
rect 27705 22883 27771 22886
rect 28206 22884 28212 22886
rect 28276 22884 28282 22948
rect 29821 22946 29887 22949
rect 31201 22946 31267 22949
rect 29821 22944 31267 22946
rect 29821 22888 29826 22944
rect 29882 22888 31206 22944
rect 31262 22888 31267 22944
rect 29821 22886 31267 22888
rect 29821 22883 29887 22886
rect 31201 22883 31267 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 13721 22674 13787 22677
rect 20110 22674 20116 22676
rect 13721 22672 20116 22674
rect 13721 22616 13726 22672
rect 13782 22616 20116 22672
rect 13721 22614 20116 22616
rect 13721 22611 13787 22614
rect 20110 22612 20116 22614
rect 20180 22612 20186 22676
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 31477 22540 31543 22541
rect 31477 22536 31524 22540
rect 31588 22538 31594 22540
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 31477 22480 31482 22536
rect 31477 22476 31524 22480
rect 31588 22478 31634 22538
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 31588 22476 31594 22478
rect 31477 22475 31543 22476
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19517 22266 19583 22269
rect 19517 22264 19994 22266
rect 19517 22208 19522 22264
rect 19578 22208 19994 22264
rect 19517 22206 19994 22208
rect 19517 22203 19583 22206
rect 19934 22130 19994 22206
rect 20069 22130 20135 22133
rect 19934 22128 20135 22130
rect 19934 22072 20074 22128
rect 20130 22072 20135 22128
rect 19934 22070 20135 22072
rect 20069 22067 20135 22070
rect 20253 22130 20319 22133
rect 20253 22128 26618 22130
rect 20253 22072 20258 22128
rect 20314 22072 26618 22128
rect 20253 22070 26618 22072
rect 20253 22067 20319 22070
rect 19333 21994 19399 21997
rect 20161 21994 20227 21997
rect 22737 21996 22803 21997
rect 19333 21992 20227 21994
rect 19333 21936 19338 21992
rect 19394 21936 20166 21992
rect 20222 21936 20227 21992
rect 19333 21934 20227 21936
rect 19333 21931 19399 21934
rect 20161 21931 20227 21934
rect 22686 21932 22692 21996
rect 22756 21994 22803 21996
rect 22756 21992 22848 21994
rect 22798 21936 22848 21992
rect 22756 21934 22848 21936
rect 22756 21932 22803 21934
rect 22737 21931 22803 21932
rect 200 21858 800 21888
rect 1761 21858 1827 21861
rect 200 21856 1827 21858
rect 200 21800 1766 21856
rect 1822 21800 1827 21856
rect 200 21798 1827 21800
rect 26558 21858 26618 22070
rect 27245 21994 27311 21997
rect 32489 21994 32555 21997
rect 27245 21992 32555 21994
rect 27245 21936 27250 21992
rect 27306 21936 32494 21992
rect 32550 21936 32555 21992
rect 27245 21934 32555 21936
rect 27245 21931 27311 21934
rect 32489 21931 32555 21934
rect 32254 21858 32260 21860
rect 26558 21798 32260 21858
rect 200 21768 800 21798
rect 1761 21795 1827 21798
rect 32254 21796 32260 21798
rect 32324 21858 32330 21860
rect 32949 21858 33015 21861
rect 32324 21856 33015 21858
rect 32324 21800 32954 21856
rect 33010 21800 33015 21856
rect 32324 21798 33015 21800
rect 32324 21796 32330 21798
rect 32949 21795 33015 21798
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 10317 21722 10383 21725
rect 16389 21722 16455 21725
rect 10317 21720 16455 21722
rect 10317 21664 10322 21720
rect 10378 21664 16394 21720
rect 16450 21664 16455 21720
rect 10317 21662 16455 21664
rect 10317 21659 10383 21662
rect 16389 21659 16455 21662
rect 22277 21722 22343 21725
rect 28809 21722 28875 21725
rect 22277 21720 28875 21722
rect 22277 21664 22282 21720
rect 22338 21664 28814 21720
rect 28870 21664 28875 21720
rect 22277 21662 28875 21664
rect 22277 21659 22343 21662
rect 28809 21659 28875 21662
rect 12525 21586 12591 21589
rect 13353 21586 13419 21589
rect 12525 21584 13419 21586
rect 12525 21528 12530 21584
rect 12586 21528 13358 21584
rect 13414 21528 13419 21584
rect 12525 21526 13419 21528
rect 12525 21523 12591 21526
rect 13353 21523 13419 21526
rect 23565 21586 23631 21589
rect 25773 21586 25839 21589
rect 23565 21584 25839 21586
rect 23565 21528 23570 21584
rect 23626 21528 25778 21584
rect 25834 21528 25839 21584
rect 23565 21526 25839 21528
rect 23565 21523 23631 21526
rect 25773 21523 25839 21526
rect 11697 21450 11763 21453
rect 11830 21450 11836 21452
rect 11697 21448 11836 21450
rect 11697 21392 11702 21448
rect 11758 21392 11836 21448
rect 11697 21390 11836 21392
rect 11697 21387 11763 21390
rect 11830 21388 11836 21390
rect 11900 21388 11906 21452
rect 20897 21450 20963 21453
rect 21398 21450 21404 21452
rect 20897 21448 21404 21450
rect 20897 21392 20902 21448
rect 20958 21392 21404 21448
rect 20897 21390 21404 21392
rect 20897 21387 20963 21390
rect 21398 21388 21404 21390
rect 21468 21388 21474 21452
rect 22553 21450 22619 21453
rect 25957 21450 26023 21453
rect 27654 21450 27660 21452
rect 22553 21448 27660 21450
rect 22553 21392 22558 21448
rect 22614 21392 25962 21448
rect 26018 21392 27660 21448
rect 22553 21390 27660 21392
rect 22553 21387 22619 21390
rect 25957 21387 26023 21390
rect 27654 21388 27660 21390
rect 27724 21388 27730 21452
rect 28257 21450 28323 21453
rect 28717 21450 28783 21453
rect 28257 21448 28783 21450
rect 28257 21392 28262 21448
rect 28318 21392 28722 21448
rect 28778 21392 28783 21448
rect 28257 21390 28783 21392
rect 28257 21387 28323 21390
rect 28717 21387 28783 21390
rect 27429 21314 27495 21317
rect 27705 21314 27771 21317
rect 28625 21314 28691 21317
rect 27429 21312 28691 21314
rect 27429 21256 27434 21312
rect 27490 21256 27710 21312
rect 27766 21256 28630 21312
rect 28686 21256 28691 21312
rect 27429 21254 28691 21256
rect 27429 21251 27495 21254
rect 27705 21251 27771 21254
rect 28625 21251 28691 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 17166 21116 17172 21180
rect 17236 21178 17242 21180
rect 20989 21178 21055 21181
rect 17236 21176 21055 21178
rect 17236 21120 20994 21176
rect 21050 21120 21055 21176
rect 17236 21118 21055 21120
rect 17236 21116 17242 21118
rect 20989 21115 21055 21118
rect 22829 21178 22895 21181
rect 23289 21178 23355 21181
rect 28533 21178 28599 21181
rect 22829 21176 28599 21178
rect 22829 21120 22834 21176
rect 22890 21120 23294 21176
rect 23350 21120 28538 21176
rect 28594 21120 28599 21176
rect 22829 21118 28599 21120
rect 22829 21115 22895 21118
rect 23289 21115 23355 21118
rect 28533 21115 28599 21118
rect 21541 21042 21607 21045
rect 25681 21042 25747 21045
rect 21541 21040 25747 21042
rect 21541 20984 21546 21040
rect 21602 20984 25686 21040
rect 25742 20984 25747 21040
rect 21541 20982 25747 20984
rect 21541 20979 21607 20982
rect 25681 20979 25747 20982
rect 30189 21042 30255 21045
rect 31937 21042 32003 21045
rect 30189 21040 32003 21042
rect 30189 20984 30194 21040
rect 30250 20984 31942 21040
rect 31998 20984 32003 21040
rect 30189 20982 32003 20984
rect 30189 20979 30255 20982
rect 31937 20979 32003 20982
rect 13629 20906 13695 20909
rect 17677 20906 17743 20909
rect 13629 20904 17743 20906
rect 13629 20848 13634 20904
rect 13690 20848 17682 20904
rect 17738 20848 17743 20904
rect 13629 20846 17743 20848
rect 13629 20843 13695 20846
rect 17677 20843 17743 20846
rect 20253 20906 20319 20909
rect 20529 20906 20595 20909
rect 20253 20904 20595 20906
rect 20253 20848 20258 20904
rect 20314 20848 20534 20904
rect 20590 20848 20595 20904
rect 20253 20846 20595 20848
rect 20253 20843 20319 20846
rect 20529 20843 20595 20846
rect 23473 20906 23539 20909
rect 23933 20906 23999 20909
rect 28206 20906 28212 20908
rect 23473 20904 28212 20906
rect 23473 20848 23478 20904
rect 23534 20848 23938 20904
rect 23994 20848 28212 20904
rect 23473 20846 28212 20848
rect 23473 20843 23539 20846
rect 23933 20843 23999 20846
rect 28206 20844 28212 20846
rect 28276 20844 28282 20908
rect 13353 20770 13419 20773
rect 22001 20772 22067 20773
rect 13486 20770 13492 20772
rect 13353 20768 13492 20770
rect 13353 20712 13358 20768
rect 13414 20712 13492 20768
rect 13353 20710 13492 20712
rect 13353 20707 13419 20710
rect 13486 20708 13492 20710
rect 13556 20708 13562 20772
rect 21950 20770 21956 20772
rect 21910 20710 21956 20770
rect 22020 20768 22067 20772
rect 22062 20712 22067 20768
rect 21950 20708 21956 20710
rect 22020 20708 22067 20712
rect 23422 20708 23428 20772
rect 23492 20770 23498 20772
rect 24710 20770 24716 20772
rect 23492 20710 24716 20770
rect 23492 20708 23498 20710
rect 24710 20708 24716 20710
rect 24780 20708 24786 20772
rect 24945 20770 25011 20773
rect 25262 20770 25268 20772
rect 24945 20768 25268 20770
rect 24945 20712 24950 20768
rect 25006 20712 25268 20768
rect 24945 20710 25268 20712
rect 22001 20707 22067 20708
rect 24945 20707 25011 20710
rect 25262 20708 25268 20710
rect 25332 20708 25338 20772
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 19057 20498 19123 20501
rect 22134 20498 22140 20500
rect 19057 20496 22140 20498
rect 19057 20440 19062 20496
rect 19118 20440 22140 20496
rect 19057 20438 22140 20440
rect 19057 20435 19123 20438
rect 22134 20436 22140 20438
rect 22204 20436 22210 20500
rect 27061 20498 27127 20501
rect 31569 20498 31635 20501
rect 27061 20496 31635 20498
rect 27061 20440 27066 20496
rect 27122 20440 31574 20496
rect 31630 20440 31635 20496
rect 27061 20438 31635 20440
rect 27061 20435 27127 20438
rect 31569 20435 31635 20438
rect 38285 20498 38351 20501
rect 39200 20498 39800 20528
rect 38285 20496 39800 20498
rect 38285 20440 38290 20496
rect 38346 20440 39800 20496
rect 38285 20438 39800 20440
rect 38285 20435 38351 20438
rect 39200 20408 39800 20438
rect 20897 20362 20963 20365
rect 21030 20362 21036 20364
rect 20897 20360 21036 20362
rect 20897 20304 20902 20360
rect 20958 20304 21036 20360
rect 20897 20302 21036 20304
rect 20897 20299 20963 20302
rect 21030 20300 21036 20302
rect 21100 20300 21106 20364
rect 30557 20362 30623 20365
rect 32949 20362 33015 20365
rect 30557 20360 33015 20362
rect 30557 20304 30562 20360
rect 30618 20304 32954 20360
rect 33010 20304 33015 20360
rect 30557 20302 33015 20304
rect 30557 20299 30623 20302
rect 32949 20299 33015 20302
rect 25865 20226 25931 20229
rect 32949 20226 33015 20229
rect 25865 20224 33015 20226
rect 25865 20168 25870 20224
rect 25926 20168 32954 20224
rect 33010 20168 33015 20224
rect 25865 20166 33015 20168
rect 25865 20163 25931 20166
rect 32949 20163 33015 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 31293 20090 31359 20093
rect 32121 20090 32187 20093
rect 31293 20088 32187 20090
rect 31293 20032 31298 20088
rect 31354 20032 32126 20088
rect 32182 20032 32187 20088
rect 31293 20030 32187 20032
rect 31293 20027 31359 20030
rect 32121 20027 32187 20030
rect 12341 19954 12407 19957
rect 12709 19954 12775 19957
rect 15837 19954 15903 19957
rect 12341 19952 15903 19954
rect 12341 19896 12346 19952
rect 12402 19896 12714 19952
rect 12770 19896 15842 19952
rect 15898 19896 15903 19952
rect 12341 19894 15903 19896
rect 12341 19891 12407 19894
rect 12709 19891 12775 19894
rect 15837 19891 15903 19894
rect 20989 19954 21055 19957
rect 27981 19954 28047 19957
rect 20989 19952 28047 19954
rect 20989 19896 20994 19952
rect 21050 19896 27986 19952
rect 28042 19896 28047 19952
rect 20989 19894 28047 19896
rect 20989 19891 21055 19894
rect 27981 19891 28047 19894
rect 30189 19954 30255 19957
rect 33041 19954 33107 19957
rect 30189 19952 33107 19954
rect 30189 19896 30194 19952
rect 30250 19896 33046 19952
rect 33102 19896 33107 19952
rect 30189 19894 33107 19896
rect 30189 19891 30255 19894
rect 33041 19891 33107 19894
rect 200 19818 800 19848
rect 1577 19818 1643 19821
rect 200 19816 1643 19818
rect 200 19760 1582 19816
rect 1638 19760 1643 19816
rect 200 19758 1643 19760
rect 200 19728 800 19758
rect 1577 19755 1643 19758
rect 5390 19756 5396 19820
rect 5460 19818 5466 19820
rect 15469 19818 15535 19821
rect 5460 19816 15535 19818
rect 5460 19760 15474 19816
rect 15530 19760 15535 19816
rect 5460 19758 15535 19760
rect 5460 19756 5466 19758
rect 15469 19755 15535 19758
rect 22369 19818 22435 19821
rect 27889 19818 27955 19821
rect 22369 19816 27955 19818
rect 22369 19760 22374 19816
rect 22430 19760 27894 19816
rect 27950 19760 27955 19816
rect 22369 19758 27955 19760
rect 22369 19755 22435 19758
rect 27889 19755 27955 19758
rect 29729 19818 29795 19821
rect 31201 19818 31267 19821
rect 29729 19816 31267 19818
rect 29729 19760 29734 19816
rect 29790 19760 31206 19816
rect 31262 19760 31267 19816
rect 29729 19758 31267 19760
rect 29729 19755 29795 19758
rect 31201 19755 31267 19758
rect 31569 19818 31635 19821
rect 32438 19818 32444 19820
rect 31569 19816 32444 19818
rect 31569 19760 31574 19816
rect 31630 19760 32444 19816
rect 31569 19758 32444 19760
rect 31569 19755 31635 19758
rect 32438 19756 32444 19758
rect 32508 19818 32514 19820
rect 32765 19818 32831 19821
rect 32508 19816 32831 19818
rect 32508 19760 32770 19816
rect 32826 19760 32831 19816
rect 32508 19758 32831 19760
rect 32508 19756 32514 19758
rect 32765 19755 32831 19758
rect 38101 19818 38167 19821
rect 39200 19818 39800 19848
rect 38101 19816 39800 19818
rect 38101 19760 38106 19816
rect 38162 19760 39800 19816
rect 38101 19758 39800 19760
rect 38101 19755 38167 19758
rect 39200 19728 39800 19758
rect 23013 19682 23079 19685
rect 27337 19682 27403 19685
rect 23013 19680 27403 19682
rect 23013 19624 23018 19680
rect 23074 19624 27342 19680
rect 27398 19624 27403 19680
rect 23013 19622 27403 19624
rect 23013 19619 23079 19622
rect 27337 19619 27403 19622
rect 30373 19682 30439 19685
rect 32305 19682 32371 19685
rect 30373 19680 32371 19682
rect 30373 19624 30378 19680
rect 30434 19624 32310 19680
rect 32366 19624 32371 19680
rect 30373 19622 32371 19624
rect 30373 19619 30439 19622
rect 32305 19619 32371 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 13629 19546 13695 19549
rect 18045 19546 18111 19549
rect 13629 19544 18111 19546
rect 13629 19488 13634 19544
rect 13690 19488 18050 19544
rect 18106 19488 18111 19544
rect 13629 19486 18111 19488
rect 13629 19483 13695 19486
rect 18045 19483 18111 19486
rect 27061 19546 27127 19549
rect 31753 19546 31819 19549
rect 27061 19544 31819 19546
rect 27061 19488 27066 19544
rect 27122 19488 31758 19544
rect 31814 19488 31819 19544
rect 27061 19486 31819 19488
rect 27061 19483 27127 19486
rect 31753 19483 31819 19486
rect 17309 19412 17375 19413
rect 17309 19408 17356 19412
rect 17420 19410 17426 19412
rect 22093 19410 22159 19413
rect 31886 19410 31892 19412
rect 17309 19352 17314 19408
rect 17309 19348 17356 19352
rect 17420 19350 17466 19410
rect 22093 19408 31892 19410
rect 22093 19352 22098 19408
rect 22154 19352 31892 19408
rect 22093 19350 31892 19352
rect 17420 19348 17426 19350
rect 17309 19347 17375 19348
rect 22093 19347 22159 19350
rect 31886 19348 31892 19350
rect 31956 19348 31962 19412
rect 32070 19348 32076 19412
rect 32140 19410 32146 19412
rect 32305 19410 32371 19413
rect 32140 19408 32371 19410
rect 32140 19352 32310 19408
rect 32366 19352 32371 19408
rect 32140 19350 32371 19352
rect 32140 19348 32146 19350
rect 32305 19347 32371 19350
rect 3550 19212 3556 19276
rect 3620 19274 3626 19276
rect 26785 19274 26851 19277
rect 3620 19272 26851 19274
rect 3620 19216 26790 19272
rect 26846 19216 26851 19272
rect 3620 19214 26851 19216
rect 3620 19212 3626 19214
rect 26785 19211 26851 19214
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 13486 19076 13492 19140
rect 13556 19138 13562 19140
rect 17718 19138 17724 19140
rect 13556 19078 17724 19138
rect 13556 19076 13562 19078
rect 17718 19076 17724 19078
rect 17788 19076 17794 19140
rect 25814 19076 25820 19140
rect 25884 19138 25890 19140
rect 26141 19138 26207 19141
rect 25884 19136 26207 19138
rect 25884 19080 26146 19136
rect 26202 19080 26207 19136
rect 25884 19078 26207 19080
rect 25884 19076 25890 19078
rect 26141 19075 26207 19078
rect 26785 19138 26851 19141
rect 31569 19138 31635 19141
rect 26785 19136 31635 19138
rect 26785 19080 26790 19136
rect 26846 19080 31574 19136
rect 31630 19080 31635 19136
rect 26785 19078 31635 19080
rect 26785 19075 26851 19078
rect 31569 19075 31635 19078
rect 38285 19138 38351 19141
rect 39200 19138 39800 19168
rect 38285 19136 39800 19138
rect 38285 19080 38290 19136
rect 38346 19080 39800 19136
rect 38285 19078 39800 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 27981 19002 28047 19005
rect 28717 19002 28783 19005
rect 27981 19000 28783 19002
rect 27981 18944 27986 19000
rect 28042 18944 28722 19000
rect 28778 18944 28783 19000
rect 27981 18942 28783 18944
rect 27981 18939 28047 18942
rect 28717 18939 28783 18942
rect 26325 18866 26391 18869
rect 28901 18866 28967 18869
rect 26325 18864 28967 18866
rect 26325 18808 26330 18864
rect 26386 18808 28906 18864
rect 28962 18808 28967 18864
rect 26325 18806 28967 18808
rect 26325 18803 26391 18806
rect 28901 18803 28967 18806
rect 5022 18668 5028 18732
rect 5092 18730 5098 18732
rect 6545 18730 6611 18733
rect 5092 18728 6611 18730
rect 5092 18672 6550 18728
rect 6606 18672 6611 18728
rect 5092 18670 6611 18672
rect 5092 18668 5098 18670
rect 6545 18667 6611 18670
rect 25681 18730 25747 18733
rect 26693 18730 26759 18733
rect 28625 18730 28691 18733
rect 29126 18730 29132 18732
rect 25681 18728 29132 18730
rect 25681 18672 25686 18728
rect 25742 18672 26698 18728
rect 26754 18672 28630 18728
rect 28686 18672 29132 18728
rect 25681 18670 29132 18672
rect 25681 18667 25747 18670
rect 26693 18667 26759 18670
rect 28625 18667 28691 18670
rect 29126 18668 29132 18670
rect 29196 18668 29202 18732
rect 2313 18594 2379 18597
rect 17534 18594 17540 18596
rect 2313 18592 17540 18594
rect 2313 18536 2318 18592
rect 2374 18536 17540 18592
rect 2313 18534 17540 18536
rect 2313 18531 2379 18534
rect 17534 18532 17540 18534
rect 17604 18532 17610 18596
rect 28441 18594 28507 18597
rect 28717 18596 28783 18597
rect 28574 18594 28580 18596
rect 28441 18592 28580 18594
rect 28441 18536 28446 18592
rect 28502 18536 28580 18592
rect 28441 18534 28580 18536
rect 28441 18531 28507 18534
rect 28574 18532 28580 18534
rect 28644 18532 28650 18596
rect 28717 18592 28764 18596
rect 28828 18594 28834 18596
rect 28717 18536 28722 18592
rect 28717 18532 28764 18536
rect 28828 18534 28874 18594
rect 28828 18532 28834 18534
rect 28717 18531 28783 18532
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 27981 18458 28047 18461
rect 28809 18458 28875 18461
rect 27981 18456 28875 18458
rect 27981 18400 27986 18456
rect 28042 18400 28814 18456
rect 28870 18400 28875 18456
rect 27981 18398 28875 18400
rect 27981 18395 28047 18398
rect 28809 18395 28875 18398
rect 19885 18322 19951 18325
rect 20161 18322 20227 18325
rect 19885 18320 20227 18322
rect 19885 18264 19890 18320
rect 19946 18264 20166 18320
rect 20222 18264 20227 18320
rect 19885 18262 20227 18264
rect 19885 18259 19951 18262
rect 20161 18259 20227 18262
rect 27470 18260 27476 18324
rect 27540 18322 27546 18324
rect 32673 18322 32739 18325
rect 33041 18322 33107 18325
rect 27540 18320 33107 18322
rect 27540 18264 32678 18320
rect 32734 18264 33046 18320
rect 33102 18264 33107 18320
rect 27540 18262 33107 18264
rect 27540 18260 27546 18262
rect 32673 18259 32739 18262
rect 33041 18259 33107 18262
rect 12801 18186 12867 18189
rect 18321 18186 18387 18189
rect 12801 18184 18387 18186
rect 12801 18128 12806 18184
rect 12862 18128 18326 18184
rect 18382 18128 18387 18184
rect 12801 18126 18387 18128
rect 12801 18123 12867 18126
rect 18321 18123 18387 18126
rect 20713 18186 20779 18189
rect 25630 18186 25636 18188
rect 20713 18184 25636 18186
rect 20713 18128 20718 18184
rect 20774 18128 25636 18184
rect 20713 18126 25636 18128
rect 20713 18123 20779 18126
rect 25630 18124 25636 18126
rect 25700 18124 25706 18188
rect 26366 18124 26372 18188
rect 26436 18186 26442 18188
rect 28257 18186 28323 18189
rect 26436 18184 28323 18186
rect 26436 18128 28262 18184
rect 28318 18128 28323 18184
rect 26436 18126 28323 18128
rect 26436 18124 26442 18126
rect 28257 18123 28323 18126
rect 28809 18186 28875 18189
rect 28942 18186 28948 18188
rect 28809 18184 28948 18186
rect 28809 18128 28814 18184
rect 28870 18128 28948 18184
rect 28809 18126 28948 18128
rect 28809 18123 28875 18126
rect 28942 18124 28948 18126
rect 29012 18124 29018 18188
rect 29453 18186 29519 18189
rect 30189 18186 30255 18189
rect 30414 18186 30420 18188
rect 29453 18184 30420 18186
rect 29453 18128 29458 18184
rect 29514 18128 30194 18184
rect 30250 18128 30420 18184
rect 29453 18126 30420 18128
rect 29453 18123 29519 18126
rect 30189 18123 30255 18126
rect 30414 18124 30420 18126
rect 30484 18124 30490 18188
rect 9489 18052 9555 18053
rect 9438 18050 9444 18052
rect 9398 17990 9444 18050
rect 9508 18048 9555 18052
rect 9550 17992 9555 18048
rect 9438 17988 9444 17990
rect 9508 17988 9555 17992
rect 9489 17987 9555 17988
rect 19425 18050 19491 18053
rect 20662 18050 20668 18052
rect 19425 18048 20668 18050
rect 19425 17992 19430 18048
rect 19486 17992 20668 18048
rect 19425 17990 20668 17992
rect 19425 17987 19491 17990
rect 20662 17988 20668 17990
rect 20732 17988 20738 18052
rect 23013 18050 23079 18053
rect 25078 18050 25084 18052
rect 23013 18048 25084 18050
rect 23013 17992 23018 18048
rect 23074 17992 25084 18048
rect 23013 17990 25084 17992
rect 23013 17987 23079 17990
rect 25078 17988 25084 17990
rect 25148 17988 25154 18052
rect 26417 18050 26483 18053
rect 26550 18050 26556 18052
rect 26417 18048 26556 18050
rect 26417 17992 26422 18048
rect 26478 17992 26556 18048
rect 26417 17990 26556 17992
rect 26417 17987 26483 17990
rect 26550 17988 26556 17990
rect 26620 17988 26626 18052
rect 26693 18050 26759 18053
rect 29177 18050 29243 18053
rect 26693 18048 29243 18050
rect 26693 17992 26698 18048
rect 26754 17992 29182 18048
rect 29238 17992 29243 18048
rect 26693 17990 29243 17992
rect 26693 17987 26759 17990
rect 29177 17987 29243 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 7598 17852 7604 17916
rect 7668 17914 7674 17916
rect 13261 17914 13327 17917
rect 7668 17912 13327 17914
rect 7668 17856 13266 17912
rect 13322 17856 13327 17912
rect 7668 17854 13327 17856
rect 7668 17852 7674 17854
rect 13261 17851 13327 17854
rect 16481 17914 16547 17917
rect 21449 17914 21515 17917
rect 16481 17912 21515 17914
rect 16481 17856 16486 17912
rect 16542 17856 21454 17912
rect 21510 17856 21515 17912
rect 16481 17854 21515 17856
rect 16481 17851 16547 17854
rect 21449 17851 21515 17854
rect 27245 17914 27311 17917
rect 28441 17914 28507 17917
rect 28901 17916 28967 17917
rect 28901 17914 28948 17916
rect 27245 17912 28507 17914
rect 27245 17856 27250 17912
rect 27306 17856 28446 17912
rect 28502 17856 28507 17912
rect 27245 17854 28507 17856
rect 28856 17912 28948 17914
rect 28856 17856 28906 17912
rect 28856 17854 28948 17856
rect 27245 17851 27311 17854
rect 28441 17851 28507 17854
rect 28901 17852 28948 17854
rect 29012 17852 29018 17916
rect 28901 17851 28967 17852
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 38101 17778 38167 17781
rect 39200 17778 39800 17808
rect 38101 17776 39800 17778
rect 38101 17720 38106 17776
rect 38162 17720 39800 17776
rect 38101 17718 39800 17720
rect 38101 17715 38167 17718
rect 39200 17688 39800 17718
rect 10593 17642 10659 17645
rect 10726 17642 10732 17644
rect 10593 17640 10732 17642
rect 10593 17584 10598 17640
rect 10654 17584 10732 17640
rect 10593 17582 10732 17584
rect 10593 17579 10659 17582
rect 10726 17580 10732 17582
rect 10796 17580 10802 17644
rect 28257 17642 28323 17645
rect 30465 17642 30531 17645
rect 28257 17640 30531 17642
rect 28257 17584 28262 17640
rect 28318 17584 30470 17640
rect 30526 17584 30531 17640
rect 28257 17582 30531 17584
rect 28257 17579 28323 17582
rect 30465 17579 30531 17582
rect 30097 17506 30163 17509
rect 30465 17506 30531 17509
rect 30097 17504 30531 17506
rect 30097 17448 30102 17504
rect 30158 17448 30470 17504
rect 30526 17448 30531 17504
rect 30097 17446 30531 17448
rect 30097 17443 30163 17446
rect 30465 17443 30531 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 25497 17370 25563 17373
rect 28758 17370 28764 17372
rect 25497 17368 28764 17370
rect 25497 17312 25502 17368
rect 25558 17312 28764 17368
rect 25497 17310 28764 17312
rect 25497 17307 25563 17310
rect 28758 17308 28764 17310
rect 28828 17308 28834 17372
rect 30833 17370 30899 17373
rect 32622 17370 32628 17372
rect 30833 17368 32628 17370
rect 30833 17312 30838 17368
rect 30894 17312 32628 17368
rect 30833 17310 32628 17312
rect 30833 17307 30899 17310
rect 32622 17308 32628 17310
rect 32692 17308 32698 17372
rect 13486 17172 13492 17236
rect 13556 17234 13562 17236
rect 24853 17234 24919 17237
rect 13556 17232 24919 17234
rect 13556 17176 24858 17232
rect 24914 17176 24919 17232
rect 13556 17174 24919 17176
rect 13556 17172 13562 17174
rect 24853 17171 24919 17174
rect 200 17098 800 17128
rect 1577 17098 1643 17101
rect 200 17096 1643 17098
rect 200 17040 1582 17096
rect 1638 17040 1643 17096
rect 200 17038 1643 17040
rect 200 17008 800 17038
rect 1577 17035 1643 17038
rect 7782 17036 7788 17100
rect 7852 17098 7858 17100
rect 14365 17098 14431 17101
rect 7852 17096 14431 17098
rect 7852 17040 14370 17096
rect 14426 17040 14431 17096
rect 7852 17038 14431 17040
rect 7852 17036 7858 17038
rect 14365 17035 14431 17038
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 12934 16900 12940 16964
rect 13004 16962 13010 16964
rect 15653 16962 15719 16965
rect 13004 16960 15719 16962
rect 13004 16904 15658 16960
rect 15714 16904 15719 16960
rect 13004 16902 15719 16904
rect 13004 16900 13010 16902
rect 15653 16899 15719 16902
rect 20529 16962 20595 16965
rect 22737 16962 22803 16965
rect 32305 16962 32371 16965
rect 20529 16960 32371 16962
rect 20529 16904 20534 16960
rect 20590 16904 22742 16960
rect 22798 16904 32310 16960
rect 32366 16904 32371 16960
rect 20529 16902 32371 16904
rect 20529 16899 20595 16902
rect 22737 16899 22803 16902
rect 32305 16899 32371 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 16430 16764 16436 16828
rect 16500 16826 16506 16828
rect 18689 16826 18755 16829
rect 16500 16824 18755 16826
rect 16500 16768 18694 16824
rect 18750 16768 18755 16824
rect 16500 16766 18755 16768
rect 16500 16764 16506 16766
rect 18689 16763 18755 16766
rect 9254 16628 9260 16692
rect 9324 16690 9330 16692
rect 9673 16690 9739 16693
rect 9324 16688 9739 16690
rect 9324 16632 9678 16688
rect 9734 16632 9739 16688
rect 9324 16630 9739 16632
rect 9324 16628 9330 16630
rect 9673 16627 9739 16630
rect 14457 16690 14523 16693
rect 14590 16690 14596 16692
rect 14457 16688 14596 16690
rect 14457 16632 14462 16688
rect 14518 16632 14596 16688
rect 14457 16630 14596 16632
rect 14457 16627 14523 16630
rect 14590 16628 14596 16630
rect 14660 16628 14666 16692
rect 14958 16628 14964 16692
rect 15028 16690 15034 16692
rect 15285 16690 15351 16693
rect 15028 16688 15351 16690
rect 15028 16632 15290 16688
rect 15346 16632 15351 16688
rect 15028 16630 15351 16632
rect 15028 16628 15034 16630
rect 15285 16627 15351 16630
rect 15837 16690 15903 16693
rect 18597 16692 18663 16693
rect 16062 16690 16068 16692
rect 15837 16688 16068 16690
rect 15837 16632 15842 16688
rect 15898 16632 16068 16688
rect 15837 16630 16068 16632
rect 15837 16627 15903 16630
rect 16062 16628 16068 16630
rect 16132 16628 16138 16692
rect 18597 16688 18644 16692
rect 18708 16690 18714 16692
rect 25681 16690 25747 16693
rect 18597 16632 18602 16688
rect 18597 16628 18644 16632
rect 18708 16630 18754 16690
rect 25681 16688 29010 16690
rect 25681 16632 25686 16688
rect 25742 16632 29010 16688
rect 25681 16630 29010 16632
rect 18708 16628 18714 16630
rect 18597 16627 18663 16628
rect 25681 16627 25747 16630
rect 11094 16492 11100 16556
rect 11164 16554 11170 16556
rect 11789 16554 11855 16557
rect 11164 16552 11855 16554
rect 11164 16496 11794 16552
rect 11850 16496 11855 16552
rect 11164 16494 11855 16496
rect 11164 16492 11170 16494
rect 11789 16491 11855 16494
rect 13629 16554 13695 16557
rect 15142 16554 15148 16556
rect 13629 16552 15148 16554
rect 13629 16496 13634 16552
rect 13690 16496 15148 16552
rect 13629 16494 15148 16496
rect 13629 16491 13695 16494
rect 15142 16492 15148 16494
rect 15212 16492 15218 16556
rect 19374 16492 19380 16556
rect 19444 16554 19450 16556
rect 20253 16554 20319 16557
rect 19444 16552 20319 16554
rect 19444 16496 20258 16552
rect 20314 16496 20319 16552
rect 19444 16494 20319 16496
rect 28950 16554 29010 16630
rect 33174 16628 33180 16692
rect 33244 16690 33250 16692
rect 33961 16690 34027 16693
rect 33244 16688 34027 16690
rect 33244 16632 33966 16688
rect 34022 16632 34027 16688
rect 33244 16630 34027 16632
rect 33244 16628 33250 16630
rect 33961 16627 34027 16630
rect 33777 16556 33843 16557
rect 28950 16494 31770 16554
rect 19444 16492 19450 16494
rect 20253 16491 20319 16494
rect 9990 16356 9996 16420
rect 10060 16418 10066 16420
rect 10225 16418 10291 16421
rect 15377 16418 15443 16421
rect 10060 16416 15443 16418
rect 10060 16360 10230 16416
rect 10286 16360 15382 16416
rect 15438 16360 15443 16416
rect 10060 16358 15443 16360
rect 31710 16418 31770 16494
rect 33726 16492 33732 16556
rect 33796 16554 33843 16556
rect 33796 16552 33888 16554
rect 33838 16496 33888 16552
rect 33796 16494 33888 16496
rect 33796 16492 33843 16494
rect 33777 16491 33843 16492
rect 38469 16418 38535 16421
rect 31710 16416 38535 16418
rect 31710 16360 38474 16416
rect 38530 16360 38535 16416
rect 31710 16358 38535 16360
rect 10060 16356 10066 16358
rect 10225 16355 10291 16358
rect 15377 16355 15443 16358
rect 38469 16355 38535 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 24117 16284 24183 16285
rect 24117 16282 24164 16284
rect 24072 16280 24164 16282
rect 24072 16224 24122 16280
rect 24072 16222 24164 16224
rect 24117 16220 24164 16222
rect 24228 16220 24234 16284
rect 24117 16219 24183 16220
rect 11421 16146 11487 16149
rect 12985 16146 13051 16149
rect 11421 16144 13051 16146
rect 11421 16088 11426 16144
rect 11482 16088 12990 16144
rect 13046 16088 13051 16144
rect 11421 16086 13051 16088
rect 11421 16083 11487 16086
rect 12985 16083 13051 16086
rect 19425 16146 19491 16149
rect 20253 16146 20319 16149
rect 19425 16144 20319 16146
rect 19425 16088 19430 16144
rect 19486 16088 20258 16144
rect 20314 16088 20319 16144
rect 19425 16086 20319 16088
rect 19425 16083 19491 16086
rect 20253 16083 20319 16086
rect 10133 16010 10199 16013
rect 10910 16010 10916 16012
rect 10133 16008 10916 16010
rect 10133 15952 10138 16008
rect 10194 15952 10916 16008
rect 10133 15950 10916 15952
rect 10133 15947 10199 15950
rect 10910 15948 10916 15950
rect 10980 15948 10986 16012
rect 12750 15948 12756 16012
rect 12820 16010 12826 16012
rect 16849 16010 16915 16013
rect 12820 16008 16915 16010
rect 12820 15952 16854 16008
rect 16910 15952 16915 16008
rect 12820 15950 16915 15952
rect 12820 15948 12826 15950
rect 16849 15947 16915 15950
rect 23105 15874 23171 15877
rect 28349 15874 28415 15877
rect 30281 15874 30347 15877
rect 23105 15872 30347 15874
rect 23105 15816 23110 15872
rect 23166 15816 28354 15872
rect 28410 15816 30286 15872
rect 30342 15816 30347 15872
rect 23105 15814 30347 15816
rect 23105 15811 23171 15814
rect 28349 15811 28415 15814
rect 30281 15811 30347 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 20345 15738 20411 15741
rect 20897 15738 20963 15741
rect 20345 15736 20963 15738
rect 20345 15680 20350 15736
rect 20406 15680 20902 15736
rect 20958 15680 20963 15736
rect 20345 15678 20963 15680
rect 20345 15675 20411 15678
rect 20897 15675 20963 15678
rect 21081 15738 21147 15741
rect 27521 15738 27587 15741
rect 21081 15736 27587 15738
rect 21081 15680 21086 15736
rect 21142 15680 27526 15736
rect 27582 15680 27587 15736
rect 21081 15678 27587 15680
rect 21081 15675 21147 15678
rect 27521 15675 27587 15678
rect 28390 15676 28396 15740
rect 28460 15738 28466 15740
rect 31017 15738 31083 15741
rect 32070 15738 32076 15740
rect 28460 15736 32076 15738
rect 28460 15680 31022 15736
rect 31078 15680 32076 15736
rect 28460 15678 32076 15680
rect 28460 15676 28466 15678
rect 31017 15675 31083 15678
rect 32070 15676 32076 15678
rect 32140 15676 32146 15740
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 4981 15602 5047 15605
rect 4981 15600 22110 15602
rect 4981 15544 4986 15600
rect 5042 15544 22110 15600
rect 4981 15542 22110 15544
rect 4981 15539 5047 15542
rect 11329 15466 11395 15469
rect 13670 15466 13676 15468
rect 11329 15464 13676 15466
rect 11329 15408 11334 15464
rect 11390 15408 13676 15464
rect 11329 15406 13676 15408
rect 11329 15403 11395 15406
rect 13670 15404 13676 15406
rect 13740 15466 13746 15468
rect 21081 15466 21147 15469
rect 13740 15464 21147 15466
rect 13740 15408 21086 15464
rect 21142 15408 21147 15464
rect 13740 15406 21147 15408
rect 22050 15466 22110 15542
rect 23054 15540 23060 15604
rect 23124 15602 23130 15604
rect 24025 15602 24091 15605
rect 23124 15600 24091 15602
rect 23124 15544 24030 15600
rect 24086 15544 24091 15600
rect 23124 15542 24091 15544
rect 23124 15540 23130 15542
rect 24025 15539 24091 15542
rect 24853 15602 24919 15605
rect 36629 15602 36695 15605
rect 24853 15600 36695 15602
rect 24853 15544 24858 15600
rect 24914 15544 36634 15600
rect 36690 15544 36695 15600
rect 24853 15542 36695 15544
rect 24853 15539 24919 15542
rect 36629 15539 36695 15542
rect 37273 15466 37339 15469
rect 22050 15464 37339 15466
rect 22050 15408 37278 15464
rect 37334 15408 37339 15464
rect 22050 15406 37339 15408
rect 13740 15404 13746 15406
rect 21081 15403 21147 15406
rect 37273 15403 37339 15406
rect 16205 15332 16271 15333
rect 16205 15328 16252 15332
rect 16316 15330 16322 15332
rect 18413 15330 18479 15333
rect 18873 15330 18939 15333
rect 16205 15272 16210 15328
rect 16205 15268 16252 15272
rect 16316 15270 16362 15330
rect 18413 15328 18939 15330
rect 18413 15272 18418 15328
rect 18474 15272 18878 15328
rect 18934 15272 18939 15328
rect 18413 15270 18939 15272
rect 16316 15268 16322 15270
rect 16205 15267 16271 15268
rect 18413 15267 18479 15270
rect 18873 15267 18939 15270
rect 24526 15268 24532 15332
rect 24596 15330 24602 15332
rect 24669 15330 24735 15333
rect 24596 15328 24735 15330
rect 24596 15272 24674 15328
rect 24730 15272 24735 15328
rect 24596 15270 24735 15272
rect 24596 15268 24602 15270
rect 24669 15267 24735 15270
rect 28942 15268 28948 15332
rect 29012 15330 29018 15332
rect 29729 15330 29795 15333
rect 29012 15328 29795 15330
rect 29012 15272 29734 15328
rect 29790 15272 29795 15328
rect 29012 15270 29795 15272
rect 29012 15268 29018 15270
rect 29729 15267 29795 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 8017 15194 8083 15197
rect 13118 15194 13124 15196
rect 8017 15192 13124 15194
rect 8017 15136 8022 15192
rect 8078 15136 13124 15192
rect 8017 15134 13124 15136
rect 8017 15131 8083 15134
rect 13118 15132 13124 15134
rect 13188 15194 13194 15196
rect 13486 15194 13492 15196
rect 13188 15134 13492 15194
rect 13188 15132 13194 15134
rect 13486 15132 13492 15134
rect 13556 15132 13562 15196
rect 28073 15192 28139 15197
rect 28073 15136 28078 15192
rect 28134 15136 28139 15192
rect 28073 15131 28139 15136
rect 200 15058 800 15088
rect 1669 15058 1735 15061
rect 200 15056 1735 15058
rect 200 15000 1674 15056
rect 1730 15000 1735 15056
rect 200 14998 1735 15000
rect 200 14968 800 14998
rect 1669 14995 1735 14998
rect 6494 14996 6500 15060
rect 6564 15058 6570 15060
rect 9949 15058 10015 15061
rect 6564 15056 10015 15058
rect 6564 15000 9954 15056
rect 10010 15000 10015 15056
rect 6564 14998 10015 15000
rect 6564 14996 6570 14998
rect 9949 14995 10015 14998
rect 19057 15058 19123 15061
rect 21766 15058 21772 15060
rect 19057 15056 21772 15058
rect 19057 15000 19062 15056
rect 19118 15000 21772 15056
rect 19057 14998 21772 15000
rect 19057 14995 19123 14998
rect 21766 14996 21772 14998
rect 21836 14996 21842 15060
rect 9765 14924 9831 14925
rect 9765 14922 9812 14924
rect 9720 14920 9812 14922
rect 9720 14864 9770 14920
rect 9720 14862 9812 14864
rect 9765 14860 9812 14862
rect 9876 14860 9882 14924
rect 12893 14922 12959 14925
rect 24209 14922 24275 14925
rect 12893 14920 24275 14922
rect 12893 14864 12898 14920
rect 12954 14864 24214 14920
rect 24270 14864 24275 14920
rect 12893 14862 24275 14864
rect 9765 14859 9831 14860
rect 12893 14859 12959 14862
rect 24209 14859 24275 14862
rect 16798 14724 16804 14788
rect 16868 14786 16874 14788
rect 17033 14786 17099 14789
rect 16868 14784 17099 14786
rect 16868 14728 17038 14784
rect 17094 14728 17099 14784
rect 16868 14726 17099 14728
rect 16868 14724 16874 14726
rect 17033 14723 17099 14726
rect 19425 14786 19491 14789
rect 28076 14786 28136 15131
rect 38193 15058 38259 15061
rect 39200 15058 39800 15088
rect 38193 15056 39800 15058
rect 38193 15000 38198 15056
rect 38254 15000 39800 15056
rect 38193 14998 39800 15000
rect 38193 14995 38259 14998
rect 39200 14968 39800 14998
rect 19425 14784 28136 14786
rect 19425 14728 19430 14784
rect 19486 14728 28136 14784
rect 19425 14726 28136 14728
rect 19425 14723 19491 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 33174 14650 33180 14652
rect 22050 14590 33180 14650
rect 12893 14514 12959 14517
rect 14457 14514 14523 14517
rect 12893 14512 14523 14514
rect 12893 14456 12898 14512
rect 12954 14456 14462 14512
rect 14518 14456 14523 14512
rect 12893 14454 14523 14456
rect 12893 14451 12959 14454
rect 14457 14451 14523 14454
rect 17718 14452 17724 14516
rect 17788 14514 17794 14516
rect 22050 14514 22110 14590
rect 33174 14588 33180 14590
rect 33244 14588 33250 14652
rect 17788 14454 22110 14514
rect 17788 14452 17794 14454
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 27337 14378 27403 14381
rect 27470 14378 27476 14380
rect 27337 14376 27476 14378
rect 27337 14320 27342 14376
rect 27398 14320 27476 14376
rect 27337 14318 27476 14320
rect 27337 14315 27403 14318
rect 27470 14316 27476 14318
rect 27540 14316 27546 14380
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 12893 14242 12959 14245
rect 13261 14242 13327 14245
rect 12893 14240 13327 14242
rect 12893 14184 12898 14240
rect 12954 14184 13266 14240
rect 13322 14184 13327 14240
rect 12893 14182 13327 14184
rect 12893 14179 12959 14182
rect 13261 14179 13327 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 20621 14106 20687 14109
rect 20846 14106 20852 14108
rect 20621 14104 20852 14106
rect 20621 14048 20626 14104
rect 20682 14048 20852 14104
rect 20621 14046 20852 14048
rect 20621 14043 20687 14046
rect 20846 14044 20852 14046
rect 20916 14044 20922 14108
rect 8845 13970 8911 13973
rect 14406 13970 14412 13972
rect 8845 13968 14412 13970
rect 8845 13912 8850 13968
rect 8906 13912 14412 13968
rect 8845 13910 14412 13912
rect 8845 13907 8911 13910
rect 14406 13908 14412 13910
rect 14476 13908 14482 13972
rect 19333 13970 19399 13973
rect 20713 13970 20779 13973
rect 19333 13968 20779 13970
rect 19333 13912 19338 13968
rect 19394 13912 20718 13968
rect 20774 13912 20779 13968
rect 19333 13910 20779 13912
rect 19333 13907 19399 13910
rect 20713 13907 20779 13910
rect 1853 13834 1919 13837
rect 19609 13834 19675 13837
rect 20805 13834 20871 13837
rect 1853 13832 6930 13834
rect 1853 13776 1858 13832
rect 1914 13776 6930 13832
rect 1853 13774 6930 13776
rect 1853 13771 1919 13774
rect 5073 13698 5139 13701
rect 5206 13698 5212 13700
rect 5073 13696 5212 13698
rect 5073 13640 5078 13696
rect 5134 13640 5212 13696
rect 5073 13638 5212 13640
rect 5073 13635 5139 13638
rect 5206 13636 5212 13638
rect 5276 13636 5282 13700
rect 6870 13698 6930 13774
rect 19609 13832 20871 13834
rect 19609 13776 19614 13832
rect 19670 13776 20810 13832
rect 20866 13776 20871 13832
rect 19609 13774 20871 13776
rect 19609 13771 19675 13774
rect 20805 13771 20871 13774
rect 9070 13698 9076 13700
rect 6870 13638 9076 13698
rect 9070 13636 9076 13638
rect 9140 13636 9146 13700
rect 16297 13698 16363 13701
rect 16941 13698 17007 13701
rect 17401 13700 17467 13701
rect 16297 13696 17007 13698
rect 16297 13640 16302 13696
rect 16358 13640 16946 13696
rect 17002 13640 17007 13696
rect 16297 13638 17007 13640
rect 16297 13635 16363 13638
rect 16941 13635 17007 13638
rect 17350 13636 17356 13700
rect 17420 13698 17467 13700
rect 17420 13696 17512 13698
rect 17462 13640 17512 13696
rect 17420 13638 17512 13640
rect 17420 13636 17467 13638
rect 20294 13636 20300 13700
rect 20364 13698 20370 13700
rect 20989 13698 21055 13701
rect 20364 13696 21055 13698
rect 20364 13640 20994 13696
rect 21050 13640 21055 13696
rect 20364 13638 21055 13640
rect 20364 13636 20370 13638
rect 17358 13635 17467 13636
rect 20989 13635 21055 13638
rect 27654 13636 27660 13700
rect 27724 13698 27730 13700
rect 28257 13698 28323 13701
rect 27724 13696 28323 13698
rect 27724 13640 28262 13696
rect 28318 13640 28323 13696
rect 27724 13638 28323 13640
rect 27724 13636 27730 13638
rect 28257 13635 28323 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 13629 13564 13695 13565
rect 13629 13562 13676 13564
rect 13584 13560 13676 13562
rect 13740 13562 13746 13564
rect 14222 13562 14228 13564
rect 13584 13504 13634 13560
rect 13584 13502 13676 13504
rect 13629 13500 13676 13502
rect 13740 13502 14228 13562
rect 13740 13500 13746 13502
rect 14222 13500 14228 13502
rect 14292 13500 14298 13564
rect 16614 13500 16620 13564
rect 16684 13562 16690 13564
rect 17358 13562 17418 13635
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 16684 13502 17418 13562
rect 20713 13562 20779 13565
rect 22870 13562 22876 13564
rect 20713 13560 22876 13562
rect 20713 13504 20718 13560
rect 20774 13504 22876 13560
rect 20713 13502 22876 13504
rect 16684 13500 16690 13502
rect 13629 13499 13695 13500
rect 20713 13499 20779 13502
rect 22870 13500 22876 13502
rect 22940 13500 22946 13564
rect 11053 13426 11119 13429
rect 12198 13426 12204 13428
rect 11053 13424 12204 13426
rect 11053 13368 11058 13424
rect 11114 13368 12204 13424
rect 11053 13366 12204 13368
rect 11053 13363 11119 13366
rect 12198 13364 12204 13366
rect 12268 13364 12274 13428
rect 23054 13426 23060 13428
rect 12390 13366 23060 13426
rect 7046 13228 7052 13292
rect 7116 13290 7122 13292
rect 9121 13290 9187 13293
rect 12390 13290 12450 13366
rect 23054 13364 23060 13366
rect 23124 13364 23130 13428
rect 7116 13288 12450 13290
rect 7116 13232 9126 13288
rect 9182 13232 12450 13288
rect 7116 13230 12450 13232
rect 14825 13290 14891 13293
rect 15561 13290 15627 13293
rect 18781 13290 18847 13293
rect 14825 13288 15394 13290
rect 14825 13232 14830 13288
rect 14886 13232 15394 13288
rect 14825 13230 15394 13232
rect 7116 13228 7122 13230
rect 9121 13227 9187 13230
rect 14825 13227 14891 13230
rect 15334 13154 15394 13230
rect 15561 13288 18847 13290
rect 15561 13232 15566 13288
rect 15622 13232 18786 13288
rect 18842 13232 18847 13288
rect 15561 13230 18847 13232
rect 15561 13227 15627 13230
rect 18781 13227 18847 13230
rect 20110 13228 20116 13292
rect 20180 13290 20186 13292
rect 20897 13290 20963 13293
rect 20180 13288 20963 13290
rect 20180 13232 20902 13288
rect 20958 13232 20963 13288
rect 20180 13230 20963 13232
rect 20180 13228 20186 13230
rect 20897 13227 20963 13230
rect 17902 13154 17908 13156
rect 15334 13094 17908 13154
rect 17902 13092 17908 13094
rect 17972 13092 17978 13156
rect 20529 13154 20595 13157
rect 20713 13154 20779 13157
rect 20529 13152 20779 13154
rect 20529 13096 20534 13152
rect 20590 13096 20718 13152
rect 20774 13096 20779 13152
rect 20529 13094 20779 13096
rect 20529 13091 20595 13094
rect 20713 13091 20779 13094
rect 30782 13092 30788 13156
rect 30852 13154 30858 13156
rect 34237 13154 34303 13157
rect 30852 13152 34303 13154
rect 30852 13096 34242 13152
rect 34298 13096 34303 13152
rect 30852 13094 34303 13096
rect 30852 13092 30858 13094
rect 34237 13091 34303 13094
rect 19570 13088 19886 13089
rect 200 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 1577 13018 1643 13021
rect 200 13016 1643 13018
rect 200 12960 1582 13016
rect 1638 12960 1643 13016
rect 200 12958 1643 12960
rect 200 12928 800 12958
rect 1577 12955 1643 12958
rect 22502 12956 22508 13020
rect 22572 13018 22578 13020
rect 32949 13018 33015 13021
rect 22572 13016 33015 13018
rect 22572 12960 32954 13016
rect 33010 12960 33015 13016
rect 22572 12958 33015 12960
rect 22572 12956 22578 12958
rect 32949 12955 33015 12958
rect 38285 13018 38351 13021
rect 39200 13018 39800 13048
rect 38285 13016 39800 13018
rect 38285 12960 38290 13016
rect 38346 12960 39800 13016
rect 38285 12958 39800 12960
rect 38285 12955 38351 12958
rect 39200 12928 39800 12958
rect 9121 12884 9187 12885
rect 9070 12820 9076 12884
rect 9140 12882 9187 12884
rect 12433 12882 12499 12885
rect 13077 12882 13143 12885
rect 9140 12880 9232 12882
rect 9182 12824 9232 12880
rect 9140 12822 9232 12824
rect 12433 12880 13143 12882
rect 12433 12824 12438 12880
rect 12494 12824 13082 12880
rect 13138 12824 13143 12880
rect 12433 12822 13143 12824
rect 9140 12820 9187 12822
rect 9121 12819 9187 12820
rect 12433 12819 12499 12822
rect 13077 12819 13143 12822
rect 16389 12882 16455 12885
rect 22134 12882 22140 12884
rect 16389 12880 22140 12882
rect 16389 12824 16394 12880
rect 16450 12824 22140 12880
rect 16389 12822 22140 12824
rect 16389 12819 16455 12822
rect 22134 12820 22140 12822
rect 22204 12820 22210 12884
rect 28349 12882 28415 12885
rect 33317 12882 33383 12885
rect 28349 12880 33383 12882
rect 28349 12824 28354 12880
rect 28410 12824 33322 12880
rect 33378 12824 33383 12880
rect 28349 12822 33383 12824
rect 28349 12819 28415 12822
rect 33317 12819 33383 12822
rect 34513 12882 34579 12885
rect 35750 12882 35756 12884
rect 34513 12880 35756 12882
rect 34513 12824 34518 12880
rect 34574 12824 35756 12880
rect 34513 12822 35756 12824
rect 34513 12819 34579 12822
rect 35750 12820 35756 12822
rect 35820 12820 35826 12884
rect 11697 12746 11763 12749
rect 19149 12746 19215 12749
rect 11697 12744 19215 12746
rect 11697 12688 11702 12744
rect 11758 12688 19154 12744
rect 19210 12688 19215 12744
rect 11697 12686 19215 12688
rect 11697 12683 11763 12686
rect 19149 12683 19215 12686
rect 19333 12746 19399 12749
rect 20529 12746 20595 12749
rect 19333 12744 20595 12746
rect 19333 12688 19338 12744
rect 19394 12688 20534 12744
rect 20590 12688 20595 12744
rect 19333 12686 20595 12688
rect 19333 12683 19399 12686
rect 20529 12683 20595 12686
rect 24894 12684 24900 12748
rect 24964 12746 24970 12748
rect 38193 12746 38259 12749
rect 24964 12744 38259 12746
rect 24964 12688 38198 12744
rect 38254 12688 38259 12744
rect 24964 12686 38259 12688
rect 24964 12684 24970 12686
rect 38193 12683 38259 12686
rect 11513 12610 11579 12613
rect 12893 12610 12959 12613
rect 20069 12610 20135 12613
rect 20345 12612 20411 12613
rect 11513 12608 12959 12610
rect 11513 12552 11518 12608
rect 11574 12552 12898 12608
rect 12954 12552 12959 12608
rect 11513 12550 12959 12552
rect 11513 12547 11579 12550
rect 12893 12547 12959 12550
rect 19566 12608 20135 12610
rect 19566 12552 20074 12608
rect 20130 12552 20135 12608
rect 19566 12550 20135 12552
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 2262 12412 2268 12476
rect 2332 12474 2338 12476
rect 4061 12474 4127 12477
rect 2332 12472 4127 12474
rect 2332 12416 4066 12472
rect 4122 12416 4127 12472
rect 2332 12414 4127 12416
rect 2332 12412 2338 12414
rect 4061 12411 4127 12414
rect 6678 12412 6684 12476
rect 6748 12474 6754 12476
rect 9990 12474 9996 12476
rect 6748 12414 9996 12474
rect 6748 12412 6754 12414
rect 9990 12412 9996 12414
rect 10060 12412 10066 12476
rect 10501 12474 10567 12477
rect 14825 12474 14891 12477
rect 10501 12472 14891 12474
rect 10501 12416 10506 12472
rect 10562 12416 14830 12472
rect 14886 12416 14891 12472
rect 10501 12414 14891 12416
rect 10501 12411 10567 12414
rect 14825 12411 14891 12414
rect 19425 12474 19491 12477
rect 19566 12474 19626 12550
rect 20069 12547 20135 12550
rect 20294 12548 20300 12612
rect 20364 12610 20411 12612
rect 20364 12608 20456 12610
rect 20406 12552 20456 12608
rect 20364 12550 20456 12552
rect 20364 12548 20411 12550
rect 22134 12548 22140 12612
rect 22204 12610 22210 12612
rect 22369 12610 22435 12613
rect 22204 12608 22435 12610
rect 22204 12552 22374 12608
rect 22430 12552 22435 12608
rect 22204 12550 22435 12552
rect 22204 12548 22210 12550
rect 20345 12547 20411 12548
rect 22369 12547 22435 12550
rect 29637 12610 29703 12613
rect 32254 12610 32260 12612
rect 29637 12608 32260 12610
rect 29637 12552 29642 12608
rect 29698 12552 32260 12608
rect 29637 12550 32260 12552
rect 29637 12547 29703 12550
rect 32254 12548 32260 12550
rect 32324 12548 32330 12612
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19425 12472 19626 12474
rect 19425 12416 19430 12472
rect 19486 12416 19626 12472
rect 19425 12414 19626 12416
rect 20069 12474 20135 12477
rect 20437 12474 20503 12477
rect 20069 12472 20503 12474
rect 20069 12416 20074 12472
rect 20130 12416 20442 12472
rect 20498 12416 20503 12472
rect 20069 12414 20503 12416
rect 19425 12411 19491 12414
rect 20069 12411 20135 12414
rect 20437 12411 20503 12414
rect 21633 12474 21699 12477
rect 23933 12474 23999 12477
rect 28625 12476 28691 12477
rect 21633 12472 23999 12474
rect 21633 12416 21638 12472
rect 21694 12416 23938 12472
rect 23994 12416 23999 12472
rect 21633 12414 23999 12416
rect 21633 12411 21699 12414
rect 23933 12411 23999 12414
rect 28574 12412 28580 12476
rect 28644 12474 28691 12476
rect 32438 12474 32444 12476
rect 28644 12472 28736 12474
rect 28686 12416 28736 12472
rect 28644 12414 28736 12416
rect 29318 12414 32444 12474
rect 28644 12412 28691 12414
rect 28625 12411 28691 12412
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 1894 12276 1900 12340
rect 1964 12338 1970 12340
rect 3877 12338 3943 12341
rect 1964 12336 3943 12338
rect 1964 12280 3882 12336
rect 3938 12280 3943 12336
rect 1964 12278 3943 12280
rect 1964 12276 1970 12278
rect 3877 12275 3943 12278
rect 9673 12338 9739 12341
rect 10225 12338 10291 12341
rect 9673 12336 10291 12338
rect 9673 12280 9678 12336
rect 9734 12280 10230 12336
rect 10286 12280 10291 12336
rect 9673 12278 10291 12280
rect 9673 12275 9739 12278
rect 10225 12275 10291 12278
rect 11697 12338 11763 12341
rect 13353 12338 13419 12341
rect 11697 12336 13419 12338
rect 11697 12280 11702 12336
rect 11758 12280 13358 12336
rect 13414 12280 13419 12336
rect 11697 12278 13419 12280
rect 11697 12275 11763 12278
rect 13353 12275 13419 12278
rect 13629 12338 13695 12341
rect 18454 12338 18460 12340
rect 13629 12336 18460 12338
rect 13629 12280 13634 12336
rect 13690 12280 18460 12336
rect 13629 12278 18460 12280
rect 13629 12275 13695 12278
rect 18454 12276 18460 12278
rect 18524 12276 18530 12340
rect 19885 12338 19951 12341
rect 21541 12338 21607 12341
rect 25313 12340 25379 12341
rect 25262 12338 25268 12340
rect 19885 12336 20546 12338
rect 19885 12280 19890 12336
rect 19946 12280 20546 12336
rect 19885 12278 20546 12280
rect 19885 12275 19951 12278
rect 20486 12205 20546 12278
rect 21541 12336 25268 12338
rect 25332 12338 25379 12340
rect 25957 12338 26023 12341
rect 29318 12340 29378 12414
rect 32438 12412 32444 12414
rect 32508 12412 32514 12476
rect 27470 12338 27476 12340
rect 25332 12336 25424 12338
rect 21541 12280 21546 12336
rect 21602 12280 25268 12336
rect 25374 12280 25424 12336
rect 21541 12278 25268 12280
rect 21541 12275 21607 12278
rect 25262 12276 25268 12278
rect 25332 12278 25424 12280
rect 25957 12336 27476 12338
rect 25957 12280 25962 12336
rect 26018 12280 27476 12336
rect 25957 12278 27476 12280
rect 25332 12276 25379 12278
rect 25313 12275 25379 12276
rect 25957 12275 26023 12278
rect 27470 12276 27476 12278
rect 27540 12276 27546 12340
rect 29310 12276 29316 12340
rect 29380 12276 29386 12340
rect 38101 12338 38167 12341
rect 39200 12338 39800 12368
rect 38101 12336 39800 12338
rect 38101 12280 38106 12336
rect 38162 12280 39800 12336
rect 38101 12278 39800 12280
rect 38101 12275 38167 12278
rect 39200 12248 39800 12278
rect 9673 12202 9739 12205
rect 9673 12200 9874 12202
rect 9673 12144 9678 12200
rect 9734 12144 9874 12200
rect 9673 12142 9874 12144
rect 9673 12139 9739 12142
rect 9438 12004 9444 12068
rect 9508 12066 9514 12068
rect 9814 12066 9874 12142
rect 11830 12140 11836 12204
rect 11900 12202 11906 12204
rect 11973 12202 12039 12205
rect 11900 12200 12039 12202
rect 11900 12144 11978 12200
rect 12034 12144 12039 12200
rect 11900 12142 12039 12144
rect 11900 12140 11906 12142
rect 11973 12139 12039 12142
rect 18270 12140 18276 12204
rect 18340 12202 18346 12204
rect 20253 12202 20319 12205
rect 18340 12200 20319 12202
rect 18340 12144 20258 12200
rect 20314 12144 20319 12200
rect 18340 12142 20319 12144
rect 20486 12200 20595 12205
rect 20486 12144 20534 12200
rect 20590 12144 20595 12200
rect 20486 12142 20595 12144
rect 18340 12140 18346 12142
rect 20253 12139 20319 12142
rect 20529 12139 20595 12142
rect 24577 12202 24643 12205
rect 27613 12202 27679 12205
rect 24577 12200 27679 12202
rect 24577 12144 24582 12200
rect 24638 12144 27618 12200
rect 27674 12144 27679 12200
rect 24577 12142 27679 12144
rect 24577 12139 24643 12142
rect 27613 12139 27679 12142
rect 29269 12202 29335 12205
rect 31518 12202 31524 12204
rect 29269 12200 31524 12202
rect 29269 12144 29274 12200
rect 29330 12144 31524 12200
rect 29269 12142 31524 12144
rect 29269 12139 29335 12142
rect 31518 12140 31524 12142
rect 31588 12202 31594 12204
rect 35893 12202 35959 12205
rect 31588 12200 35959 12202
rect 31588 12144 35898 12200
rect 35954 12144 35959 12200
rect 31588 12142 35959 12144
rect 31588 12140 31594 12142
rect 35893 12139 35959 12142
rect 11053 12066 11119 12069
rect 17125 12066 17191 12069
rect 9508 12006 9690 12066
rect 9814 12064 17191 12066
rect 9814 12008 11058 12064
rect 11114 12008 17130 12064
rect 17186 12008 17191 12064
rect 9814 12006 17191 12008
rect 9508 12004 9514 12006
rect 8477 11930 8543 11933
rect 9305 11932 9371 11933
rect 9254 11930 9260 11932
rect 8477 11928 9260 11930
rect 9324 11928 9371 11932
rect 8477 11872 8482 11928
rect 8538 11872 9260 11928
rect 9366 11872 9371 11928
rect 8477 11870 9260 11872
rect 8477 11867 8543 11870
rect 9254 11868 9260 11870
rect 9324 11868 9371 11872
rect 9305 11867 9371 11868
rect 7189 11794 7255 11797
rect 9489 11794 9555 11797
rect 7189 11792 9555 11794
rect 7189 11736 7194 11792
rect 7250 11736 9494 11792
rect 9550 11736 9555 11792
rect 7189 11734 9555 11736
rect 9630 11794 9690 12006
rect 11053 12003 11119 12006
rect 17125 12003 17191 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 11697 11930 11763 11933
rect 14733 11930 14799 11933
rect 16481 11930 16547 11933
rect 11697 11928 16547 11930
rect 11697 11872 11702 11928
rect 11758 11872 14738 11928
rect 14794 11872 16486 11928
rect 16542 11872 16547 11928
rect 11697 11870 16547 11872
rect 11697 11867 11763 11870
rect 14733 11867 14799 11870
rect 16481 11867 16547 11870
rect 22553 11794 22619 11797
rect 22686 11794 22692 11796
rect 9630 11734 11346 11794
rect 7189 11731 7255 11734
rect 9489 11731 9555 11734
rect 6177 11658 6243 11661
rect 8702 11658 8708 11660
rect 6177 11656 8708 11658
rect 6177 11600 6182 11656
rect 6238 11600 8708 11656
rect 6177 11598 8708 11600
rect 6177 11595 6243 11598
rect 8702 11596 8708 11598
rect 8772 11596 8778 11660
rect 9806 11596 9812 11660
rect 9876 11658 9882 11660
rect 10133 11658 10199 11661
rect 10593 11660 10659 11661
rect 10542 11658 10548 11660
rect 9876 11656 10199 11658
rect 9876 11600 10138 11656
rect 10194 11600 10199 11656
rect 9876 11598 10199 11600
rect 10502 11598 10548 11658
rect 10612 11656 10659 11660
rect 10654 11600 10659 11656
rect 9876 11596 9882 11598
rect 10133 11595 10199 11598
rect 10542 11596 10548 11598
rect 10612 11596 10659 11600
rect 11286 11658 11346 11734
rect 22553 11792 22692 11794
rect 22553 11736 22558 11792
rect 22614 11736 22692 11792
rect 22553 11734 22692 11736
rect 22553 11731 22619 11734
rect 22686 11732 22692 11734
rect 22756 11732 22762 11796
rect 29913 11794 29979 11797
rect 30046 11794 30052 11796
rect 29913 11792 30052 11794
rect 29913 11736 29918 11792
rect 29974 11736 30052 11792
rect 29913 11734 30052 11736
rect 29913 11731 29979 11734
rect 30046 11732 30052 11734
rect 30116 11732 30122 11796
rect 12617 11658 12683 11661
rect 11286 11656 12683 11658
rect 11286 11600 12622 11656
rect 12678 11600 12683 11656
rect 11286 11598 12683 11600
rect 10593 11595 10659 11596
rect 12617 11595 12683 11598
rect 20621 11660 20687 11661
rect 20621 11656 20668 11660
rect 20732 11658 20738 11660
rect 20621 11600 20626 11656
rect 20621 11596 20668 11600
rect 20732 11598 20778 11658
rect 20732 11596 20738 11598
rect 26550 11596 26556 11660
rect 26620 11658 26626 11660
rect 28942 11658 28948 11660
rect 26620 11598 28948 11658
rect 26620 11596 26626 11598
rect 28942 11596 28948 11598
rect 29012 11596 29018 11660
rect 29453 11658 29519 11661
rect 30414 11658 30420 11660
rect 29453 11656 30420 11658
rect 29453 11600 29458 11656
rect 29514 11600 30420 11656
rect 29453 11598 30420 11600
rect 20621 11595 20687 11596
rect 29453 11595 29519 11598
rect 30414 11596 30420 11598
rect 30484 11596 30490 11660
rect 31518 11596 31524 11660
rect 31588 11658 31594 11660
rect 33685 11658 33751 11661
rect 31588 11656 33751 11658
rect 31588 11600 33690 11656
rect 33746 11600 33751 11656
rect 31588 11598 33751 11600
rect 31588 11596 31594 11598
rect 33685 11595 33751 11598
rect 5349 11522 5415 11525
rect 5349 11520 11346 11522
rect 5349 11464 5354 11520
rect 5410 11464 11346 11520
rect 5349 11462 11346 11464
rect 5349 11459 5415 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 7925 11386 7991 11389
rect 11053 11386 11119 11389
rect 7925 11384 11119 11386
rect 7925 11328 7930 11384
rect 7986 11328 11058 11384
rect 11114 11328 11119 11384
rect 7925 11326 11119 11328
rect 7925 11323 7991 11326
rect 11053 11323 11119 11326
rect 6637 11114 6703 11117
rect 10041 11116 10107 11117
rect 8334 11114 8340 11116
rect 6637 11112 8340 11114
rect 6637 11056 6642 11112
rect 6698 11056 8340 11112
rect 6637 11054 8340 11056
rect 6637 11051 6703 11054
rect 8334 11052 8340 11054
rect 8404 11052 8410 11116
rect 9990 11114 9996 11116
rect 9950 11054 9996 11114
rect 10060 11112 10107 11116
rect 10102 11056 10107 11112
rect 9990 11052 9996 11054
rect 10060 11052 10107 11056
rect 11286 11114 11346 11462
rect 18454 11460 18460 11524
rect 18524 11522 18530 11524
rect 22318 11522 22324 11524
rect 18524 11462 22324 11522
rect 18524 11460 18530 11462
rect 22318 11460 22324 11462
rect 22388 11460 22394 11524
rect 28073 11522 28139 11525
rect 28625 11522 28691 11525
rect 30741 11522 30807 11525
rect 28073 11520 30807 11522
rect 28073 11464 28078 11520
rect 28134 11464 28630 11520
rect 28686 11464 30746 11520
rect 30802 11464 30807 11520
rect 28073 11462 30807 11464
rect 28073 11459 28139 11462
rect 28625 11459 28691 11462
rect 30741 11459 30807 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 13905 11386 13971 11389
rect 15469 11386 15535 11389
rect 13905 11384 15535 11386
rect 13905 11328 13910 11384
rect 13966 11328 15474 11384
rect 15530 11328 15535 11384
rect 13905 11326 15535 11328
rect 13905 11323 13971 11326
rect 15469 11323 15535 11326
rect 26601 11386 26667 11389
rect 27981 11386 28047 11389
rect 26601 11384 28047 11386
rect 26601 11328 26606 11384
rect 26662 11328 27986 11384
rect 28042 11328 28047 11384
rect 26601 11326 28047 11328
rect 26601 11323 26667 11326
rect 27981 11323 28047 11326
rect 28165 11386 28231 11389
rect 29637 11386 29703 11389
rect 28165 11384 29703 11386
rect 28165 11328 28170 11384
rect 28226 11328 29642 11384
rect 29698 11328 29703 11384
rect 28165 11326 29703 11328
rect 28165 11323 28231 11326
rect 29637 11323 29703 11326
rect 14089 11250 14155 11253
rect 15469 11250 15535 11253
rect 14089 11248 15535 11250
rect 14089 11192 14094 11248
rect 14150 11192 15474 11248
rect 15530 11192 15535 11248
rect 14089 11190 15535 11192
rect 14089 11187 14155 11190
rect 15469 11187 15535 11190
rect 16757 11250 16823 11253
rect 18137 11250 18203 11253
rect 16757 11248 18203 11250
rect 16757 11192 16762 11248
rect 16818 11192 18142 11248
rect 18198 11192 18203 11248
rect 16757 11190 18203 11192
rect 16757 11187 16823 11190
rect 18137 11187 18203 11190
rect 20989 11250 21055 11253
rect 30465 11250 30531 11253
rect 37457 11250 37523 11253
rect 20989 11248 30531 11250
rect 20989 11192 20994 11248
rect 21050 11192 30470 11248
rect 30526 11192 30531 11248
rect 20989 11190 30531 11192
rect 20989 11187 21055 11190
rect 30465 11187 30531 11190
rect 31710 11248 37523 11250
rect 31710 11192 37462 11248
rect 37518 11192 37523 11248
rect 31710 11190 37523 11192
rect 16941 11114 17007 11117
rect 11286 11112 17007 11114
rect 11286 11056 16946 11112
rect 17002 11056 17007 11112
rect 11286 11054 17007 11056
rect 10041 11051 10107 11052
rect 16941 11051 17007 11054
rect 25497 11114 25563 11117
rect 26366 11114 26372 11116
rect 25497 11112 26372 11114
rect 25497 11056 25502 11112
rect 25558 11056 26372 11112
rect 25497 11054 26372 11056
rect 25497 11051 25563 11054
rect 26366 11052 26372 11054
rect 26436 11052 26442 11116
rect 31710 11114 31770 11190
rect 37457 11187 37523 11190
rect 27846 11054 31770 11114
rect 36077 11116 36143 11117
rect 36077 11112 36124 11116
rect 36188 11114 36194 11116
rect 36077 11056 36082 11112
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 6361 10978 6427 10981
rect 7741 10978 7807 10981
rect 6361 10976 7807 10978
rect 6361 10920 6366 10976
rect 6422 10920 7746 10976
rect 7802 10920 7807 10976
rect 6361 10918 7807 10920
rect 6361 10915 6427 10918
rect 7741 10915 7807 10918
rect 10225 10978 10291 10981
rect 12934 10978 12940 10980
rect 10225 10976 12940 10978
rect 10225 10920 10230 10976
rect 10286 10920 12940 10976
rect 10225 10918 12940 10920
rect 10225 10915 10291 10918
rect 12934 10916 12940 10918
rect 13004 10916 13010 10980
rect 14222 10916 14228 10980
rect 14292 10978 14298 10980
rect 14825 10978 14891 10981
rect 14292 10976 14891 10978
rect 14292 10920 14830 10976
rect 14886 10920 14891 10976
rect 14292 10918 14891 10920
rect 14292 10916 14298 10918
rect 14825 10915 14891 10918
rect 20437 10980 20503 10981
rect 20437 10976 20484 10980
rect 20548 10978 20554 10980
rect 27846 10978 27906 11054
rect 36077 11052 36124 11056
rect 36188 11054 36234 11114
rect 36188 11052 36194 11054
rect 36077 11051 36143 11052
rect 20437 10920 20442 10976
rect 20437 10916 20484 10920
rect 20548 10918 20594 10978
rect 22050 10918 27906 10978
rect 20548 10916 20554 10918
rect 20437 10915 20503 10916
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 5901 10842 5967 10845
rect 11329 10842 11395 10845
rect 5901 10840 11395 10842
rect 5901 10784 5906 10840
rect 5962 10784 11334 10840
rect 11390 10784 11395 10840
rect 5901 10782 11395 10784
rect 5901 10779 5967 10782
rect 11329 10779 11395 10782
rect 15878 10780 15884 10844
rect 15948 10842 15954 10844
rect 16430 10842 16436 10844
rect 15948 10782 16436 10842
rect 15948 10780 15954 10782
rect 16430 10780 16436 10782
rect 16500 10780 16506 10844
rect 22050 10842 22110 10918
rect 29126 10916 29132 10980
rect 29196 10978 29202 10980
rect 29453 10978 29519 10981
rect 29196 10976 29519 10978
rect 29196 10920 29458 10976
rect 29514 10920 29519 10976
rect 29196 10918 29519 10920
rect 29196 10916 29202 10918
rect 29453 10915 29519 10918
rect 30281 10978 30347 10981
rect 37365 10978 37431 10981
rect 30281 10976 37431 10978
rect 30281 10920 30286 10976
rect 30342 10920 37370 10976
rect 37426 10920 37431 10976
rect 30281 10918 37431 10920
rect 30281 10915 30347 10918
rect 37365 10915 37431 10918
rect 38101 10978 38167 10981
rect 39200 10978 39800 11008
rect 38101 10976 39800 10978
rect 38101 10920 38106 10976
rect 38162 10920 39800 10976
rect 38101 10918 39800 10920
rect 38101 10915 38167 10918
rect 39200 10888 39800 10918
rect 20072 10782 22110 10842
rect 28165 10842 28231 10845
rect 30741 10842 30807 10845
rect 31017 10842 31083 10845
rect 28165 10840 31083 10842
rect 28165 10784 28170 10840
rect 28226 10784 30746 10840
rect 30802 10784 31022 10840
rect 31078 10784 31083 10840
rect 28165 10782 31083 10784
rect 6913 10706 6979 10709
rect 8201 10706 8267 10709
rect 6913 10704 8267 10706
rect 6913 10648 6918 10704
rect 6974 10648 8206 10704
rect 8262 10648 8267 10704
rect 6913 10646 8267 10648
rect 6913 10643 6979 10646
rect 8201 10643 8267 10646
rect 9673 10706 9739 10709
rect 11094 10706 11100 10708
rect 9673 10704 11100 10706
rect 9673 10648 9678 10704
rect 9734 10648 11100 10704
rect 9673 10646 11100 10648
rect 9673 10643 9739 10646
rect 11094 10644 11100 10646
rect 11164 10644 11170 10708
rect 12617 10706 12683 10709
rect 13445 10706 13511 10709
rect 12617 10704 13511 10706
rect 12617 10648 12622 10704
rect 12678 10648 13450 10704
rect 13506 10648 13511 10704
rect 12617 10646 13511 10648
rect 12617 10643 12683 10646
rect 13445 10643 13511 10646
rect 16430 10644 16436 10708
rect 16500 10706 16506 10708
rect 20072 10706 20132 10782
rect 28165 10779 28231 10782
rect 30741 10779 30807 10782
rect 31017 10779 31083 10782
rect 20345 10708 20411 10709
rect 16500 10646 20132 10706
rect 16500 10644 16506 10646
rect 20294 10644 20300 10708
rect 20364 10706 20411 10708
rect 20713 10706 20779 10709
rect 21449 10706 21515 10709
rect 32029 10706 32095 10709
rect 20364 10704 20456 10706
rect 20406 10648 20456 10704
rect 20364 10646 20456 10648
rect 20713 10704 32095 10706
rect 20713 10648 20718 10704
rect 20774 10648 21454 10704
rect 21510 10648 32034 10704
rect 32090 10648 32095 10704
rect 20713 10646 32095 10648
rect 20364 10644 20411 10646
rect 20345 10643 20411 10644
rect 20713 10643 20779 10646
rect 21449 10643 21515 10646
rect 32029 10643 32095 10646
rect 10501 10570 10567 10573
rect 13813 10570 13879 10573
rect 10501 10568 13879 10570
rect 10501 10512 10506 10568
rect 10562 10512 13818 10568
rect 13874 10512 13879 10568
rect 10501 10510 13879 10512
rect 10501 10507 10567 10510
rect 13813 10507 13879 10510
rect 24577 10570 24643 10573
rect 25814 10570 25820 10572
rect 24577 10568 25820 10570
rect 24577 10512 24582 10568
rect 24638 10512 25820 10568
rect 24577 10510 25820 10512
rect 24577 10507 24643 10510
rect 25814 10508 25820 10510
rect 25884 10570 25890 10572
rect 26049 10570 26115 10573
rect 25884 10568 26115 10570
rect 25884 10512 26054 10568
rect 26110 10512 26115 10568
rect 25884 10510 26115 10512
rect 25884 10508 25890 10510
rect 26049 10507 26115 10510
rect 31017 10570 31083 10573
rect 31201 10570 31267 10573
rect 31017 10568 31267 10570
rect 31017 10512 31022 10568
rect 31078 10512 31206 10568
rect 31262 10512 31267 10568
rect 31017 10510 31267 10512
rect 31017 10507 31083 10510
rect 31201 10507 31267 10510
rect 9765 10434 9831 10437
rect 13997 10434 14063 10437
rect 9765 10432 14063 10434
rect 9765 10376 9770 10432
rect 9826 10376 14002 10432
rect 14058 10376 14063 10432
rect 9765 10374 14063 10376
rect 9765 10371 9831 10374
rect 13997 10371 14063 10374
rect 30833 10434 30899 10437
rect 31661 10434 31727 10437
rect 30833 10432 31727 10434
rect 30833 10376 30838 10432
rect 30894 10376 31666 10432
rect 31722 10376 31727 10432
rect 30833 10374 31727 10376
rect 30833 10371 30899 10374
rect 31661 10371 31727 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1761 10298 1827 10301
rect 200 10296 1827 10298
rect 200 10240 1766 10296
rect 1822 10240 1827 10296
rect 200 10238 1827 10240
rect 200 10208 800 10238
rect 1761 10235 1827 10238
rect 29085 10298 29151 10301
rect 32213 10298 32279 10301
rect 29085 10296 32279 10298
rect 29085 10240 29090 10296
rect 29146 10240 32218 10296
rect 32274 10240 32279 10296
rect 29085 10238 32279 10240
rect 29085 10235 29151 10238
rect 32213 10235 32279 10238
rect 38101 10298 38167 10301
rect 39200 10298 39800 10328
rect 38101 10296 39800 10298
rect 38101 10240 38106 10296
rect 38162 10240 39800 10296
rect 38101 10238 39800 10240
rect 38101 10235 38167 10238
rect 39200 10208 39800 10238
rect 4061 10162 4127 10165
rect 7465 10162 7531 10165
rect 4061 10160 7531 10162
rect 4061 10104 4066 10160
rect 4122 10104 7470 10160
rect 7526 10104 7531 10160
rect 4061 10102 7531 10104
rect 4061 10099 4127 10102
rect 7465 10099 7531 10102
rect 31477 10162 31543 10165
rect 33593 10162 33659 10165
rect 31477 10160 33659 10162
rect 31477 10104 31482 10160
rect 31538 10104 33598 10160
rect 33654 10104 33659 10160
rect 31477 10102 33659 10104
rect 31477 10099 31543 10102
rect 33593 10099 33659 10102
rect 5809 10028 5875 10029
rect 5758 9964 5764 10028
rect 5828 10026 5875 10028
rect 6729 10026 6795 10029
rect 7649 10026 7715 10029
rect 11973 10028 12039 10029
rect 11973 10026 12020 10028
rect 5828 10024 5920 10026
rect 5870 9968 5920 10024
rect 5828 9966 5920 9968
rect 6729 10024 7715 10026
rect 6729 9968 6734 10024
rect 6790 9968 7654 10024
rect 7710 9968 7715 10024
rect 6729 9966 7715 9968
rect 11928 10024 12020 10026
rect 11928 9968 11978 10024
rect 11928 9966 12020 9968
rect 5828 9964 5875 9966
rect 5809 9963 5875 9964
rect 6729 9963 6795 9966
rect 7649 9963 7715 9966
rect 11973 9964 12020 9966
rect 12084 9964 12090 10028
rect 16665 10026 16731 10029
rect 17585 10026 17651 10029
rect 35617 10026 35683 10029
rect 16665 10024 17651 10026
rect 16665 9968 16670 10024
rect 16726 9968 17590 10024
rect 17646 9968 17651 10024
rect 16665 9966 17651 9968
rect 11973 9963 12039 9964
rect 16665 9963 16731 9966
rect 17585 9963 17651 9966
rect 31710 10024 35683 10026
rect 31710 9968 35622 10024
rect 35678 9968 35683 10024
rect 31710 9966 35683 9968
rect 6269 9890 6335 9893
rect 8385 9890 8451 9893
rect 6269 9888 8451 9890
rect 6269 9832 6274 9888
rect 6330 9832 8390 9888
rect 8446 9832 8451 9888
rect 6269 9830 8451 9832
rect 6269 9827 6335 9830
rect 8385 9827 8451 9830
rect 12433 9890 12499 9893
rect 14089 9890 14155 9893
rect 19374 9890 19380 9892
rect 12433 9888 19380 9890
rect 12433 9832 12438 9888
rect 12494 9832 14094 9888
rect 14150 9832 19380 9888
rect 12433 9830 19380 9832
rect 12433 9827 12499 9830
rect 14089 9827 14155 9830
rect 19374 9828 19380 9830
rect 19444 9828 19450 9892
rect 20437 9890 20503 9893
rect 26785 9892 26851 9893
rect 20846 9890 20852 9892
rect 20437 9888 20852 9890
rect 20437 9832 20442 9888
rect 20498 9832 20852 9888
rect 20437 9830 20852 9832
rect 20437 9827 20503 9830
rect 20846 9828 20852 9830
rect 20916 9828 20922 9892
rect 26734 9890 26740 9892
rect 26694 9830 26740 9890
rect 26804 9888 26851 9892
rect 26846 9832 26851 9888
rect 26734 9828 26740 9830
rect 26804 9828 26851 9832
rect 28942 9828 28948 9892
rect 29012 9890 29018 9892
rect 30598 9890 30604 9892
rect 29012 9830 30604 9890
rect 29012 9828 29018 9830
rect 30598 9828 30604 9830
rect 30668 9890 30674 9892
rect 31569 9890 31635 9893
rect 30668 9888 31635 9890
rect 30668 9832 31574 9888
rect 31630 9832 31635 9888
rect 30668 9830 31635 9832
rect 30668 9828 30674 9830
rect 26785 9827 26851 9828
rect 31569 9827 31635 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 6453 9754 6519 9757
rect 9857 9754 9923 9757
rect 10726 9754 10732 9756
rect 6453 9752 6930 9754
rect 6453 9696 6458 9752
rect 6514 9696 6930 9752
rect 6453 9694 6930 9696
rect 6453 9691 6519 9694
rect 200 9618 800 9648
rect 1761 9618 1827 9621
rect 5901 9620 5967 9621
rect 5901 9618 5948 9620
rect 200 9616 1827 9618
rect 200 9560 1766 9616
rect 1822 9560 1827 9616
rect 200 9558 1827 9560
rect 5856 9616 5948 9618
rect 5856 9560 5906 9616
rect 5856 9558 5948 9560
rect 200 9528 800 9558
rect 1761 9555 1827 9558
rect 5901 9556 5948 9558
rect 6012 9556 6018 9620
rect 6361 9618 6427 9621
rect 6870 9620 6930 9694
rect 9857 9752 10732 9754
rect 9857 9696 9862 9752
rect 9918 9696 10732 9752
rect 9857 9694 10732 9696
rect 9857 9691 9923 9694
rect 10726 9692 10732 9694
rect 10796 9692 10802 9756
rect 16246 9692 16252 9756
rect 16316 9754 16322 9756
rect 18045 9754 18111 9757
rect 18597 9756 18663 9757
rect 18597 9754 18644 9756
rect 16316 9752 18111 9754
rect 16316 9696 18050 9752
rect 18106 9696 18111 9752
rect 16316 9694 18111 9696
rect 18552 9752 18644 9754
rect 18552 9696 18602 9752
rect 18552 9694 18644 9696
rect 16316 9692 16322 9694
rect 18045 9691 18111 9694
rect 18597 9692 18644 9694
rect 18708 9692 18714 9756
rect 26049 9754 26115 9757
rect 26918 9754 26924 9756
rect 26049 9752 26924 9754
rect 26049 9696 26054 9752
rect 26110 9696 26924 9752
rect 26049 9694 26924 9696
rect 18597 9691 18663 9692
rect 26049 9691 26115 9694
rect 26918 9692 26924 9694
rect 26988 9754 26994 9756
rect 27429 9754 27495 9757
rect 31710 9754 31770 9966
rect 35617 9963 35683 9966
rect 33317 9890 33383 9893
rect 34237 9890 34303 9893
rect 33317 9888 34303 9890
rect 33317 9832 33322 9888
rect 33378 9832 34242 9888
rect 34298 9832 34303 9888
rect 33317 9830 34303 9832
rect 33317 9827 33383 9830
rect 34237 9827 34303 9830
rect 26988 9752 31770 9754
rect 26988 9696 27434 9752
rect 27490 9696 31770 9752
rect 26988 9694 31770 9696
rect 26988 9692 26994 9694
rect 27429 9691 27495 9694
rect 6678 9618 6684 9620
rect 6361 9616 6684 9618
rect 6361 9560 6366 9616
rect 6422 9560 6684 9616
rect 6361 9558 6684 9560
rect 5901 9555 5967 9556
rect 6361 9555 6427 9558
rect 6678 9556 6684 9558
rect 6748 9556 6754 9620
rect 6862 9556 6868 9620
rect 6932 9556 6938 9620
rect 7925 9618 7991 9621
rect 10501 9620 10567 9621
rect 7925 9616 8034 9618
rect 7925 9560 7930 9616
rect 7986 9560 8034 9616
rect 7925 9555 8034 9560
rect 10501 9616 10548 9620
rect 10612 9618 10618 9620
rect 20989 9618 21055 9621
rect 22134 9618 22140 9620
rect 10501 9560 10506 9616
rect 10501 9556 10548 9560
rect 10612 9558 10658 9618
rect 20989 9616 22140 9618
rect 20989 9560 20994 9616
rect 21050 9560 22140 9616
rect 20989 9558 22140 9560
rect 10612 9556 10618 9558
rect 10501 9555 10567 9556
rect 20989 9555 21055 9558
rect 22134 9556 22140 9558
rect 22204 9556 22210 9620
rect 30373 9618 30439 9621
rect 31477 9618 31543 9621
rect 30373 9616 31543 9618
rect 30373 9560 30378 9616
rect 30434 9560 31482 9616
rect 31538 9560 31543 9616
rect 30373 9558 31543 9560
rect 30373 9555 30439 9558
rect 31477 9555 31543 9558
rect 5533 9482 5599 9485
rect 7974 9482 8034 9555
rect 5533 9480 8034 9482
rect 5533 9424 5538 9480
rect 5594 9424 8034 9480
rect 5533 9422 8034 9424
rect 5533 9419 5599 9422
rect 7974 9346 8034 9422
rect 8385 9482 8451 9485
rect 16113 9482 16179 9485
rect 8385 9480 16179 9482
rect 8385 9424 8390 9480
rect 8446 9424 16118 9480
rect 16174 9424 16179 9480
rect 8385 9422 16179 9424
rect 8385 9419 8451 9422
rect 16113 9419 16179 9422
rect 18413 9482 18479 9485
rect 19241 9482 19307 9485
rect 18413 9480 19307 9482
rect 18413 9424 18418 9480
rect 18474 9424 19246 9480
rect 19302 9424 19307 9480
rect 18413 9422 19307 9424
rect 18413 9419 18479 9422
rect 19241 9419 19307 9422
rect 19885 9482 19951 9485
rect 21030 9482 21036 9484
rect 19885 9480 21036 9482
rect 19885 9424 19890 9480
rect 19946 9424 21036 9480
rect 19885 9422 21036 9424
rect 19885 9419 19951 9422
rect 21030 9420 21036 9422
rect 21100 9420 21106 9484
rect 22829 9482 22895 9485
rect 23606 9482 23612 9484
rect 22829 9480 23612 9482
rect 22829 9424 22834 9480
rect 22890 9424 23612 9480
rect 22829 9422 23612 9424
rect 22829 9419 22895 9422
rect 23606 9420 23612 9422
rect 23676 9420 23682 9484
rect 24761 9482 24827 9485
rect 30557 9482 30623 9485
rect 24761 9480 30623 9482
rect 24761 9424 24766 9480
rect 24822 9424 30562 9480
rect 30618 9424 30623 9480
rect 24761 9422 30623 9424
rect 24761 9419 24827 9422
rect 30557 9419 30623 9422
rect 10593 9346 10659 9349
rect 7974 9344 10659 9346
rect 7974 9288 10598 9344
rect 10654 9288 10659 9344
rect 7974 9286 10659 9288
rect 10593 9283 10659 9286
rect 14825 9346 14891 9349
rect 14958 9346 14964 9348
rect 14825 9344 14964 9346
rect 14825 9288 14830 9344
rect 14886 9288 14964 9344
rect 14825 9286 14964 9288
rect 14825 9283 14891 9286
rect 14958 9284 14964 9286
rect 15028 9284 15034 9348
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 6177 9210 6243 9213
rect 6310 9210 6316 9212
rect 6177 9208 6316 9210
rect 6177 9152 6182 9208
rect 6238 9152 6316 9208
rect 6177 9150 6316 9152
rect 6177 9147 6243 9150
rect 6310 9148 6316 9150
rect 6380 9148 6386 9212
rect 6729 9210 6795 9213
rect 8385 9210 8451 9213
rect 6729 9208 8451 9210
rect 6729 9152 6734 9208
rect 6790 9152 8390 9208
rect 8446 9152 8451 9208
rect 6729 9150 8451 9152
rect 6729 9147 6795 9150
rect 8385 9147 8451 9150
rect 15837 9210 15903 9213
rect 25078 9210 25084 9212
rect 15837 9208 25084 9210
rect 15837 9152 15842 9208
rect 15898 9152 25084 9208
rect 15837 9150 25084 9152
rect 15837 9147 15903 9150
rect 25078 9148 25084 9150
rect 25148 9148 25154 9212
rect 31017 9210 31083 9213
rect 31937 9210 32003 9213
rect 32765 9210 32831 9213
rect 31017 9208 32831 9210
rect 31017 9152 31022 9208
rect 31078 9152 31942 9208
rect 31998 9152 32770 9208
rect 32826 9152 32831 9208
rect 31017 9150 32831 9152
rect 31017 9147 31083 9150
rect 31937 9147 32003 9150
rect 32765 9147 32831 9150
rect 5533 9074 5599 9077
rect 17401 9074 17467 9077
rect 5533 9072 17467 9074
rect 5533 9016 5538 9072
rect 5594 9016 17406 9072
rect 17462 9016 17467 9072
rect 5533 9014 17467 9016
rect 5533 9011 5599 9014
rect 17401 9011 17467 9014
rect 24669 9074 24735 9077
rect 33225 9074 33291 9077
rect 24669 9072 33291 9074
rect 24669 9016 24674 9072
rect 24730 9016 33230 9072
rect 33286 9016 33291 9072
rect 24669 9014 33291 9016
rect 24669 9011 24735 9014
rect 33225 9011 33291 9014
rect 5390 8876 5396 8940
rect 5460 8938 5466 8940
rect 10225 8938 10291 8941
rect 5460 8936 10291 8938
rect 5460 8880 10230 8936
rect 10286 8880 10291 8936
rect 5460 8878 10291 8880
rect 5460 8876 5466 8878
rect 10225 8875 10291 8878
rect 10961 8938 11027 8941
rect 16941 8938 17007 8941
rect 10961 8936 17007 8938
rect 10961 8880 10966 8936
rect 11022 8880 16946 8936
rect 17002 8880 17007 8936
rect 10961 8878 17007 8880
rect 10961 8875 11027 8878
rect 16941 8875 17007 8878
rect 17125 8938 17191 8941
rect 17718 8938 17724 8940
rect 17125 8936 17724 8938
rect 17125 8880 17130 8936
rect 17186 8880 17724 8936
rect 17125 8878 17724 8880
rect 17125 8875 17191 8878
rect 17718 8876 17724 8878
rect 17788 8876 17794 8940
rect 18505 8938 18571 8941
rect 30782 8938 30788 8940
rect 18505 8936 30788 8938
rect 18505 8880 18510 8936
rect 18566 8880 30788 8936
rect 18505 8878 30788 8880
rect 18505 8875 18571 8878
rect 30782 8876 30788 8878
rect 30852 8876 30858 8940
rect 31845 8938 31911 8941
rect 32070 8938 32076 8940
rect 31845 8936 32076 8938
rect 31845 8880 31850 8936
rect 31906 8880 32076 8936
rect 31845 8878 32076 8880
rect 31845 8875 31911 8878
rect 32070 8876 32076 8878
rect 32140 8938 32146 8940
rect 36813 8938 36879 8941
rect 32140 8936 36879 8938
rect 32140 8880 36818 8936
rect 36874 8880 36879 8936
rect 32140 8878 36879 8880
rect 32140 8876 32146 8878
rect 36813 8875 36879 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 3049 8802 3115 8805
rect 3918 8802 3924 8804
rect 3049 8800 3924 8802
rect 3049 8744 3054 8800
rect 3110 8744 3924 8800
rect 3049 8742 3924 8744
rect 3049 8739 3115 8742
rect 3918 8740 3924 8742
rect 3988 8740 3994 8804
rect 4705 8802 4771 8805
rect 10869 8802 10935 8805
rect 4705 8800 10935 8802
rect 4705 8744 4710 8800
rect 4766 8744 10874 8800
rect 10930 8744 10935 8800
rect 4705 8742 10935 8744
rect 4705 8739 4771 8742
rect 10869 8739 10935 8742
rect 11513 8802 11579 8805
rect 13169 8802 13235 8805
rect 11513 8800 13235 8802
rect 11513 8744 11518 8800
rect 11574 8744 13174 8800
rect 13230 8744 13235 8800
rect 11513 8742 13235 8744
rect 11513 8739 11579 8742
rect 13169 8739 13235 8742
rect 14549 8802 14615 8805
rect 15745 8802 15811 8805
rect 14549 8800 15811 8802
rect 14549 8744 14554 8800
rect 14610 8744 15750 8800
rect 15806 8744 15811 8800
rect 14549 8742 15811 8744
rect 14549 8739 14615 8742
rect 15745 8739 15811 8742
rect 26877 8802 26943 8805
rect 27705 8802 27771 8805
rect 26877 8800 27771 8802
rect 26877 8744 26882 8800
rect 26938 8744 27710 8800
rect 27766 8744 27771 8800
rect 26877 8742 27771 8744
rect 26877 8739 26943 8742
rect 27705 8739 27771 8742
rect 32673 8802 32739 8805
rect 33225 8802 33291 8805
rect 32673 8800 33291 8802
rect 32673 8744 32678 8800
rect 32734 8744 33230 8800
rect 33286 8744 33291 8800
rect 32673 8742 33291 8744
rect 32673 8739 32739 8742
rect 33225 8739 33291 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4245 8666 4311 8669
rect 9857 8666 9923 8669
rect 4245 8664 9923 8666
rect 4245 8608 4250 8664
rect 4306 8608 9862 8664
rect 9918 8608 9923 8664
rect 4245 8606 9923 8608
rect 4245 8603 4311 8606
rect 9857 8603 9923 8606
rect 12433 8666 12499 8669
rect 15929 8666 15995 8669
rect 12433 8664 15995 8666
rect 12433 8608 12438 8664
rect 12494 8608 15934 8664
rect 15990 8608 15995 8664
rect 12433 8606 15995 8608
rect 12433 8603 12499 8606
rect 15929 8603 15995 8606
rect 23105 8666 23171 8669
rect 32029 8666 32095 8669
rect 23105 8664 32095 8666
rect 23105 8608 23110 8664
rect 23166 8608 32034 8664
rect 32090 8608 32095 8664
rect 23105 8606 32095 8608
rect 23105 8603 23171 8606
rect 32029 8603 32095 8606
rect 32765 8666 32831 8669
rect 33685 8666 33751 8669
rect 32765 8664 33751 8666
rect 32765 8608 32770 8664
rect 32826 8608 33690 8664
rect 33746 8608 33751 8664
rect 32765 8606 33751 8608
rect 32765 8603 32831 8606
rect 33685 8603 33751 8606
rect 6361 8532 6427 8533
rect 6310 8530 6316 8532
rect 6270 8470 6316 8530
rect 6380 8528 6427 8532
rect 6422 8472 6427 8528
rect 6310 8468 6316 8470
rect 6380 8468 6427 8472
rect 6361 8467 6427 8468
rect 7373 8530 7439 8533
rect 11145 8530 11211 8533
rect 16614 8530 16620 8532
rect 7373 8528 9138 8530
rect 7373 8472 7378 8528
rect 7434 8472 9138 8528
rect 7373 8470 9138 8472
rect 7373 8467 7439 8470
rect 6085 8394 6151 8397
rect 7925 8394 7991 8397
rect 6085 8392 7991 8394
rect 6085 8336 6090 8392
rect 6146 8336 7930 8392
rect 7986 8336 7991 8392
rect 6085 8334 7991 8336
rect 9078 8394 9138 8470
rect 11145 8528 16620 8530
rect 11145 8472 11150 8528
rect 11206 8472 16620 8528
rect 11145 8470 16620 8472
rect 11145 8467 11211 8470
rect 16614 8468 16620 8470
rect 16684 8468 16690 8532
rect 24117 8530 24183 8533
rect 27337 8530 27403 8533
rect 28257 8530 28323 8533
rect 24117 8528 28323 8530
rect 24117 8472 24122 8528
rect 24178 8472 27342 8528
rect 27398 8472 28262 8528
rect 28318 8472 28323 8528
rect 24117 8470 28323 8472
rect 24117 8467 24183 8470
rect 27337 8467 27403 8470
rect 28257 8467 28323 8470
rect 30414 8468 30420 8532
rect 30484 8530 30490 8532
rect 30557 8530 30623 8533
rect 30782 8530 30788 8532
rect 30484 8528 30788 8530
rect 30484 8472 30562 8528
rect 30618 8472 30788 8528
rect 30484 8470 30788 8472
rect 30484 8468 30490 8470
rect 30557 8467 30623 8470
rect 30782 8468 30788 8470
rect 30852 8468 30858 8532
rect 9305 8394 9371 8397
rect 9078 8392 9371 8394
rect 9078 8336 9310 8392
rect 9366 8336 9371 8392
rect 9078 8334 9371 8336
rect 6085 8331 6151 8334
rect 7925 8331 7991 8334
rect 9305 8331 9371 8334
rect 15285 8394 15351 8397
rect 16798 8394 16804 8396
rect 15285 8392 16804 8394
rect 15285 8336 15290 8392
rect 15346 8336 16804 8392
rect 15285 8334 16804 8336
rect 15285 8331 15351 8334
rect 16798 8332 16804 8334
rect 16868 8332 16874 8396
rect 17902 8332 17908 8396
rect 17972 8394 17978 8396
rect 19149 8394 19215 8397
rect 17972 8392 19215 8394
rect 17972 8336 19154 8392
rect 19210 8336 19215 8392
rect 17972 8334 19215 8336
rect 17972 8332 17978 8334
rect 19149 8331 19215 8334
rect 22737 8394 22803 8397
rect 24894 8394 24900 8396
rect 22737 8392 24900 8394
rect 22737 8336 22742 8392
rect 22798 8336 24900 8392
rect 22737 8334 24900 8336
rect 22737 8331 22803 8334
rect 24894 8332 24900 8334
rect 24964 8332 24970 8396
rect 29821 8394 29887 8397
rect 34421 8394 34487 8397
rect 29821 8392 34487 8394
rect 29821 8336 29826 8392
rect 29882 8336 34426 8392
rect 34482 8336 34487 8392
rect 29821 8334 34487 8336
rect 29821 8331 29887 8334
rect 34421 8331 34487 8334
rect 200 8258 800 8288
rect 1393 8258 1459 8261
rect 200 8256 1459 8258
rect 200 8200 1398 8256
rect 1454 8200 1459 8256
rect 200 8198 1459 8200
rect 200 8168 800 8198
rect 1393 8195 1459 8198
rect 4981 8258 5047 8261
rect 7741 8258 7807 8261
rect 4981 8256 7807 8258
rect 4981 8200 4986 8256
rect 5042 8200 7746 8256
rect 7802 8200 7807 8256
rect 4981 8198 7807 8200
rect 4981 8195 5047 8198
rect 7741 8195 7807 8198
rect 9949 8258 10015 8261
rect 18229 8258 18295 8261
rect 9949 8256 18295 8258
rect 9949 8200 9954 8256
rect 10010 8200 18234 8256
rect 18290 8200 18295 8256
rect 9949 8198 18295 8200
rect 9949 8195 10015 8198
rect 18229 8195 18295 8198
rect 22277 8260 22343 8261
rect 22277 8256 22324 8260
rect 22388 8258 22394 8260
rect 31201 8258 31267 8261
rect 31661 8258 31727 8261
rect 22277 8200 22282 8256
rect 22277 8196 22324 8200
rect 22388 8198 22434 8258
rect 31201 8256 31727 8258
rect 31201 8200 31206 8256
rect 31262 8200 31666 8256
rect 31722 8200 31727 8256
rect 31201 8198 31727 8200
rect 22388 8196 22394 8198
rect 22277 8195 22343 8196
rect 31201 8195 31267 8198
rect 31661 8195 31727 8198
rect 38193 8258 38259 8261
rect 39200 8258 39800 8288
rect 38193 8256 39800 8258
rect 38193 8200 38198 8256
rect 38254 8200 39800 8256
rect 38193 8198 39800 8200
rect 38193 8195 38259 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 5349 8122 5415 8125
rect 7833 8122 7899 8125
rect 5349 8120 7899 8122
rect 5349 8064 5354 8120
rect 5410 8064 7838 8120
rect 7894 8064 7899 8120
rect 5349 8062 7899 8064
rect 5349 8059 5415 8062
rect 7833 8059 7899 8062
rect 16297 8122 16363 8125
rect 16430 8122 16436 8124
rect 16297 8120 16436 8122
rect 16297 8064 16302 8120
rect 16358 8064 16436 8120
rect 16297 8062 16436 8064
rect 16297 8059 16363 8062
rect 16430 8060 16436 8062
rect 16500 8060 16506 8124
rect 17861 8122 17927 8125
rect 21173 8122 21239 8125
rect 17861 8120 21239 8122
rect 17861 8064 17866 8120
rect 17922 8064 21178 8120
rect 21234 8064 21239 8120
rect 17861 8062 21239 8064
rect 17861 8059 17927 8062
rect 21173 8059 21239 8062
rect 27061 8122 27127 8125
rect 27521 8122 27587 8125
rect 27061 8120 27587 8122
rect 27061 8064 27066 8120
rect 27122 8064 27526 8120
rect 27582 8064 27587 8120
rect 27061 8062 27587 8064
rect 27061 8059 27127 8062
rect 27521 8059 27587 8062
rect 30465 8122 30531 8125
rect 32857 8122 32923 8125
rect 30465 8120 32923 8122
rect 30465 8064 30470 8120
rect 30526 8064 32862 8120
rect 32918 8064 32923 8120
rect 30465 8062 32923 8064
rect 30465 8059 30531 8062
rect 32857 8059 32923 8062
rect 3325 7986 3391 7989
rect 30414 7986 30420 7988
rect 3325 7984 30420 7986
rect 3325 7928 3330 7984
rect 3386 7928 30420 7984
rect 3325 7926 30420 7928
rect 3325 7923 3391 7926
rect 30414 7924 30420 7926
rect 30484 7924 30490 7988
rect 5349 7850 5415 7853
rect 7833 7850 7899 7853
rect 5349 7848 7899 7850
rect 5349 7792 5354 7848
rect 5410 7792 7838 7848
rect 7894 7792 7899 7848
rect 5349 7790 7899 7792
rect 5349 7787 5415 7790
rect 7833 7787 7899 7790
rect 21173 7850 21239 7853
rect 22502 7850 22508 7852
rect 21173 7848 22508 7850
rect 21173 7792 21178 7848
rect 21234 7792 22508 7848
rect 21173 7790 22508 7792
rect 21173 7787 21239 7790
rect 22502 7788 22508 7790
rect 22572 7788 22578 7852
rect 26141 7850 26207 7853
rect 33593 7850 33659 7853
rect 26141 7848 33659 7850
rect 26141 7792 26146 7848
rect 26202 7792 33598 7848
rect 33654 7792 33659 7848
rect 26141 7790 33659 7792
rect 26141 7787 26207 7790
rect 33593 7787 33659 7790
rect 5022 7714 5028 7716
rect 2270 7654 5028 7714
rect 200 7578 800 7608
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 2270 7173 2330 7654
rect 5022 7652 5028 7654
rect 5092 7652 5098 7716
rect 7005 7714 7071 7717
rect 8569 7714 8635 7717
rect 7005 7712 8635 7714
rect 7005 7656 7010 7712
rect 7066 7656 8574 7712
rect 8630 7656 8635 7712
rect 7005 7654 8635 7656
rect 7005 7651 7071 7654
rect 8569 7651 8635 7654
rect 22185 7714 22251 7717
rect 26693 7714 26759 7717
rect 27429 7716 27495 7717
rect 27429 7714 27476 7716
rect 22185 7712 26759 7714
rect 22185 7656 22190 7712
rect 22246 7656 26698 7712
rect 26754 7656 26759 7712
rect 22185 7654 26759 7656
rect 27384 7712 27476 7714
rect 27384 7656 27434 7712
rect 27384 7654 27476 7656
rect 22185 7651 22251 7654
rect 26693 7651 26759 7654
rect 27429 7652 27476 7654
rect 27540 7652 27546 7716
rect 28901 7714 28967 7717
rect 31017 7714 31083 7717
rect 28901 7712 31083 7714
rect 28901 7656 28906 7712
rect 28962 7656 31022 7712
rect 31078 7656 31083 7712
rect 28901 7654 31083 7656
rect 27429 7651 27495 7652
rect 28901 7651 28967 7654
rect 31017 7651 31083 7654
rect 31569 7712 31635 7717
rect 31569 7656 31574 7712
rect 31630 7656 31635 7712
rect 31569 7651 31635 7656
rect 32070 7652 32076 7716
rect 32140 7714 32146 7716
rect 33133 7714 33199 7717
rect 32140 7712 33199 7714
rect 32140 7656 33138 7712
rect 33194 7656 33199 7712
rect 32140 7654 33199 7656
rect 32140 7652 32146 7654
rect 33133 7651 33199 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4613 7578 4679 7581
rect 8845 7578 8911 7581
rect 4613 7576 8911 7578
rect 4613 7520 4618 7576
rect 4674 7520 8850 7576
rect 8906 7520 8911 7576
rect 4613 7518 8911 7520
rect 4613 7515 4679 7518
rect 8845 7515 8911 7518
rect 17401 7578 17467 7581
rect 18505 7578 18571 7581
rect 17401 7576 18571 7578
rect 17401 7520 17406 7576
rect 17462 7520 18510 7576
rect 18566 7520 18571 7576
rect 17401 7518 18571 7520
rect 17401 7515 17467 7518
rect 18505 7515 18571 7518
rect 26693 7578 26759 7581
rect 27337 7578 27403 7581
rect 26693 7576 27403 7578
rect 26693 7520 26698 7576
rect 26754 7520 27342 7576
rect 27398 7520 27403 7576
rect 26693 7518 27403 7520
rect 31572 7578 31632 7651
rect 34053 7578 34119 7581
rect 31572 7576 34119 7578
rect 31572 7520 34058 7576
rect 34114 7520 34119 7576
rect 31572 7518 34119 7520
rect 26693 7515 26759 7518
rect 27337 7515 27403 7518
rect 34053 7515 34119 7518
rect 38193 7578 38259 7581
rect 39200 7578 39800 7608
rect 38193 7576 39800 7578
rect 38193 7520 38198 7576
rect 38254 7520 39800 7576
rect 38193 7518 39800 7520
rect 38193 7515 38259 7518
rect 39200 7488 39800 7518
rect 3509 7442 3575 7445
rect 8017 7442 8083 7445
rect 3509 7440 8083 7442
rect 3509 7384 3514 7440
rect 3570 7384 8022 7440
rect 8078 7384 8083 7440
rect 3509 7382 8083 7384
rect 3509 7379 3575 7382
rect 8017 7379 8083 7382
rect 16941 7442 17007 7445
rect 20161 7442 20227 7445
rect 16941 7440 20227 7442
rect 16941 7384 16946 7440
rect 17002 7384 20166 7440
rect 20222 7384 20227 7440
rect 16941 7382 20227 7384
rect 16941 7379 17007 7382
rect 20161 7379 20227 7382
rect 23381 7442 23447 7445
rect 35709 7442 35775 7445
rect 23381 7440 35775 7442
rect 23381 7384 23386 7440
rect 23442 7384 35714 7440
rect 35770 7384 35775 7440
rect 23381 7382 35775 7384
rect 23381 7379 23447 7382
rect 35709 7379 35775 7382
rect 4521 7306 4587 7309
rect 14590 7306 14596 7308
rect 4521 7304 14596 7306
rect 4521 7248 4526 7304
rect 4582 7248 14596 7304
rect 4521 7246 14596 7248
rect 4521 7243 4587 7246
rect 14590 7244 14596 7246
rect 14660 7244 14666 7308
rect 14733 7306 14799 7309
rect 16021 7306 16087 7309
rect 14733 7304 16087 7306
rect 14733 7248 14738 7304
rect 14794 7248 16026 7304
rect 16082 7248 16087 7304
rect 14733 7246 16087 7248
rect 14733 7243 14799 7246
rect 16021 7243 16087 7246
rect 21081 7306 21147 7309
rect 32949 7306 33015 7309
rect 21081 7304 33015 7306
rect 21081 7248 21086 7304
rect 21142 7248 32954 7304
rect 33010 7248 33015 7304
rect 21081 7246 33015 7248
rect 21081 7243 21147 7246
rect 32949 7243 33015 7246
rect 2221 7168 2330 7173
rect 2221 7112 2226 7168
rect 2282 7112 2330 7168
rect 2221 7110 2330 7112
rect 6269 7170 6335 7173
rect 9673 7170 9739 7173
rect 6269 7168 9739 7170
rect 6269 7112 6274 7168
rect 6330 7112 9678 7168
rect 9734 7112 9739 7168
rect 6269 7110 9739 7112
rect 2221 7107 2287 7110
rect 6269 7107 6335 7110
rect 9673 7107 9739 7110
rect 11605 7170 11671 7173
rect 13813 7170 13879 7173
rect 18965 7170 19031 7173
rect 11605 7168 13600 7170
rect 11605 7112 11610 7168
rect 11666 7112 13600 7168
rect 11605 7110 13600 7112
rect 11605 7107 11671 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 13540 7037 13600 7110
rect 13813 7168 19031 7170
rect 13813 7112 13818 7168
rect 13874 7112 18970 7168
rect 19026 7112 19031 7168
rect 13813 7110 19031 7112
rect 13813 7107 13879 7110
rect 18965 7107 19031 7110
rect 26601 7170 26667 7173
rect 27521 7170 27587 7173
rect 26601 7168 27587 7170
rect 26601 7112 26606 7168
rect 26662 7112 27526 7168
rect 27582 7112 27587 7168
rect 26601 7110 27587 7112
rect 26601 7107 26667 7110
rect 27521 7107 27587 7110
rect 31477 7170 31543 7173
rect 34237 7170 34303 7173
rect 31477 7168 34303 7170
rect 31477 7112 31482 7168
rect 31538 7112 34242 7168
rect 34298 7112 34303 7168
rect 31477 7110 34303 7112
rect 31477 7107 31543 7110
rect 34237 7107 34303 7110
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 5073 7034 5139 7037
rect 7833 7034 7899 7037
rect 5073 7032 7899 7034
rect 5073 6976 5078 7032
rect 5134 6976 7838 7032
rect 7894 6976 7899 7032
rect 5073 6974 7899 6976
rect 5073 6971 5139 6974
rect 7833 6971 7899 6974
rect 11881 7034 11947 7037
rect 12433 7034 12499 7037
rect 11881 7032 12499 7034
rect 11881 6976 11886 7032
rect 11942 6976 12438 7032
rect 12494 6976 12499 7032
rect 11881 6974 12499 6976
rect 11881 6971 11947 6974
rect 12433 6971 12499 6974
rect 13537 7034 13603 7037
rect 17585 7034 17651 7037
rect 13537 7032 17651 7034
rect 13537 6976 13542 7032
rect 13598 6976 17590 7032
rect 17646 6976 17651 7032
rect 13537 6974 17651 6976
rect 13537 6971 13603 6974
rect 17585 6971 17651 6974
rect 18873 7034 18939 7037
rect 20529 7034 20595 7037
rect 18873 7032 20595 7034
rect 18873 6976 18878 7032
rect 18934 6976 20534 7032
rect 20590 6976 20595 7032
rect 18873 6974 20595 6976
rect 18873 6971 18939 6974
rect 20529 6971 20595 6974
rect 24761 7034 24827 7037
rect 26325 7034 26391 7037
rect 31569 7036 31635 7037
rect 31518 7034 31524 7036
rect 24761 7032 26250 7034
rect 24761 6976 24766 7032
rect 24822 6976 26250 7032
rect 24761 6974 26250 6976
rect 24761 6971 24827 6974
rect 5073 6898 5139 6901
rect 7833 6900 7899 6901
rect 5206 6898 5212 6900
rect 5073 6896 5212 6898
rect 5073 6840 5078 6896
rect 5134 6840 5212 6896
rect 5073 6838 5212 6840
rect 5073 6835 5139 6838
rect 5206 6836 5212 6838
rect 5276 6836 5282 6900
rect 7782 6898 7788 6900
rect 7742 6838 7788 6898
rect 7852 6896 7899 6900
rect 7894 6840 7899 6896
rect 7782 6836 7788 6838
rect 7852 6836 7899 6840
rect 7833 6835 7899 6836
rect 8201 6898 8267 6901
rect 8753 6900 8819 6901
rect 8334 6898 8340 6900
rect 8201 6896 8340 6898
rect 8201 6840 8206 6896
rect 8262 6840 8340 6896
rect 8201 6838 8340 6840
rect 8201 6835 8267 6838
rect 8334 6836 8340 6838
rect 8404 6836 8410 6900
rect 8702 6898 8708 6900
rect 8662 6838 8708 6898
rect 8772 6896 8819 6900
rect 8814 6840 8819 6896
rect 8702 6836 8708 6838
rect 8772 6836 8819 6840
rect 8753 6835 8819 6836
rect 9305 6898 9371 6901
rect 12617 6900 12683 6901
rect 9305 6896 12450 6898
rect 9305 6840 9310 6896
rect 9366 6840 12450 6896
rect 9305 6838 12450 6840
rect 9305 6835 9371 6838
rect 2589 6762 2655 6765
rect 6862 6762 6868 6764
rect 2589 6760 6868 6762
rect 2589 6704 2594 6760
rect 2650 6704 6868 6760
rect 2589 6702 6868 6704
rect 2589 6699 2655 6702
rect 6862 6700 6868 6702
rect 6932 6700 6938 6764
rect 8518 6700 8524 6764
rect 8588 6762 8594 6764
rect 10593 6762 10659 6765
rect 8588 6760 10659 6762
rect 8588 6704 10598 6760
rect 10654 6704 10659 6760
rect 8588 6702 10659 6704
rect 12390 6762 12450 6838
rect 12566 6836 12572 6900
rect 12636 6898 12683 6900
rect 13077 6900 13143 6901
rect 13077 6898 13124 6900
rect 12636 6896 12728 6898
rect 12678 6840 12728 6896
rect 12636 6838 12728 6840
rect 13032 6896 13124 6898
rect 13032 6840 13082 6896
rect 13032 6838 13124 6840
rect 12636 6836 12683 6838
rect 12617 6835 12683 6836
rect 13077 6836 13124 6838
rect 13188 6836 13194 6900
rect 17401 6898 17467 6901
rect 20437 6898 20503 6901
rect 17401 6896 20503 6898
rect 17401 6840 17406 6896
rect 17462 6840 20442 6896
rect 20498 6840 20503 6896
rect 17401 6838 20503 6840
rect 13077 6835 13143 6836
rect 17401 6835 17467 6838
rect 20437 6835 20503 6838
rect 21950 6836 21956 6900
rect 22020 6898 22026 6900
rect 22737 6898 22803 6901
rect 22020 6896 22803 6898
rect 22020 6840 22742 6896
rect 22798 6840 22803 6896
rect 22020 6838 22803 6840
rect 22020 6836 22026 6838
rect 22737 6835 22803 6838
rect 25589 6900 25655 6901
rect 25589 6896 25636 6900
rect 25700 6898 25706 6900
rect 26190 6898 26250 6974
rect 26325 7032 31524 7034
rect 31588 7032 31635 7036
rect 26325 6976 26330 7032
rect 26386 6976 31524 7032
rect 31630 6976 31635 7032
rect 26325 6974 31524 6976
rect 26325 6971 26391 6974
rect 31518 6972 31524 6974
rect 31588 6972 31635 6976
rect 31569 6971 31635 6972
rect 31937 7034 32003 7037
rect 32949 7034 33015 7037
rect 31937 7032 33015 7034
rect 31937 6976 31942 7032
rect 31998 6976 32954 7032
rect 33010 6976 33015 7032
rect 31937 6974 33015 6976
rect 31937 6971 32003 6974
rect 32949 6971 33015 6974
rect 26785 6898 26851 6901
rect 28625 6898 28691 6901
rect 25589 6840 25594 6896
rect 25589 6836 25636 6840
rect 25700 6838 25746 6898
rect 26190 6896 28691 6898
rect 26190 6840 26790 6896
rect 26846 6840 28630 6896
rect 28686 6840 28691 6896
rect 26190 6838 28691 6840
rect 25700 6836 25706 6838
rect 25589 6835 25655 6836
rect 26785 6835 26851 6838
rect 28625 6835 28691 6838
rect 30414 6836 30420 6900
rect 30484 6898 30490 6900
rect 33501 6898 33567 6901
rect 30484 6896 33567 6898
rect 30484 6840 33506 6896
rect 33562 6840 33567 6896
rect 30484 6838 33567 6840
rect 30484 6836 30490 6838
rect 33501 6835 33567 6838
rect 30373 6762 30439 6765
rect 12390 6760 30439 6762
rect 12390 6704 30378 6760
rect 30434 6704 30439 6760
rect 12390 6702 30439 6704
rect 8588 6700 8594 6702
rect 10593 6699 10659 6702
rect 30373 6699 30439 6702
rect 36261 6762 36327 6765
rect 36445 6762 36511 6765
rect 36261 6760 36511 6762
rect 36261 6704 36266 6760
rect 36322 6704 36450 6760
rect 36506 6704 36511 6760
rect 36261 6702 36511 6704
rect 36261 6699 36327 6702
rect 36445 6699 36511 6702
rect 3877 6626 3943 6629
rect 9622 6626 9628 6628
rect 3877 6624 9628 6626
rect 3877 6568 3882 6624
rect 3938 6568 9628 6624
rect 3877 6566 9628 6568
rect 3877 6563 3943 6566
rect 9622 6564 9628 6566
rect 9692 6564 9698 6628
rect 24301 6626 24367 6629
rect 30557 6626 30623 6629
rect 24301 6624 30623 6626
rect 24301 6568 24306 6624
rect 24362 6568 30562 6624
rect 30618 6568 30623 6624
rect 24301 6566 30623 6568
rect 24301 6563 24367 6566
rect 30557 6563 30623 6566
rect 30782 6564 30788 6628
rect 30852 6626 30858 6628
rect 32305 6626 32371 6629
rect 30852 6624 32371 6626
rect 30852 6568 32310 6624
rect 32366 6568 32371 6624
rect 30852 6566 32371 6568
rect 30852 6564 30858 6566
rect 32305 6563 32371 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 7741 6490 7807 6493
rect 9489 6490 9555 6493
rect 7741 6488 9555 6490
rect 7741 6432 7746 6488
rect 7802 6432 9494 6488
rect 9550 6432 9555 6488
rect 7741 6430 9555 6432
rect 7741 6427 7807 6430
rect 9489 6427 9555 6430
rect 11329 6490 11395 6493
rect 19149 6490 19215 6493
rect 11329 6488 19215 6490
rect 11329 6432 11334 6488
rect 11390 6432 19154 6488
rect 19210 6432 19215 6488
rect 11329 6430 19215 6432
rect 11329 6427 11395 6430
rect 19149 6427 19215 6430
rect 20253 6490 20319 6493
rect 23197 6490 23263 6493
rect 20253 6488 23263 6490
rect 20253 6432 20258 6488
rect 20314 6432 23202 6488
rect 23258 6432 23263 6488
rect 20253 6430 23263 6432
rect 20253 6427 20319 6430
rect 23197 6427 23263 6430
rect 27429 6492 27495 6493
rect 27429 6488 27476 6492
rect 27540 6490 27546 6492
rect 28073 6490 28139 6493
rect 35709 6490 35775 6493
rect 27429 6432 27434 6488
rect 27429 6428 27476 6432
rect 27540 6430 27586 6490
rect 28073 6488 35775 6490
rect 28073 6432 28078 6488
rect 28134 6432 35714 6488
rect 35770 6432 35775 6488
rect 28073 6430 35775 6432
rect 27540 6428 27546 6430
rect 27429 6427 27495 6428
rect 28073 6427 28139 6430
rect 35709 6427 35775 6430
rect 4245 6354 4311 6357
rect 5758 6354 5764 6356
rect 4245 6352 5764 6354
rect 4245 6296 4250 6352
rect 4306 6296 5764 6352
rect 4245 6294 5764 6296
rect 4245 6291 4311 6294
rect 5758 6292 5764 6294
rect 5828 6354 5834 6356
rect 10685 6354 10751 6357
rect 5828 6352 10751 6354
rect 5828 6296 10690 6352
rect 10746 6296 10751 6352
rect 5828 6294 10751 6296
rect 5828 6292 5834 6294
rect 10685 6291 10751 6294
rect 21449 6354 21515 6357
rect 30189 6354 30255 6357
rect 32397 6354 32463 6357
rect 21449 6352 22110 6354
rect 21449 6296 21454 6352
rect 21510 6296 22110 6352
rect 21449 6294 22110 6296
rect 21449 6291 21515 6294
rect 200 6218 800 6248
rect 1761 6218 1827 6221
rect 200 6216 1827 6218
rect 200 6160 1766 6216
rect 1822 6160 1827 6216
rect 200 6158 1827 6160
rect 200 6128 800 6158
rect 1761 6155 1827 6158
rect 6821 6218 6887 6221
rect 18229 6218 18295 6221
rect 6821 6216 18295 6218
rect 6821 6160 6826 6216
rect 6882 6160 18234 6216
rect 18290 6160 18295 6216
rect 6821 6158 18295 6160
rect 22050 6218 22110 6294
rect 30189 6352 32463 6354
rect 30189 6296 30194 6352
rect 30250 6296 32402 6352
rect 32458 6296 32463 6352
rect 30189 6294 32463 6296
rect 30189 6291 30255 6294
rect 32397 6291 32463 6294
rect 33685 6354 33751 6357
rect 34789 6354 34855 6357
rect 33685 6352 34855 6354
rect 33685 6296 33690 6352
rect 33746 6296 34794 6352
rect 34850 6296 34855 6352
rect 33685 6294 34855 6296
rect 33685 6291 33751 6294
rect 34789 6291 34855 6294
rect 35801 6354 35867 6357
rect 35801 6352 38394 6354
rect 35801 6296 35806 6352
rect 35862 6296 38394 6352
rect 35801 6294 38394 6296
rect 35801 6291 35867 6294
rect 38193 6218 38259 6221
rect 22050 6216 38259 6218
rect 22050 6160 38198 6216
rect 38254 6160 38259 6216
rect 22050 6158 38259 6160
rect 38334 6218 38394 6294
rect 39200 6218 39800 6248
rect 38334 6158 39800 6218
rect 6821 6155 6887 6158
rect 18229 6155 18295 6158
rect 38193 6155 38259 6158
rect 39200 6128 39800 6158
rect 7373 6082 7439 6085
rect 8753 6082 8819 6085
rect 7373 6080 8819 6082
rect 7373 6024 7378 6080
rect 7434 6024 8758 6080
rect 8814 6024 8819 6080
rect 7373 6022 8819 6024
rect 7373 6019 7439 6022
rect 8753 6019 8819 6022
rect 21817 6082 21883 6085
rect 22277 6082 22343 6085
rect 21817 6080 22343 6082
rect 21817 6024 21822 6080
rect 21878 6024 22282 6080
rect 22338 6024 22343 6080
rect 21817 6022 22343 6024
rect 21817 6019 21883 6022
rect 22277 6019 22343 6022
rect 29545 6082 29611 6085
rect 29545 6080 33978 6082
rect 29545 6024 29550 6080
rect 29606 6024 33978 6080
rect 29545 6022 33978 6024
rect 29545 6019 29611 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 1853 5948 1919 5949
rect 1853 5946 1900 5948
rect 1808 5944 1900 5946
rect 1808 5888 1858 5944
rect 1808 5886 1900 5888
rect 1853 5884 1900 5886
rect 1964 5884 1970 5948
rect 22645 5946 22711 5949
rect 27521 5946 27587 5949
rect 22645 5944 27587 5946
rect 22645 5888 22650 5944
rect 22706 5888 27526 5944
rect 27582 5888 27587 5944
rect 22645 5886 27587 5888
rect 1853 5883 1919 5884
rect 22645 5883 22711 5886
rect 27521 5883 27587 5886
rect 30281 5946 30347 5949
rect 30649 5946 30715 5949
rect 30281 5944 30715 5946
rect 30281 5888 30286 5944
rect 30342 5888 30654 5944
rect 30710 5888 30715 5944
rect 30281 5886 30715 5888
rect 30281 5883 30347 5886
rect 30649 5883 30715 5886
rect 4245 5810 4311 5813
rect 8293 5810 8359 5813
rect 4245 5808 8359 5810
rect 4245 5752 4250 5808
rect 4306 5752 8298 5808
rect 8354 5752 8359 5808
rect 4245 5750 8359 5752
rect 4245 5747 4311 5750
rect 8293 5747 8359 5750
rect 9765 5810 9831 5813
rect 12750 5810 12756 5812
rect 9765 5808 12756 5810
rect 9765 5752 9770 5808
rect 9826 5752 12756 5808
rect 9765 5750 12756 5752
rect 9765 5747 9831 5750
rect 12750 5748 12756 5750
rect 12820 5748 12826 5812
rect 16573 5810 16639 5813
rect 17677 5810 17743 5813
rect 16573 5808 17743 5810
rect 16573 5752 16578 5808
rect 16634 5752 17682 5808
rect 17738 5752 17743 5808
rect 16573 5750 17743 5752
rect 16573 5747 16639 5750
rect 17677 5747 17743 5750
rect 24577 5810 24643 5813
rect 28257 5812 28323 5813
rect 28206 5810 28212 5812
rect 24577 5808 28212 5810
rect 28276 5810 28323 5812
rect 30373 5810 30439 5813
rect 32121 5810 32187 5813
rect 28276 5808 28368 5810
rect 24577 5752 24582 5808
rect 24638 5752 28212 5808
rect 28318 5752 28368 5808
rect 24577 5750 28212 5752
rect 24577 5747 24643 5750
rect 28206 5748 28212 5750
rect 28276 5750 28368 5752
rect 30373 5808 32187 5810
rect 30373 5752 30378 5808
rect 30434 5752 32126 5808
rect 32182 5752 32187 5808
rect 30373 5750 32187 5752
rect 33918 5810 33978 6022
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 36169 5810 36235 5813
rect 33918 5808 36235 5810
rect 33918 5752 36174 5808
rect 36230 5752 36235 5808
rect 33918 5750 36235 5752
rect 28276 5748 28323 5750
rect 28257 5747 28323 5748
rect 30373 5747 30439 5750
rect 32121 5747 32187 5750
rect 36169 5747 36235 5750
rect 6361 5674 6427 5677
rect 6494 5674 6500 5676
rect 6361 5672 6500 5674
rect 6361 5616 6366 5672
rect 6422 5616 6500 5672
rect 6361 5614 6500 5616
rect 6361 5611 6427 5614
rect 6494 5612 6500 5614
rect 6564 5612 6570 5676
rect 6862 5612 6868 5676
rect 6932 5674 6938 5676
rect 11421 5674 11487 5677
rect 6932 5672 11487 5674
rect 6932 5616 11426 5672
rect 11482 5616 11487 5672
rect 6932 5614 11487 5616
rect 6932 5612 6938 5614
rect 11421 5611 11487 5614
rect 26785 5674 26851 5677
rect 31569 5674 31635 5677
rect 26785 5672 31635 5674
rect 26785 5616 26790 5672
rect 26846 5616 31574 5672
rect 31630 5616 31635 5672
rect 26785 5614 31635 5616
rect 26785 5611 26851 5614
rect 31569 5611 31635 5614
rect 31753 5674 31819 5677
rect 34329 5674 34395 5677
rect 31753 5672 34395 5674
rect 31753 5616 31758 5672
rect 31814 5616 34334 5672
rect 34390 5616 34395 5672
rect 31753 5614 34395 5616
rect 31753 5611 31819 5614
rect 34329 5611 34395 5614
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 2129 5538 2195 5541
rect 7005 5540 7071 5541
rect 7557 5540 7623 5541
rect 16113 5540 16179 5541
rect 7005 5538 7052 5540
rect 2129 5536 2790 5538
rect 2129 5480 2134 5536
rect 2190 5480 2790 5536
rect 2129 5478 2790 5480
rect 6960 5536 7052 5538
rect 6960 5480 7010 5536
rect 6960 5478 7052 5480
rect 2129 5475 2195 5478
rect 2730 5402 2790 5478
rect 7005 5476 7052 5478
rect 7116 5476 7122 5540
rect 7557 5536 7604 5540
rect 7668 5538 7674 5540
rect 16062 5538 16068 5540
rect 7557 5480 7562 5536
rect 7557 5476 7604 5480
rect 7668 5478 7714 5538
rect 16022 5478 16068 5538
rect 16132 5536 16179 5540
rect 16174 5480 16179 5536
rect 7668 5476 7674 5478
rect 16062 5476 16068 5478
rect 16132 5476 16179 5480
rect 7005 5475 7071 5476
rect 7557 5475 7623 5476
rect 16113 5475 16179 5476
rect 22277 5538 22343 5541
rect 28390 5538 28396 5540
rect 22277 5536 28396 5538
rect 22277 5480 22282 5536
rect 22338 5480 28396 5536
rect 22277 5478 28396 5480
rect 22277 5475 22343 5478
rect 28390 5476 28396 5478
rect 28460 5476 28466 5540
rect 29637 5538 29703 5541
rect 30465 5538 30531 5541
rect 29637 5536 30531 5538
rect 29637 5480 29642 5536
rect 29698 5480 30470 5536
rect 30526 5480 30531 5536
rect 29637 5478 30531 5480
rect 29637 5475 29703 5478
rect 30465 5475 30531 5478
rect 33726 5476 33732 5540
rect 33796 5538 33802 5540
rect 34329 5538 34395 5541
rect 33796 5536 34395 5538
rect 33796 5480 34334 5536
rect 34390 5480 34395 5536
rect 33796 5478 34395 5480
rect 33796 5476 33802 5478
rect 34329 5475 34395 5478
rect 36721 5538 36787 5541
rect 36854 5538 36860 5540
rect 36721 5536 36860 5538
rect 36721 5480 36726 5536
rect 36782 5480 36860 5536
rect 36721 5478 36860 5480
rect 36721 5475 36787 5478
rect 36854 5476 36860 5478
rect 36924 5476 36930 5540
rect 38377 5538 38443 5541
rect 39200 5538 39800 5568
rect 38377 5536 39800 5538
rect 38377 5480 38382 5536
rect 38438 5480 39800 5536
rect 38377 5478 39800 5480
rect 38377 5475 38443 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 13721 5402 13787 5405
rect 15101 5404 15167 5405
rect 15101 5402 15148 5404
rect 2730 5400 13787 5402
rect 2730 5344 13726 5400
rect 13782 5344 13787 5400
rect 2730 5342 13787 5344
rect 15056 5400 15148 5402
rect 15056 5344 15106 5400
rect 15056 5342 15148 5344
rect 13721 5339 13787 5342
rect 15101 5340 15148 5342
rect 15212 5340 15218 5404
rect 15878 5340 15884 5404
rect 15948 5402 15954 5404
rect 16297 5402 16363 5405
rect 15948 5400 16363 5402
rect 15948 5344 16302 5400
rect 16358 5344 16363 5400
rect 15948 5342 16363 5344
rect 15948 5340 15954 5342
rect 15101 5339 15167 5340
rect 16297 5339 16363 5342
rect 30189 5402 30255 5405
rect 31477 5402 31543 5405
rect 30189 5400 31543 5402
rect 30189 5344 30194 5400
rect 30250 5344 31482 5400
rect 31538 5344 31543 5400
rect 30189 5342 31543 5344
rect 30189 5339 30255 5342
rect 31477 5339 31543 5342
rect 31845 5402 31911 5405
rect 33869 5402 33935 5405
rect 31845 5400 33935 5402
rect 31845 5344 31850 5400
rect 31906 5344 33874 5400
rect 33930 5344 33935 5400
rect 31845 5342 33935 5344
rect 31845 5339 31911 5342
rect 33869 5339 33935 5342
rect 7005 5266 7071 5269
rect 9121 5266 9187 5269
rect 7005 5264 9187 5266
rect 7005 5208 7010 5264
rect 7066 5208 9126 5264
rect 9182 5208 9187 5264
rect 7005 5206 9187 5208
rect 7005 5203 7071 5206
rect 9121 5203 9187 5206
rect 31569 5266 31635 5269
rect 32305 5266 32371 5269
rect 31569 5264 32371 5266
rect 31569 5208 31574 5264
rect 31630 5208 32310 5264
rect 32366 5208 32371 5264
rect 31569 5206 32371 5208
rect 31569 5203 31635 5206
rect 32305 5203 32371 5206
rect 5625 5130 5691 5133
rect 8109 5130 8175 5133
rect 5625 5128 8175 5130
rect 5625 5072 5630 5128
rect 5686 5072 8114 5128
rect 8170 5072 8175 5128
rect 5625 5070 8175 5072
rect 5625 5067 5691 5070
rect 8109 5067 8175 5070
rect 9397 5130 9463 5133
rect 28942 5130 28948 5132
rect 9397 5128 28948 5130
rect 9397 5072 9402 5128
rect 9458 5072 28948 5128
rect 9397 5070 28948 5072
rect 9397 5067 9463 5070
rect 28942 5068 28948 5070
rect 29012 5068 29018 5132
rect 32213 5130 32279 5133
rect 34053 5130 34119 5133
rect 34881 5130 34947 5133
rect 32213 5128 34947 5130
rect 32213 5072 32218 5128
rect 32274 5072 34058 5128
rect 34114 5072 34886 5128
rect 34942 5072 34947 5128
rect 32213 5070 34947 5072
rect 32213 5067 32279 5070
rect 34053 5067 34119 5070
rect 34881 5067 34947 5070
rect 5717 4994 5783 4997
rect 7833 4994 7899 4997
rect 5717 4992 7899 4994
rect 5717 4936 5722 4992
rect 5778 4936 7838 4992
rect 7894 4936 7899 4992
rect 5717 4934 7899 4936
rect 5717 4931 5783 4934
rect 7833 4931 7899 4934
rect 13997 4994 14063 4997
rect 15101 4994 15167 4997
rect 17309 4994 17375 4997
rect 13997 4992 17375 4994
rect 13997 4936 14002 4992
rect 14058 4936 15106 4992
rect 15162 4936 17314 4992
rect 17370 4936 17375 4992
rect 13997 4934 17375 4936
rect 13997 4931 14063 4934
rect 15101 4931 15167 4934
rect 17309 4931 17375 4934
rect 17585 4994 17651 4997
rect 22369 4994 22435 4997
rect 17585 4992 22435 4994
rect 17585 4936 17590 4992
rect 17646 4936 22374 4992
rect 22430 4936 22435 4992
rect 17585 4934 22435 4936
rect 17585 4931 17651 4934
rect 22369 4931 22435 4934
rect 24393 4994 24459 4997
rect 32857 4994 32923 4997
rect 24393 4992 32923 4994
rect 24393 4936 24398 4992
rect 24454 4936 32862 4992
rect 32918 4936 32923 4992
rect 24393 4934 32923 4936
rect 24393 4931 24459 4934
rect 32857 4931 32923 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 2865 4858 2931 4861
rect 200 4856 2931 4858
rect 200 4800 2870 4856
rect 2926 4800 2931 4856
rect 200 4798 2931 4800
rect 200 4768 800 4798
rect 2865 4795 2931 4798
rect 13721 4858 13787 4861
rect 24396 4858 24456 4931
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 13721 4856 24456 4858
rect 13721 4800 13726 4856
rect 13782 4800 24456 4856
rect 13721 4798 24456 4800
rect 30373 4858 30439 4861
rect 34237 4858 34303 4861
rect 30373 4856 34303 4858
rect 30373 4800 30378 4856
rect 30434 4800 34242 4856
rect 34298 4800 34303 4856
rect 30373 4798 34303 4800
rect 13721 4795 13787 4798
rect 30373 4795 30439 4798
rect 34237 4795 34303 4798
rect 3049 4722 3115 4725
rect 26785 4722 26851 4725
rect 3049 4720 26851 4722
rect 3049 4664 3054 4720
rect 3110 4664 26790 4720
rect 26846 4664 26851 4720
rect 3049 4662 26851 4664
rect 3049 4659 3115 4662
rect 26785 4659 26851 4662
rect 30097 4722 30163 4725
rect 36629 4722 36695 4725
rect 30097 4720 36695 4722
rect 30097 4664 30102 4720
rect 30158 4664 36634 4720
rect 36690 4664 36695 4720
rect 30097 4662 36695 4664
rect 30097 4659 30163 4662
rect 36629 4659 36695 4662
rect 13905 4586 13971 4589
rect 17401 4586 17467 4589
rect 18873 4586 18939 4589
rect 13905 4584 18939 4586
rect 13905 4528 13910 4584
rect 13966 4528 17406 4584
rect 17462 4528 18878 4584
rect 18934 4528 18939 4584
rect 13905 4526 18939 4528
rect 13905 4523 13971 4526
rect 17401 4523 17467 4526
rect 18873 4523 18939 4526
rect 10961 4450 11027 4453
rect 19425 4450 19491 4453
rect 10961 4448 19491 4450
rect 10961 4392 10966 4448
rect 11022 4392 19430 4448
rect 19486 4392 19491 4448
rect 10961 4390 19491 4392
rect 10961 4387 11027 4390
rect 19425 4387 19491 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4521 4314 4587 4317
rect 6637 4314 6703 4317
rect 14641 4316 14707 4317
rect 14590 4314 14596 4316
rect 4521 4312 6703 4314
rect 4521 4256 4526 4312
rect 4582 4256 6642 4312
rect 6698 4256 6703 4312
rect 4521 4254 6703 4256
rect 14514 4254 14596 4314
rect 14660 4314 14707 4316
rect 15101 4314 15167 4317
rect 14660 4312 15167 4314
rect 14702 4256 15106 4312
rect 15162 4256 15167 4312
rect 4521 4251 4587 4254
rect 6637 4251 6703 4254
rect 14590 4252 14596 4254
rect 14660 4254 15167 4256
rect 14660 4252 14707 4254
rect 14641 4251 14707 4252
rect 15101 4251 15167 4254
rect 30281 4314 30347 4317
rect 30925 4314 30991 4317
rect 30281 4312 30991 4314
rect 30281 4256 30286 4312
rect 30342 4256 30930 4312
rect 30986 4256 30991 4312
rect 30281 4254 30991 4256
rect 30281 4251 30347 4254
rect 30925 4251 30991 4254
rect 3601 4178 3667 4181
rect 8937 4178 9003 4181
rect 3601 4176 9003 4178
rect 3601 4120 3606 4176
rect 3662 4120 8942 4176
rect 8998 4120 9003 4176
rect 3601 4118 9003 4120
rect 3601 4115 3667 4118
rect 8937 4115 9003 4118
rect 14089 4178 14155 4181
rect 21449 4178 21515 4181
rect 36813 4178 36879 4181
rect 39200 4178 39800 4208
rect 14089 4176 20730 4178
rect 14089 4120 14094 4176
rect 14150 4120 20730 4176
rect 14089 4118 20730 4120
rect 14089 4115 14155 4118
rect 3969 4042 4035 4045
rect 6361 4042 6427 4045
rect 3969 4040 6427 4042
rect 3969 3984 3974 4040
rect 4030 3984 6366 4040
rect 6422 3984 6427 4040
rect 3969 3982 6427 3984
rect 3969 3979 4035 3982
rect 6361 3979 6427 3982
rect 10777 4042 10843 4045
rect 10910 4042 10916 4044
rect 10777 4040 10916 4042
rect 10777 3984 10782 4040
rect 10838 3984 10916 4040
rect 10777 3982 10916 3984
rect 10777 3979 10843 3982
rect 10910 3980 10916 3982
rect 10980 3980 10986 4044
rect 16297 4042 16363 4045
rect 17166 4042 17172 4044
rect 16297 4040 17172 4042
rect 16297 3984 16302 4040
rect 16358 3984 17172 4040
rect 16297 3982 17172 3984
rect 16297 3979 16363 3982
rect 17166 3980 17172 3982
rect 17236 3980 17242 4044
rect 20670 4042 20730 4118
rect 21449 4176 26250 4178
rect 21449 4120 21454 4176
rect 21510 4120 26250 4176
rect 21449 4118 26250 4120
rect 21449 4115 21515 4118
rect 21398 4042 21404 4044
rect 20670 3982 21404 4042
rect 21398 3980 21404 3982
rect 21468 3980 21474 4044
rect 24577 4042 24643 4045
rect 24710 4042 24716 4044
rect 24577 4040 24716 4042
rect 24577 3984 24582 4040
rect 24638 3984 24716 4040
rect 24577 3982 24716 3984
rect 24577 3979 24643 3982
rect 24710 3980 24716 3982
rect 24780 3980 24786 4044
rect 26190 4042 26250 4118
rect 36813 4176 39800 4178
rect 36813 4120 36818 4176
rect 36874 4120 39800 4176
rect 36813 4118 39800 4120
rect 36813 4115 36879 4118
rect 39200 4088 39800 4118
rect 26550 4042 26556 4044
rect 26190 3982 26556 4042
rect 26550 3980 26556 3982
rect 26620 3980 26626 4044
rect 27521 4042 27587 4045
rect 29177 4042 29243 4045
rect 29310 4042 29316 4044
rect 27521 4040 29316 4042
rect 27521 3984 27526 4040
rect 27582 3984 29182 4040
rect 29238 3984 29316 4040
rect 27521 3982 29316 3984
rect 27521 3979 27587 3982
rect 29177 3979 29243 3982
rect 29310 3980 29316 3982
rect 29380 3980 29386 4044
rect 35617 4042 35683 4045
rect 35750 4042 35756 4044
rect 35617 4040 35756 4042
rect 35617 3984 35622 4040
rect 35678 3984 35756 4040
rect 35617 3982 35756 3984
rect 35617 3979 35683 3982
rect 35750 3980 35756 3982
rect 35820 3980 35826 4044
rect 14406 3844 14412 3908
rect 14476 3906 14482 3908
rect 17493 3906 17559 3909
rect 14476 3904 17559 3906
rect 14476 3848 17498 3904
rect 17554 3848 17559 3904
rect 14476 3846 17559 3848
rect 14476 3844 14482 3846
rect 17493 3843 17559 3846
rect 24209 3906 24275 3909
rect 27889 3906 27955 3909
rect 24209 3904 27955 3906
rect 24209 3848 24214 3904
rect 24270 3848 27894 3904
rect 27950 3848 27955 3904
rect 24209 3846 27955 3848
rect 24209 3843 24275 3846
rect 27889 3843 27955 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 21725 3772 21791 3773
rect 21725 3770 21772 3772
rect 21680 3768 21772 3770
rect 21836 3770 21842 3772
rect 24485 3770 24551 3773
rect 32581 3772 32647 3773
rect 32581 3770 32628 3772
rect 21836 3768 24551 3770
rect 21680 3712 21730 3768
rect 21836 3712 24490 3768
rect 24546 3712 24551 3768
rect 21680 3710 21772 3712
rect 21725 3708 21772 3710
rect 21836 3710 24551 3712
rect 32536 3768 32628 3770
rect 32536 3712 32586 3768
rect 32536 3710 32628 3712
rect 21836 3708 21842 3710
rect 21725 3707 21791 3708
rect 24485 3707 24551 3710
rect 32581 3708 32628 3710
rect 32692 3708 32698 3772
rect 32581 3707 32647 3708
rect 1945 3634 2011 3637
rect 38193 3634 38259 3637
rect 1945 3632 38259 3634
rect 1945 3576 1950 3632
rect 2006 3576 38198 3632
rect 38254 3576 38259 3632
rect 1945 3574 38259 3576
rect 1945 3571 2011 3574
rect 38193 3571 38259 3574
rect 200 3498 800 3528
rect 1761 3498 1827 3501
rect 2221 3500 2287 3501
rect 2221 3498 2268 3500
rect 200 3496 1827 3498
rect 200 3440 1766 3496
rect 1822 3440 1827 3496
rect 200 3438 1827 3440
rect 2176 3496 2268 3498
rect 2176 3440 2226 3496
rect 2176 3438 2268 3440
rect 200 3408 800 3438
rect 1761 3435 1827 3438
rect 2221 3436 2268 3438
rect 2332 3436 2338 3500
rect 3918 3436 3924 3500
rect 3988 3498 3994 3500
rect 7557 3498 7623 3501
rect 3988 3496 7623 3498
rect 3988 3440 7562 3496
rect 7618 3440 7623 3496
rect 3988 3438 7623 3440
rect 3988 3436 3994 3438
rect 2221 3435 2287 3436
rect 7557 3435 7623 3438
rect 8661 3498 8727 3501
rect 35249 3498 35315 3501
rect 8661 3496 35315 3498
rect 8661 3440 8666 3496
rect 8722 3440 35254 3496
rect 35310 3440 35315 3496
rect 8661 3438 35315 3440
rect 8661 3435 8727 3438
rect 35249 3435 35315 3438
rect 38285 3498 38351 3501
rect 39200 3498 39800 3528
rect 38285 3496 39800 3498
rect 38285 3440 38290 3496
rect 38346 3440 39800 3496
rect 38285 3438 39800 3440
rect 38285 3435 38351 3438
rect 39200 3408 39800 3438
rect 5073 3362 5139 3365
rect 7833 3362 7899 3365
rect 5073 3360 7899 3362
rect 5073 3304 5078 3360
rect 5134 3304 7838 3360
rect 7894 3304 7899 3360
rect 5073 3302 7899 3304
rect 5073 3299 5139 3302
rect 7833 3299 7899 3302
rect 16021 3362 16087 3365
rect 19057 3362 19123 3365
rect 16021 3360 19123 3362
rect 16021 3304 16026 3360
rect 16082 3304 19062 3360
rect 19118 3304 19123 3360
rect 16021 3302 19123 3304
rect 16021 3299 16087 3302
rect 19057 3299 19123 3302
rect 22461 3362 22527 3365
rect 27429 3362 27495 3365
rect 22461 3360 27495 3362
rect 22461 3304 22466 3360
rect 22522 3304 27434 3360
rect 27490 3304 27495 3360
rect 22461 3302 27495 3304
rect 22461 3299 22527 3302
rect 27429 3299 27495 3302
rect 34421 3362 34487 3365
rect 38929 3362 38995 3365
rect 34421 3360 38995 3362
rect 34421 3304 34426 3360
rect 34482 3304 38934 3360
rect 38990 3304 38995 3360
rect 34421 3302 38995 3304
rect 34421 3299 34487 3302
rect 38929 3299 38995 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 3969 3226 4035 3229
rect 5942 3226 5948 3228
rect 3969 3224 5948 3226
rect 3969 3168 3974 3224
rect 4030 3168 5948 3224
rect 3969 3166 5948 3168
rect 3969 3163 4035 3166
rect 5942 3164 5948 3166
rect 6012 3226 6018 3228
rect 9397 3226 9463 3229
rect 6012 3224 9463 3226
rect 6012 3168 9402 3224
rect 9458 3168 9463 3224
rect 6012 3166 9463 3168
rect 6012 3164 6018 3166
rect 9397 3163 9463 3166
rect 21265 3226 21331 3229
rect 21398 3226 21404 3228
rect 21265 3224 21404 3226
rect 21265 3168 21270 3224
rect 21326 3168 21404 3224
rect 21265 3166 21404 3168
rect 21265 3163 21331 3166
rect 21398 3164 21404 3166
rect 21468 3164 21474 3228
rect 21817 3226 21883 3229
rect 25221 3226 25287 3229
rect 21817 3224 25287 3226
rect 21817 3168 21822 3224
rect 21878 3168 25226 3224
rect 25282 3168 25287 3224
rect 21817 3166 25287 3168
rect 21817 3163 21883 3166
rect 25221 3163 25287 3166
rect 26417 3226 26483 3229
rect 26550 3226 26556 3228
rect 26417 3224 26556 3226
rect 26417 3168 26422 3224
rect 26478 3168 26556 3224
rect 26417 3166 26556 3168
rect 26417 3163 26483 3166
rect 26550 3164 26556 3166
rect 26620 3164 26626 3228
rect 32581 3090 32647 3093
rect 22050 3088 32647 3090
rect 22050 3032 32586 3088
rect 32642 3032 32647 3088
rect 22050 3030 32647 3032
rect 4797 2954 4863 2957
rect 4981 2954 5047 2957
rect 5993 2954 6059 2957
rect 4797 2952 6059 2954
rect 4797 2896 4802 2952
rect 4858 2896 4986 2952
rect 5042 2896 5998 2952
rect 6054 2896 6059 2952
rect 4797 2894 6059 2896
rect 4797 2891 4863 2894
rect 4981 2891 5047 2894
rect 5993 2891 6059 2894
rect 10777 2954 10843 2957
rect 22050 2954 22110 3030
rect 32581 3027 32647 3030
rect 10777 2952 22110 2954
rect 10777 2896 10782 2952
rect 10838 2896 22110 2952
rect 10777 2894 22110 2896
rect 26969 2954 27035 2957
rect 34789 2954 34855 2957
rect 26969 2952 34855 2954
rect 26969 2896 26974 2952
rect 27030 2896 34794 2952
rect 34850 2896 34855 2952
rect 26969 2894 34855 2896
rect 10777 2891 10843 2894
rect 26969 2891 27035 2894
rect 34789 2891 34855 2894
rect 200 2818 800 2848
rect 1669 2818 1735 2821
rect 200 2816 1735 2818
rect 200 2760 1674 2816
rect 1730 2760 1735 2816
rect 200 2758 1735 2760
rect 200 2728 800 2758
rect 1669 2755 1735 2758
rect 7189 2818 7255 2821
rect 7649 2818 7715 2821
rect 10961 2818 11027 2821
rect 7189 2816 11027 2818
rect 7189 2760 7194 2816
rect 7250 2760 7654 2816
rect 7710 2760 10966 2816
rect 11022 2760 11027 2816
rect 7189 2758 11027 2760
rect 7189 2755 7255 2758
rect 7649 2755 7715 2758
rect 10961 2755 11027 2758
rect 35801 2818 35867 2821
rect 39200 2818 39800 2848
rect 35801 2816 39800 2818
rect 35801 2760 35806 2816
rect 35862 2760 39800 2816
rect 35801 2758 39800 2760
rect 35801 2755 35867 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 2313 2682 2379 2685
rect 3550 2682 3556 2684
rect 2313 2680 3556 2682
rect 2313 2624 2318 2680
rect 2374 2624 3556 2680
rect 2313 2622 3556 2624
rect 2313 2619 2379 2622
rect 3550 2620 3556 2622
rect 3620 2620 3626 2684
rect 16665 2682 16731 2685
rect 24526 2682 24532 2684
rect 16665 2680 24532 2682
rect 16665 2624 16670 2680
rect 16726 2624 24532 2680
rect 16665 2622 24532 2624
rect 16665 2619 16731 2622
rect 24526 2620 24532 2622
rect 24596 2682 24602 2684
rect 29913 2682 29979 2685
rect 24596 2680 29979 2682
rect 24596 2624 29918 2680
rect 29974 2624 29979 2680
rect 24596 2622 29979 2624
rect 24596 2620 24602 2622
rect 29913 2619 29979 2622
rect 4153 2546 4219 2549
rect 4838 2546 4844 2548
rect 4153 2544 4844 2546
rect 4153 2488 4158 2544
rect 4214 2488 4844 2544
rect 4153 2486 4844 2488
rect 4153 2483 4219 2486
rect 4838 2484 4844 2486
rect 4908 2484 4914 2548
rect 31293 2546 31359 2549
rect 31702 2546 31708 2548
rect 31293 2544 31708 2546
rect 31293 2488 31298 2544
rect 31354 2488 31708 2544
rect 31293 2486 31708 2488
rect 31293 2483 31359 2486
rect 31702 2484 31708 2486
rect 31772 2484 31778 2548
rect 27429 2410 27495 2413
rect 36118 2410 36124 2412
rect 27429 2408 36124 2410
rect 27429 2352 27434 2408
rect 27490 2352 36124 2408
rect 27429 2350 36124 2352
rect 27429 2347 27495 2350
rect 36118 2348 36124 2350
rect 36188 2348 36194 2412
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1485 1458 1551 1461
rect 200 1456 1551 1458
rect 200 1400 1490 1456
rect 1546 1400 1551 1456
rect 200 1398 1551 1400
rect 200 1368 800 1398
rect 1485 1395 1551 1398
rect 35709 1458 35775 1461
rect 39200 1458 39800 1488
rect 35709 1456 39800 1458
rect 35709 1400 35714 1456
rect 35770 1400 39800 1456
rect 35709 1398 39800 1400
rect 35709 1395 35775 1398
rect 39200 1368 39800 1398
rect 200 778 800 808
rect 1853 778 1919 781
rect 200 776 1919 778
rect 200 720 1858 776
rect 1914 720 1919 776
rect 200 718 1919 720
rect 200 688 800 718
rect 1853 715 1919 718
rect 37549 778 37615 781
rect 39200 778 39800 808
rect 37549 776 39800 778
rect 37549 720 37554 776
rect 37610 720 39800 776
rect 37549 718 39800 720
rect 37549 715 37615 718
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 24164 32540 24228 32604
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4844 30092 4908 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 9076 29684 9140 29748
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 23428 27644 23492 27708
rect 8524 27296 8588 27300
rect 8524 27240 8538 27296
rect 8538 27240 8588 27296
rect 8524 27236 8588 27240
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 20300 25332 20364 25396
rect 20484 25196 20548 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 17540 24924 17604 24988
rect 12020 24788 12084 24852
rect 18460 24712 18524 24716
rect 18460 24656 18474 24712
rect 18474 24656 18524 24712
rect 18460 24652 18524 24656
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 1900 23428 1964 23492
rect 18276 23428 18340 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 22876 23700 22940 23764
rect 23612 23564 23676 23628
rect 30052 23488 30116 23492
rect 30052 23432 30102 23488
rect 30102 23432 30116 23488
rect 30052 23428 30116 23432
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 36860 23020 36924 23084
rect 26924 22884 26988 22948
rect 28212 22884 28276 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 20116 22612 20180 22676
rect 31524 22536 31588 22540
rect 31524 22480 31538 22536
rect 31538 22480 31588 22536
rect 31524 22476 31588 22480
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 22692 21992 22756 21996
rect 22692 21936 22742 21992
rect 22742 21936 22756 21992
rect 22692 21932 22756 21936
rect 32260 21796 32324 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 11836 21388 11900 21452
rect 21404 21388 21468 21452
rect 27660 21388 27724 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 17172 21116 17236 21180
rect 28212 20844 28276 20908
rect 13492 20708 13556 20772
rect 21956 20768 22020 20772
rect 21956 20712 22006 20768
rect 22006 20712 22020 20768
rect 21956 20708 22020 20712
rect 23428 20708 23492 20772
rect 24716 20708 24780 20772
rect 25268 20708 25332 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 22140 20436 22204 20500
rect 21036 20300 21100 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 5396 19756 5460 19820
rect 32444 19756 32508 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 17356 19408 17420 19412
rect 17356 19352 17370 19408
rect 17370 19352 17420 19408
rect 17356 19348 17420 19352
rect 31892 19348 31956 19412
rect 32076 19348 32140 19412
rect 3556 19212 3620 19276
rect 13492 19076 13556 19140
rect 17724 19076 17788 19140
rect 25820 19076 25884 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 5028 18668 5092 18732
rect 29132 18668 29196 18732
rect 17540 18532 17604 18596
rect 28580 18532 28644 18596
rect 28764 18592 28828 18596
rect 28764 18536 28778 18592
rect 28778 18536 28828 18592
rect 28764 18532 28828 18536
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 27476 18260 27540 18324
rect 25636 18124 25700 18188
rect 26372 18124 26436 18188
rect 28948 18124 29012 18188
rect 30420 18124 30484 18188
rect 9444 18048 9508 18052
rect 9444 17992 9494 18048
rect 9494 17992 9508 18048
rect 9444 17988 9508 17992
rect 20668 17988 20732 18052
rect 25084 17988 25148 18052
rect 26556 17988 26620 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 7604 17852 7668 17916
rect 28948 17912 29012 17916
rect 28948 17856 28962 17912
rect 28962 17856 29012 17912
rect 28948 17852 29012 17856
rect 10732 17580 10796 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 28764 17308 28828 17372
rect 32628 17308 32692 17372
rect 13492 17172 13556 17236
rect 7788 17036 7852 17100
rect 12940 16900 13004 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 16436 16764 16500 16828
rect 9260 16628 9324 16692
rect 14596 16628 14660 16692
rect 14964 16628 15028 16692
rect 16068 16628 16132 16692
rect 18644 16688 18708 16692
rect 18644 16632 18658 16688
rect 18658 16632 18708 16688
rect 18644 16628 18708 16632
rect 11100 16492 11164 16556
rect 15148 16492 15212 16556
rect 19380 16492 19444 16556
rect 33180 16628 33244 16692
rect 9996 16356 10060 16420
rect 33732 16552 33796 16556
rect 33732 16496 33782 16552
rect 33782 16496 33796 16552
rect 33732 16492 33796 16496
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 24164 16280 24228 16284
rect 24164 16224 24178 16280
rect 24178 16224 24228 16280
rect 24164 16220 24228 16224
rect 10916 15948 10980 16012
rect 12756 15948 12820 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 28396 15676 28460 15740
rect 32076 15676 32140 15740
rect 13676 15404 13740 15468
rect 23060 15540 23124 15604
rect 16252 15328 16316 15332
rect 16252 15272 16266 15328
rect 16266 15272 16316 15328
rect 16252 15268 16316 15272
rect 24532 15268 24596 15332
rect 28948 15268 29012 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 13124 15132 13188 15196
rect 13492 15132 13556 15196
rect 6500 14996 6564 15060
rect 21772 14996 21836 15060
rect 9812 14920 9876 14924
rect 9812 14864 9826 14920
rect 9826 14864 9876 14920
rect 9812 14860 9876 14864
rect 16804 14724 16868 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 17724 14452 17788 14516
rect 33180 14588 33244 14652
rect 27476 14316 27540 14380
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 20852 14044 20916 14108
rect 14412 13908 14476 13972
rect 5212 13636 5276 13700
rect 9076 13636 9140 13700
rect 17356 13696 17420 13700
rect 17356 13640 17406 13696
rect 17406 13640 17420 13696
rect 17356 13636 17420 13640
rect 20300 13636 20364 13700
rect 27660 13636 27724 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 13676 13560 13740 13564
rect 13676 13504 13690 13560
rect 13690 13504 13740 13560
rect 13676 13500 13740 13504
rect 14228 13500 14292 13564
rect 16620 13500 16684 13564
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 22876 13500 22940 13564
rect 12204 13364 12268 13428
rect 7052 13228 7116 13292
rect 23060 13364 23124 13428
rect 20116 13228 20180 13292
rect 17908 13092 17972 13156
rect 30788 13092 30852 13156
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 22508 12956 22572 13020
rect 9076 12880 9140 12884
rect 9076 12824 9126 12880
rect 9126 12824 9140 12880
rect 9076 12820 9140 12824
rect 22140 12820 22204 12884
rect 35756 12820 35820 12884
rect 24900 12684 24964 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 2268 12412 2332 12476
rect 6684 12412 6748 12476
rect 9996 12412 10060 12476
rect 20300 12608 20364 12612
rect 20300 12552 20350 12608
rect 20350 12552 20364 12608
rect 20300 12548 20364 12552
rect 22140 12548 22204 12612
rect 32260 12548 32324 12612
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 28580 12472 28644 12476
rect 28580 12416 28630 12472
rect 28630 12416 28644 12472
rect 28580 12412 28644 12416
rect 1900 12276 1964 12340
rect 18460 12276 18524 12340
rect 25268 12336 25332 12340
rect 32444 12412 32508 12476
rect 25268 12280 25318 12336
rect 25318 12280 25332 12336
rect 25268 12276 25332 12280
rect 27476 12276 27540 12340
rect 29316 12276 29380 12340
rect 9444 12004 9508 12068
rect 11836 12140 11900 12204
rect 18276 12140 18340 12204
rect 31524 12140 31588 12204
rect 9260 11928 9324 11932
rect 9260 11872 9310 11928
rect 9310 11872 9324 11928
rect 9260 11868 9324 11872
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 8708 11596 8772 11660
rect 9812 11596 9876 11660
rect 10548 11656 10612 11660
rect 10548 11600 10598 11656
rect 10598 11600 10612 11656
rect 10548 11596 10612 11600
rect 22692 11732 22756 11796
rect 30052 11732 30116 11796
rect 20668 11656 20732 11660
rect 20668 11600 20682 11656
rect 20682 11600 20732 11656
rect 20668 11596 20732 11600
rect 26556 11596 26620 11660
rect 28948 11596 29012 11660
rect 30420 11596 30484 11660
rect 31524 11596 31588 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 8340 11052 8404 11116
rect 9996 11112 10060 11116
rect 9996 11056 10046 11112
rect 10046 11056 10060 11112
rect 9996 11052 10060 11056
rect 18460 11460 18524 11524
rect 22324 11460 22388 11524
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 26372 11052 26436 11116
rect 36124 11112 36188 11116
rect 36124 11056 36138 11112
rect 36138 11056 36188 11112
rect 12940 10916 13004 10980
rect 14228 10916 14292 10980
rect 20484 10976 20548 10980
rect 36124 11052 36188 11056
rect 20484 10920 20498 10976
rect 20498 10920 20548 10976
rect 20484 10916 20548 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 15884 10780 15948 10844
rect 16436 10780 16500 10844
rect 29132 10916 29196 10980
rect 11100 10644 11164 10708
rect 16436 10644 16500 10708
rect 20300 10704 20364 10708
rect 20300 10648 20350 10704
rect 20350 10648 20364 10704
rect 20300 10644 20364 10648
rect 25820 10508 25884 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 5764 10024 5828 10028
rect 5764 9968 5814 10024
rect 5814 9968 5828 10024
rect 5764 9964 5828 9968
rect 12020 10024 12084 10028
rect 12020 9968 12034 10024
rect 12034 9968 12084 10024
rect 12020 9964 12084 9968
rect 19380 9828 19444 9892
rect 20852 9828 20916 9892
rect 26740 9888 26804 9892
rect 26740 9832 26790 9888
rect 26790 9832 26804 9888
rect 26740 9828 26804 9832
rect 28948 9828 29012 9892
rect 30604 9828 30668 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 5948 9616 6012 9620
rect 5948 9560 5962 9616
rect 5962 9560 6012 9616
rect 5948 9556 6012 9560
rect 10732 9692 10796 9756
rect 16252 9692 16316 9756
rect 18644 9752 18708 9756
rect 18644 9696 18658 9752
rect 18658 9696 18708 9752
rect 18644 9692 18708 9696
rect 26924 9692 26988 9756
rect 6684 9556 6748 9620
rect 6868 9556 6932 9620
rect 10548 9616 10612 9620
rect 10548 9560 10562 9616
rect 10562 9560 10612 9616
rect 10548 9556 10612 9560
rect 22140 9556 22204 9620
rect 21036 9420 21100 9484
rect 23612 9420 23676 9484
rect 14964 9284 15028 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 6316 9148 6380 9212
rect 25084 9148 25148 9212
rect 5396 8876 5460 8940
rect 17724 8876 17788 8940
rect 30788 8876 30852 8940
rect 32076 8876 32140 8940
rect 3924 8740 3988 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 6316 8528 6380 8532
rect 6316 8472 6366 8528
rect 6366 8472 6380 8528
rect 6316 8468 6380 8472
rect 16620 8468 16684 8532
rect 30420 8468 30484 8532
rect 30788 8468 30852 8532
rect 16804 8332 16868 8396
rect 17908 8332 17972 8396
rect 24900 8332 24964 8396
rect 22324 8256 22388 8260
rect 22324 8200 22338 8256
rect 22338 8200 22388 8256
rect 22324 8196 22388 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 16436 8060 16500 8124
rect 30420 7924 30484 7988
rect 22508 7788 22572 7852
rect 5028 7652 5092 7716
rect 27476 7712 27540 7716
rect 27476 7656 27490 7712
rect 27490 7656 27540 7712
rect 27476 7652 27540 7656
rect 32076 7652 32140 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 14596 7244 14660 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 5212 6836 5276 6900
rect 7788 6896 7852 6900
rect 7788 6840 7838 6896
rect 7838 6840 7852 6896
rect 7788 6836 7852 6840
rect 8340 6836 8404 6900
rect 8708 6896 8772 6900
rect 8708 6840 8758 6896
rect 8758 6840 8772 6896
rect 8708 6836 8772 6840
rect 6868 6700 6932 6764
rect 8524 6700 8588 6764
rect 12572 6896 12636 6900
rect 12572 6840 12622 6896
rect 12622 6840 12636 6896
rect 12572 6836 12636 6840
rect 13124 6896 13188 6900
rect 13124 6840 13138 6896
rect 13138 6840 13188 6896
rect 13124 6836 13188 6840
rect 21956 6836 22020 6900
rect 25636 6896 25700 6900
rect 31524 7032 31588 7036
rect 31524 6976 31574 7032
rect 31574 6976 31588 7032
rect 31524 6972 31588 6976
rect 25636 6840 25650 6896
rect 25650 6840 25700 6896
rect 25636 6836 25700 6840
rect 30420 6836 30484 6900
rect 9628 6564 9692 6628
rect 30788 6564 30852 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 27476 6488 27540 6492
rect 27476 6432 27490 6488
rect 27490 6432 27540 6488
rect 27476 6428 27540 6432
rect 5764 6292 5828 6356
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 1900 5944 1964 5948
rect 1900 5888 1914 5944
rect 1914 5888 1964 5944
rect 1900 5884 1964 5888
rect 12756 5748 12820 5812
rect 28212 5808 28276 5812
rect 28212 5752 28262 5808
rect 28262 5752 28276 5808
rect 28212 5748 28276 5752
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 6500 5612 6564 5676
rect 6868 5612 6932 5676
rect 7052 5536 7116 5540
rect 7052 5480 7066 5536
rect 7066 5480 7116 5536
rect 7052 5476 7116 5480
rect 7604 5536 7668 5540
rect 7604 5480 7618 5536
rect 7618 5480 7668 5536
rect 7604 5476 7668 5480
rect 16068 5536 16132 5540
rect 16068 5480 16118 5536
rect 16118 5480 16132 5536
rect 16068 5476 16132 5480
rect 28396 5476 28460 5540
rect 33732 5476 33796 5540
rect 36860 5476 36924 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 15148 5400 15212 5404
rect 15148 5344 15162 5400
rect 15162 5344 15212 5400
rect 15148 5340 15212 5344
rect 15884 5340 15948 5404
rect 28948 5068 29012 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 14596 4312 14660 4316
rect 14596 4256 14646 4312
rect 14646 4256 14660 4312
rect 14596 4252 14660 4256
rect 10916 3980 10980 4044
rect 17172 3980 17236 4044
rect 21404 3980 21468 4044
rect 24716 3980 24780 4044
rect 26556 3980 26620 4044
rect 29316 3980 29380 4044
rect 35756 3980 35820 4044
rect 14412 3844 14476 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 21772 3768 21836 3772
rect 21772 3712 21786 3768
rect 21786 3712 21836 3768
rect 21772 3708 21836 3712
rect 32628 3768 32692 3772
rect 32628 3712 32642 3768
rect 32642 3712 32692 3768
rect 32628 3708 32692 3712
rect 2268 3496 2332 3500
rect 2268 3440 2282 3496
rect 2282 3440 2332 3496
rect 2268 3436 2332 3440
rect 3924 3436 3988 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 5948 3164 6012 3228
rect 21404 3164 21468 3228
rect 26556 3164 26620 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 3556 2620 3620 2684
rect 24532 2620 24596 2684
rect 4844 2484 4908 2548
rect 31708 2484 31772 2548
rect 36124 2348 36188 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 24163 32604 24229 32605
rect 24163 32540 24164 32604
rect 24228 32540 24229 32604
rect 24163 32539 24229 32540
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 4843 30156 4909 30157
rect 4843 30092 4844 30156
rect 4908 30092 4909 30156
rect 4843 30091 4909 30092
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 1899 23492 1965 23493
rect 1899 23428 1900 23492
rect 1964 23428 1965 23492
rect 1899 23427 1965 23428
rect 1902 12341 1962 23427
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3555 19276 3621 19277
rect 3555 19212 3556 19276
rect 3620 19212 3621 19276
rect 3555 19211 3621 19212
rect 2267 12476 2333 12477
rect 2267 12412 2268 12476
rect 2332 12412 2333 12476
rect 2267 12411 2333 12412
rect 1899 12340 1965 12341
rect 1899 12276 1900 12340
rect 1964 12276 1965 12340
rect 1899 12275 1965 12276
rect 1902 5949 1962 12275
rect 1899 5948 1965 5949
rect 1899 5884 1900 5948
rect 1964 5884 1965 5948
rect 1899 5883 1965 5884
rect 2270 3501 2330 12411
rect 2267 3500 2333 3501
rect 2267 3436 2268 3500
rect 2332 3436 2333 3500
rect 2267 3435 2333 3436
rect 3558 2685 3618 19211
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 3923 8804 3989 8805
rect 3923 8740 3924 8804
rect 3988 8740 3989 8804
rect 3923 8739 3989 8740
rect 3926 3501 3986 8739
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 3923 3500 3989 3501
rect 3923 3436 3924 3500
rect 3988 3436 3989 3500
rect 3923 3435 3989 3436
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 3555 2684 3621 2685
rect 3555 2620 3556 2684
rect 3620 2620 3621 2684
rect 3555 2619 3621 2620
rect 4208 2128 4528 2688
rect 4846 2549 4906 30091
rect 9075 29748 9141 29749
rect 9075 29684 9076 29748
rect 9140 29684 9141 29748
rect 9075 29683 9141 29684
rect 8523 27300 8589 27301
rect 8523 27236 8524 27300
rect 8588 27236 8589 27300
rect 8523 27235 8589 27236
rect 5395 19820 5461 19821
rect 5395 19756 5396 19820
rect 5460 19756 5461 19820
rect 5395 19755 5461 19756
rect 5027 18732 5093 18733
rect 5027 18668 5028 18732
rect 5092 18668 5093 18732
rect 5027 18667 5093 18668
rect 5030 7717 5090 18667
rect 5211 13700 5277 13701
rect 5211 13636 5212 13700
rect 5276 13636 5277 13700
rect 5211 13635 5277 13636
rect 5027 7716 5093 7717
rect 5027 7652 5028 7716
rect 5092 7652 5093 7716
rect 5027 7651 5093 7652
rect 5214 6901 5274 13635
rect 5398 8941 5458 19755
rect 7603 17916 7669 17917
rect 7603 17852 7604 17916
rect 7668 17852 7669 17916
rect 7603 17851 7669 17852
rect 6499 15060 6565 15061
rect 6499 14996 6500 15060
rect 6564 14996 6565 15060
rect 6499 14995 6565 14996
rect 5763 10028 5829 10029
rect 5763 9964 5764 10028
rect 5828 9964 5829 10028
rect 5763 9963 5829 9964
rect 5395 8940 5461 8941
rect 5395 8876 5396 8940
rect 5460 8876 5461 8940
rect 5395 8875 5461 8876
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 5766 6357 5826 9963
rect 5947 9620 6013 9621
rect 5947 9556 5948 9620
rect 6012 9556 6013 9620
rect 5947 9555 6013 9556
rect 5763 6356 5829 6357
rect 5763 6292 5764 6356
rect 5828 6292 5829 6356
rect 5763 6291 5829 6292
rect 5950 3229 6010 9555
rect 6315 9212 6381 9213
rect 6315 9148 6316 9212
rect 6380 9148 6381 9212
rect 6315 9147 6381 9148
rect 6318 8533 6378 9147
rect 6315 8532 6381 8533
rect 6315 8468 6316 8532
rect 6380 8468 6381 8532
rect 6315 8467 6381 8468
rect 6502 5677 6562 14995
rect 7051 13292 7117 13293
rect 7051 13228 7052 13292
rect 7116 13228 7117 13292
rect 7051 13227 7117 13228
rect 6683 12476 6749 12477
rect 6683 12412 6684 12476
rect 6748 12412 6749 12476
rect 6683 12411 6749 12412
rect 6686 9621 6746 12411
rect 6683 9620 6749 9621
rect 6683 9556 6684 9620
rect 6748 9556 6749 9620
rect 6683 9555 6749 9556
rect 6867 9620 6933 9621
rect 6867 9556 6868 9620
rect 6932 9556 6933 9620
rect 6867 9555 6933 9556
rect 6870 6765 6930 9555
rect 6867 6764 6933 6765
rect 6867 6700 6868 6764
rect 6932 6700 6933 6764
rect 6867 6699 6933 6700
rect 6870 5677 6930 6699
rect 6499 5676 6565 5677
rect 6499 5612 6500 5676
rect 6564 5612 6565 5676
rect 6499 5611 6565 5612
rect 6867 5676 6933 5677
rect 6867 5612 6868 5676
rect 6932 5612 6933 5676
rect 6867 5611 6933 5612
rect 7054 5541 7114 13227
rect 7606 5541 7666 17851
rect 7787 17100 7853 17101
rect 7787 17036 7788 17100
rect 7852 17036 7853 17100
rect 7787 17035 7853 17036
rect 7790 6901 7850 17035
rect 8339 11116 8405 11117
rect 8339 11052 8340 11116
rect 8404 11052 8405 11116
rect 8339 11051 8405 11052
rect 8342 6901 8402 11051
rect 7787 6900 7853 6901
rect 7787 6836 7788 6900
rect 7852 6836 7853 6900
rect 7787 6835 7853 6836
rect 8339 6900 8405 6901
rect 8339 6836 8340 6900
rect 8404 6836 8405 6900
rect 8339 6835 8405 6836
rect 8526 6765 8586 27235
rect 9078 13701 9138 29683
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 23427 27708 23493 27709
rect 23427 27644 23428 27708
rect 23492 27644 23493 27708
rect 23427 27643 23493 27644
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 20299 25396 20365 25397
rect 20299 25332 20300 25396
rect 20364 25332 20365 25396
rect 20299 25331 20365 25332
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 17539 24988 17605 24989
rect 17539 24924 17540 24988
rect 17604 24924 17605 24988
rect 17539 24923 17605 24924
rect 12019 24852 12085 24853
rect 12019 24788 12020 24852
rect 12084 24788 12085 24852
rect 12019 24787 12085 24788
rect 11835 21452 11901 21453
rect 11835 21388 11836 21452
rect 11900 21388 11901 21452
rect 11835 21387 11901 21388
rect 9443 18052 9509 18053
rect 9443 17988 9444 18052
rect 9508 17988 9509 18052
rect 9443 17987 9509 17988
rect 9259 16692 9325 16693
rect 9259 16628 9260 16692
rect 9324 16628 9325 16692
rect 9259 16627 9325 16628
rect 9075 13700 9141 13701
rect 9075 13636 9076 13700
rect 9140 13636 9141 13700
rect 9075 13635 9141 13636
rect 9078 12885 9138 13635
rect 9075 12884 9141 12885
rect 9075 12820 9076 12884
rect 9140 12820 9141 12884
rect 9075 12819 9141 12820
rect 9262 11933 9322 16627
rect 9446 12069 9506 17987
rect 10731 17644 10797 17645
rect 10731 17580 10732 17644
rect 10796 17580 10797 17644
rect 10731 17579 10797 17580
rect 9995 16420 10061 16421
rect 9995 16356 9996 16420
rect 10060 16356 10061 16420
rect 9995 16355 10061 16356
rect 9811 14924 9877 14925
rect 9811 14860 9812 14924
rect 9876 14860 9877 14924
rect 9811 14859 9877 14860
rect 9443 12068 9509 12069
rect 9443 12004 9444 12068
rect 9508 12004 9509 12068
rect 9443 12003 9509 12004
rect 9259 11932 9325 11933
rect 9259 11868 9260 11932
rect 9324 11868 9325 11932
rect 9259 11867 9325 11868
rect 9814 11661 9874 14859
rect 9998 12477 10058 16355
rect 9995 12476 10061 12477
rect 9995 12412 9996 12476
rect 10060 12412 10061 12476
rect 9995 12411 10061 12412
rect 8707 11660 8773 11661
rect 8707 11596 8708 11660
rect 8772 11596 8773 11660
rect 8707 11595 8773 11596
rect 9811 11660 9877 11661
rect 9811 11596 9812 11660
rect 9876 11596 9877 11660
rect 9811 11595 9877 11596
rect 8710 6901 8770 11595
rect 9814 9690 9874 11595
rect 9998 11117 10058 12411
rect 10547 11660 10613 11661
rect 10547 11596 10548 11660
rect 10612 11596 10613 11660
rect 10547 11595 10613 11596
rect 9995 11116 10061 11117
rect 9995 11052 9996 11116
rect 10060 11052 10061 11116
rect 9995 11051 10061 11052
rect 9630 9630 9874 9690
rect 8707 6900 8773 6901
rect 8707 6836 8708 6900
rect 8772 6836 8773 6900
rect 8707 6835 8773 6836
rect 8523 6764 8589 6765
rect 8523 6700 8524 6764
rect 8588 6700 8589 6764
rect 8523 6699 8589 6700
rect 9630 6629 9690 9630
rect 10550 9621 10610 11595
rect 10734 9757 10794 17579
rect 11099 16556 11165 16557
rect 11099 16492 11100 16556
rect 11164 16492 11165 16556
rect 11099 16491 11165 16492
rect 10915 16012 10981 16013
rect 10915 15948 10916 16012
rect 10980 15948 10981 16012
rect 10915 15947 10981 15948
rect 10731 9756 10797 9757
rect 10731 9692 10732 9756
rect 10796 9692 10797 9756
rect 10731 9691 10797 9692
rect 10547 9620 10613 9621
rect 10547 9556 10548 9620
rect 10612 9556 10613 9620
rect 10547 9555 10613 9556
rect 9627 6628 9693 6629
rect 9627 6564 9628 6628
rect 9692 6564 9693 6628
rect 9627 6563 9693 6564
rect 7051 5540 7117 5541
rect 7051 5476 7052 5540
rect 7116 5476 7117 5540
rect 7051 5475 7117 5476
rect 7603 5540 7669 5541
rect 7603 5476 7604 5540
rect 7668 5476 7669 5540
rect 7603 5475 7669 5476
rect 10918 4045 10978 15947
rect 11102 10709 11162 16491
rect 11838 12205 11898 21387
rect 11835 12204 11901 12205
rect 11835 12140 11836 12204
rect 11900 12140 11901 12204
rect 11835 12139 11901 12140
rect 11099 10708 11165 10709
rect 11099 10644 11100 10708
rect 11164 10644 11165 10708
rect 11099 10643 11165 10644
rect 12022 10029 12082 24787
rect 17171 21180 17237 21181
rect 17171 21116 17172 21180
rect 17236 21116 17237 21180
rect 17171 21115 17237 21116
rect 13491 20772 13557 20773
rect 13491 20708 13492 20772
rect 13556 20708 13557 20772
rect 13491 20707 13557 20708
rect 13494 19141 13554 20707
rect 13491 19140 13557 19141
rect 13491 19076 13492 19140
rect 13556 19076 13557 19140
rect 13491 19075 13557 19076
rect 13491 17236 13557 17237
rect 13491 17172 13492 17236
rect 13556 17172 13557 17236
rect 13491 17171 13557 17172
rect 12939 16964 13005 16965
rect 12939 16900 12940 16964
rect 13004 16900 13005 16964
rect 12939 16899 13005 16900
rect 12755 16012 12821 16013
rect 12755 15948 12756 16012
rect 12820 15948 12821 16012
rect 12755 15947 12821 15948
rect 12203 13428 12269 13429
rect 12203 13364 12204 13428
rect 12268 13364 12269 13428
rect 12203 13363 12269 13364
rect 12019 10028 12085 10029
rect 12019 9964 12020 10028
rect 12084 9964 12085 10028
rect 12019 9963 12085 9964
rect 12206 9690 12266 13363
rect 12206 9630 12634 9690
rect 12574 6901 12634 9630
rect 12571 6900 12637 6901
rect 12571 6836 12572 6900
rect 12636 6836 12637 6900
rect 12571 6835 12637 6836
rect 12758 5813 12818 15947
rect 12942 10981 13002 16899
rect 13494 15197 13554 17171
rect 16435 16828 16501 16829
rect 16435 16764 16436 16828
rect 16500 16764 16501 16828
rect 16435 16763 16501 16764
rect 14595 16692 14661 16693
rect 14595 16628 14596 16692
rect 14660 16628 14661 16692
rect 14595 16627 14661 16628
rect 14963 16692 15029 16693
rect 14963 16628 14964 16692
rect 15028 16628 15029 16692
rect 14963 16627 15029 16628
rect 16067 16692 16133 16693
rect 16067 16628 16068 16692
rect 16132 16628 16133 16692
rect 16067 16627 16133 16628
rect 13675 15468 13741 15469
rect 13675 15404 13676 15468
rect 13740 15404 13741 15468
rect 13675 15403 13741 15404
rect 13123 15196 13189 15197
rect 13123 15132 13124 15196
rect 13188 15132 13189 15196
rect 13123 15131 13189 15132
rect 13491 15196 13557 15197
rect 13491 15132 13492 15196
rect 13556 15132 13557 15196
rect 13491 15131 13557 15132
rect 12939 10980 13005 10981
rect 12939 10916 12940 10980
rect 13004 10916 13005 10980
rect 12939 10915 13005 10916
rect 13126 6901 13186 15131
rect 13678 13565 13738 15403
rect 14411 13972 14477 13973
rect 14411 13908 14412 13972
rect 14476 13908 14477 13972
rect 14411 13907 14477 13908
rect 13675 13564 13741 13565
rect 13675 13500 13676 13564
rect 13740 13500 13741 13564
rect 13675 13499 13741 13500
rect 14227 13564 14293 13565
rect 14227 13500 14228 13564
rect 14292 13500 14293 13564
rect 14227 13499 14293 13500
rect 14230 10981 14290 13499
rect 14227 10980 14293 10981
rect 14227 10916 14228 10980
rect 14292 10916 14293 10980
rect 14227 10915 14293 10916
rect 13123 6900 13189 6901
rect 13123 6836 13124 6900
rect 13188 6836 13189 6900
rect 13123 6835 13189 6836
rect 12755 5812 12821 5813
rect 12755 5748 12756 5812
rect 12820 5748 12821 5812
rect 12755 5747 12821 5748
rect 10915 4044 10981 4045
rect 10915 3980 10916 4044
rect 10980 3980 10981 4044
rect 10915 3979 10981 3980
rect 14414 3909 14474 13907
rect 14598 7309 14658 16627
rect 14966 9349 15026 16627
rect 15147 16556 15213 16557
rect 15147 16492 15148 16556
rect 15212 16492 15213 16556
rect 15147 16491 15213 16492
rect 14963 9348 15029 9349
rect 14963 9284 14964 9348
rect 15028 9284 15029 9348
rect 14963 9283 15029 9284
rect 14595 7308 14661 7309
rect 14595 7244 14596 7308
rect 14660 7244 14661 7308
rect 14595 7243 14661 7244
rect 14598 4317 14658 7243
rect 15150 5405 15210 16491
rect 15883 10844 15949 10845
rect 15883 10780 15884 10844
rect 15948 10780 15949 10844
rect 15883 10779 15949 10780
rect 15886 5405 15946 10779
rect 16070 5541 16130 16627
rect 16251 15332 16317 15333
rect 16251 15268 16252 15332
rect 16316 15268 16317 15332
rect 16251 15267 16317 15268
rect 16254 9757 16314 15267
rect 16438 10845 16498 16763
rect 16803 14788 16869 14789
rect 16803 14724 16804 14788
rect 16868 14724 16869 14788
rect 16803 14723 16869 14724
rect 16619 13564 16685 13565
rect 16619 13500 16620 13564
rect 16684 13500 16685 13564
rect 16619 13499 16685 13500
rect 16435 10844 16501 10845
rect 16435 10780 16436 10844
rect 16500 10780 16501 10844
rect 16435 10779 16501 10780
rect 16435 10708 16501 10709
rect 16435 10644 16436 10708
rect 16500 10644 16501 10708
rect 16435 10643 16501 10644
rect 16251 9756 16317 9757
rect 16251 9692 16252 9756
rect 16316 9692 16317 9756
rect 16251 9691 16317 9692
rect 16438 8125 16498 10643
rect 16622 8533 16682 13499
rect 16619 8532 16685 8533
rect 16619 8468 16620 8532
rect 16684 8468 16685 8532
rect 16619 8467 16685 8468
rect 16806 8397 16866 14723
rect 16803 8396 16869 8397
rect 16803 8332 16804 8396
rect 16868 8332 16869 8396
rect 16803 8331 16869 8332
rect 16435 8124 16501 8125
rect 16435 8060 16436 8124
rect 16500 8060 16501 8124
rect 16435 8059 16501 8060
rect 16067 5540 16133 5541
rect 16067 5476 16068 5540
rect 16132 5476 16133 5540
rect 16067 5475 16133 5476
rect 15147 5404 15213 5405
rect 15147 5340 15148 5404
rect 15212 5340 15213 5404
rect 15147 5339 15213 5340
rect 15883 5404 15949 5405
rect 15883 5340 15884 5404
rect 15948 5340 15949 5404
rect 15883 5339 15949 5340
rect 14595 4316 14661 4317
rect 14595 4252 14596 4316
rect 14660 4252 14661 4316
rect 14595 4251 14661 4252
rect 17174 4045 17234 21115
rect 17355 19412 17421 19413
rect 17355 19348 17356 19412
rect 17420 19348 17421 19412
rect 17355 19347 17421 19348
rect 17358 13701 17418 19347
rect 17542 18597 17602 24923
rect 18459 24716 18525 24717
rect 18459 24652 18460 24716
rect 18524 24652 18525 24716
rect 18459 24651 18525 24652
rect 18275 23492 18341 23493
rect 18275 23428 18276 23492
rect 18340 23428 18341 23492
rect 18275 23427 18341 23428
rect 17723 19140 17789 19141
rect 17723 19076 17724 19140
rect 17788 19076 17789 19140
rect 17723 19075 17789 19076
rect 17539 18596 17605 18597
rect 17539 18532 17540 18596
rect 17604 18532 17605 18596
rect 17539 18531 17605 18532
rect 17726 14517 17786 19075
rect 17723 14516 17789 14517
rect 17723 14452 17724 14516
rect 17788 14452 17789 14516
rect 17723 14451 17789 14452
rect 17355 13700 17421 13701
rect 17355 13636 17356 13700
rect 17420 13636 17421 13700
rect 17355 13635 17421 13636
rect 17726 8941 17786 14451
rect 17907 13156 17973 13157
rect 17907 13092 17908 13156
rect 17972 13092 17973 13156
rect 17907 13091 17973 13092
rect 17723 8940 17789 8941
rect 17723 8876 17724 8940
rect 17788 8876 17789 8940
rect 17723 8875 17789 8876
rect 17910 8397 17970 13091
rect 18278 12205 18338 23427
rect 18462 12341 18522 24651
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 20115 22676 20181 22677
rect 20115 22612 20116 22676
rect 20180 22612 20181 22676
rect 20115 22611 20181 22612
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 18643 16692 18709 16693
rect 18643 16628 18644 16692
rect 18708 16628 18709 16692
rect 18643 16627 18709 16628
rect 18459 12340 18525 12341
rect 18459 12276 18460 12340
rect 18524 12276 18525 12340
rect 18459 12275 18525 12276
rect 18275 12204 18341 12205
rect 18275 12140 18276 12204
rect 18340 12140 18341 12204
rect 18275 12139 18341 12140
rect 18462 11525 18522 12275
rect 18459 11524 18525 11525
rect 18459 11460 18460 11524
rect 18524 11460 18525 11524
rect 18459 11459 18525 11460
rect 18646 9757 18706 16627
rect 19379 16556 19445 16557
rect 19379 16492 19380 16556
rect 19444 16492 19445 16556
rect 19379 16491 19445 16492
rect 19382 9893 19442 16491
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 20118 13293 20178 22611
rect 20302 13701 20362 25331
rect 20483 25260 20549 25261
rect 20483 25196 20484 25260
rect 20548 25196 20549 25260
rect 20483 25195 20549 25196
rect 20299 13700 20365 13701
rect 20299 13636 20300 13700
rect 20364 13636 20365 13700
rect 20299 13635 20365 13636
rect 20115 13292 20181 13293
rect 20115 13228 20116 13292
rect 20180 13228 20181 13292
rect 20115 13227 20181 13228
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 20299 12612 20365 12613
rect 20299 12548 20300 12612
rect 20364 12548 20365 12612
rect 20299 12547 20365 12548
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19379 9892 19445 9893
rect 19379 9828 19380 9892
rect 19444 9828 19445 9892
rect 19379 9827 19445 9828
rect 19568 9824 19888 10848
rect 20302 10709 20362 12547
rect 20486 10981 20546 25195
rect 22875 23764 22941 23765
rect 22875 23700 22876 23764
rect 22940 23700 22941 23764
rect 22875 23699 22941 23700
rect 22691 21996 22757 21997
rect 22691 21932 22692 21996
rect 22756 21932 22757 21996
rect 22691 21931 22757 21932
rect 21403 21452 21469 21453
rect 21403 21388 21404 21452
rect 21468 21388 21469 21452
rect 21403 21387 21469 21388
rect 21035 20364 21101 20365
rect 21035 20300 21036 20364
rect 21100 20300 21101 20364
rect 21035 20299 21101 20300
rect 20667 18052 20733 18053
rect 20667 17988 20668 18052
rect 20732 17988 20733 18052
rect 20667 17987 20733 17988
rect 20670 11661 20730 17987
rect 20851 14108 20917 14109
rect 20851 14044 20852 14108
rect 20916 14044 20917 14108
rect 20851 14043 20917 14044
rect 20667 11660 20733 11661
rect 20667 11596 20668 11660
rect 20732 11596 20733 11660
rect 20667 11595 20733 11596
rect 20483 10980 20549 10981
rect 20483 10916 20484 10980
rect 20548 10916 20549 10980
rect 20483 10915 20549 10916
rect 20299 10708 20365 10709
rect 20299 10644 20300 10708
rect 20364 10644 20365 10708
rect 20299 10643 20365 10644
rect 20854 9893 20914 14043
rect 20851 9892 20917 9893
rect 20851 9828 20852 9892
rect 20916 9828 20917 9892
rect 20851 9827 20917 9828
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 18643 9756 18709 9757
rect 18643 9692 18644 9756
rect 18708 9692 18709 9756
rect 18643 9691 18709 9692
rect 19568 8736 19888 9760
rect 21038 9485 21098 20299
rect 21035 9484 21101 9485
rect 21035 9420 21036 9484
rect 21100 9420 21101 9484
rect 21035 9419 21101 9420
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 17907 8396 17973 8397
rect 17907 8332 17908 8396
rect 17972 8332 17973 8396
rect 17907 8331 17973 8332
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 17171 4044 17237 4045
rect 17171 3980 17172 4044
rect 17236 3980 17237 4044
rect 17171 3979 17237 3980
rect 14411 3908 14477 3909
rect 14411 3844 14412 3908
rect 14476 3844 14477 3908
rect 14411 3843 14477 3844
rect 19568 3296 19888 4320
rect 21406 4045 21466 21387
rect 21955 20772 22021 20773
rect 21955 20708 21956 20772
rect 22020 20708 22021 20772
rect 21955 20707 22021 20708
rect 21771 15060 21837 15061
rect 21771 14996 21772 15060
rect 21836 14996 21837 15060
rect 21771 14995 21837 14996
rect 21403 4044 21469 4045
rect 21403 3980 21404 4044
rect 21468 3980 21469 4044
rect 21403 3979 21469 3980
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 5947 3228 6013 3229
rect 5947 3164 5948 3228
rect 6012 3164 6013 3228
rect 5947 3163 6013 3164
rect 4843 2548 4909 2549
rect 4843 2484 4844 2548
rect 4908 2484 4909 2548
rect 4843 2483 4909 2484
rect 19568 2208 19888 3232
rect 21406 3229 21466 3979
rect 21774 3773 21834 14995
rect 21958 6901 22018 20707
rect 22139 20500 22205 20501
rect 22139 20436 22140 20500
rect 22204 20436 22205 20500
rect 22139 20435 22205 20436
rect 22142 12885 22202 20435
rect 22507 13020 22573 13021
rect 22507 12956 22508 13020
rect 22572 12956 22573 13020
rect 22507 12955 22573 12956
rect 22139 12884 22205 12885
rect 22139 12820 22140 12884
rect 22204 12820 22205 12884
rect 22139 12819 22205 12820
rect 22139 12612 22205 12613
rect 22139 12548 22140 12612
rect 22204 12548 22205 12612
rect 22139 12547 22205 12548
rect 22142 9621 22202 12547
rect 22323 11524 22389 11525
rect 22323 11460 22324 11524
rect 22388 11460 22389 11524
rect 22323 11459 22389 11460
rect 22139 9620 22205 9621
rect 22139 9556 22140 9620
rect 22204 9556 22205 9620
rect 22139 9555 22205 9556
rect 22326 8261 22386 11459
rect 22323 8260 22389 8261
rect 22323 8196 22324 8260
rect 22388 8196 22389 8260
rect 22323 8195 22389 8196
rect 22510 7853 22570 12955
rect 22694 11797 22754 21931
rect 22878 13565 22938 23699
rect 23430 20773 23490 27643
rect 23611 23628 23677 23629
rect 23611 23564 23612 23628
rect 23676 23564 23677 23628
rect 23611 23563 23677 23564
rect 23427 20772 23493 20773
rect 23427 20708 23428 20772
rect 23492 20708 23493 20772
rect 23427 20707 23493 20708
rect 23059 15604 23125 15605
rect 23059 15540 23060 15604
rect 23124 15540 23125 15604
rect 23059 15539 23125 15540
rect 22875 13564 22941 13565
rect 22875 13500 22876 13564
rect 22940 13500 22941 13564
rect 22875 13499 22941 13500
rect 23062 13429 23122 15539
rect 23059 13428 23125 13429
rect 23059 13364 23060 13428
rect 23124 13364 23125 13428
rect 23059 13363 23125 13364
rect 22691 11796 22757 11797
rect 22691 11732 22692 11796
rect 22756 11732 22757 11796
rect 22691 11731 22757 11732
rect 23614 9485 23674 23563
rect 24166 16285 24226 32539
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 30051 23492 30117 23493
rect 30051 23428 30052 23492
rect 30116 23428 30117 23492
rect 30051 23427 30117 23428
rect 26923 22948 26989 22949
rect 26923 22884 26924 22948
rect 26988 22884 26989 22948
rect 26923 22883 26989 22884
rect 28211 22948 28277 22949
rect 28211 22884 28212 22948
rect 28276 22884 28277 22948
rect 28211 22883 28277 22884
rect 24715 20772 24781 20773
rect 24715 20708 24716 20772
rect 24780 20708 24781 20772
rect 24715 20707 24781 20708
rect 25267 20772 25333 20773
rect 25267 20708 25268 20772
rect 25332 20708 25333 20772
rect 25267 20707 25333 20708
rect 24163 16284 24229 16285
rect 24163 16220 24164 16284
rect 24228 16220 24229 16284
rect 24163 16219 24229 16220
rect 24531 15332 24597 15333
rect 24531 15268 24532 15332
rect 24596 15268 24597 15332
rect 24531 15267 24597 15268
rect 23611 9484 23677 9485
rect 23611 9420 23612 9484
rect 23676 9420 23677 9484
rect 23611 9419 23677 9420
rect 22507 7852 22573 7853
rect 22507 7788 22508 7852
rect 22572 7788 22573 7852
rect 22507 7787 22573 7788
rect 21955 6900 22021 6901
rect 21955 6836 21956 6900
rect 22020 6836 22021 6900
rect 21955 6835 22021 6836
rect 21771 3772 21837 3773
rect 21771 3708 21772 3772
rect 21836 3708 21837 3772
rect 21771 3707 21837 3708
rect 21403 3228 21469 3229
rect 21403 3164 21404 3228
rect 21468 3164 21469 3228
rect 21403 3163 21469 3164
rect 24534 2685 24594 15267
rect 24718 4045 24778 20707
rect 25083 18052 25149 18053
rect 25083 17988 25084 18052
rect 25148 17988 25149 18052
rect 25083 17987 25149 17988
rect 24899 12748 24965 12749
rect 24899 12684 24900 12748
rect 24964 12684 24965 12748
rect 24899 12683 24965 12684
rect 24902 8397 24962 12683
rect 25086 9213 25146 17987
rect 25270 12341 25330 20707
rect 25819 19140 25885 19141
rect 25819 19076 25820 19140
rect 25884 19076 25885 19140
rect 25819 19075 25885 19076
rect 25635 18188 25701 18189
rect 25635 18124 25636 18188
rect 25700 18124 25701 18188
rect 25635 18123 25701 18124
rect 25267 12340 25333 12341
rect 25267 12276 25268 12340
rect 25332 12276 25333 12340
rect 25267 12275 25333 12276
rect 25083 9212 25149 9213
rect 25083 9148 25084 9212
rect 25148 9148 25149 9212
rect 25083 9147 25149 9148
rect 24899 8396 24965 8397
rect 24899 8332 24900 8396
rect 24964 8332 24965 8396
rect 24899 8331 24965 8332
rect 25638 6901 25698 18123
rect 25822 10573 25882 19075
rect 26371 18188 26437 18189
rect 26371 18124 26372 18188
rect 26436 18124 26437 18188
rect 26371 18123 26437 18124
rect 26374 11117 26434 18123
rect 26555 18052 26621 18053
rect 26555 17988 26556 18052
rect 26620 17988 26621 18052
rect 26555 17987 26621 17988
rect 26558 12450 26618 17987
rect 26558 12390 26802 12450
rect 26555 11660 26621 11661
rect 26555 11596 26556 11660
rect 26620 11596 26621 11660
rect 26555 11595 26621 11596
rect 26371 11116 26437 11117
rect 26371 11052 26372 11116
rect 26436 11052 26437 11116
rect 26371 11051 26437 11052
rect 25819 10572 25885 10573
rect 25819 10508 25820 10572
rect 25884 10508 25885 10572
rect 25819 10507 25885 10508
rect 25635 6900 25701 6901
rect 25635 6836 25636 6900
rect 25700 6836 25701 6900
rect 25635 6835 25701 6836
rect 26558 4045 26618 11595
rect 26742 9893 26802 12390
rect 26739 9892 26805 9893
rect 26739 9828 26740 9892
rect 26804 9828 26805 9892
rect 26739 9827 26805 9828
rect 26926 9757 26986 22883
rect 27659 21452 27725 21453
rect 27659 21388 27660 21452
rect 27724 21388 27725 21452
rect 27659 21387 27725 21388
rect 27475 18324 27541 18325
rect 27475 18260 27476 18324
rect 27540 18260 27541 18324
rect 27475 18259 27541 18260
rect 27478 14381 27538 18259
rect 27475 14380 27541 14381
rect 27475 14316 27476 14380
rect 27540 14316 27541 14380
rect 27475 14315 27541 14316
rect 27478 12341 27538 14315
rect 27662 13701 27722 21387
rect 28214 20909 28274 22883
rect 28211 20908 28277 20909
rect 28211 20844 28212 20908
rect 28276 20844 28277 20908
rect 28211 20843 28277 20844
rect 27659 13700 27725 13701
rect 27659 13636 27660 13700
rect 27724 13636 27725 13700
rect 27659 13635 27725 13636
rect 27475 12340 27541 12341
rect 27475 12276 27476 12340
rect 27540 12276 27541 12340
rect 27475 12275 27541 12276
rect 26923 9756 26989 9757
rect 26923 9692 26924 9756
rect 26988 9692 26989 9756
rect 26923 9691 26989 9692
rect 27475 7716 27541 7717
rect 27475 7652 27476 7716
rect 27540 7652 27541 7716
rect 27475 7651 27541 7652
rect 27478 6493 27538 7651
rect 27475 6492 27541 6493
rect 27475 6428 27476 6492
rect 27540 6428 27541 6492
rect 27475 6427 27541 6428
rect 28214 5813 28274 20843
rect 29131 18732 29197 18733
rect 29131 18668 29132 18732
rect 29196 18668 29197 18732
rect 29131 18667 29197 18668
rect 28579 18596 28645 18597
rect 28579 18532 28580 18596
rect 28644 18532 28645 18596
rect 28579 18531 28645 18532
rect 28763 18596 28829 18597
rect 28763 18532 28764 18596
rect 28828 18532 28829 18596
rect 28763 18531 28829 18532
rect 28395 15740 28461 15741
rect 28395 15676 28396 15740
rect 28460 15676 28461 15740
rect 28395 15675 28461 15676
rect 28211 5812 28277 5813
rect 28211 5748 28212 5812
rect 28276 5748 28277 5812
rect 28211 5747 28277 5748
rect 28398 5541 28458 15675
rect 28582 12477 28642 18531
rect 28766 17373 28826 18531
rect 28947 18188 29013 18189
rect 28947 18124 28948 18188
rect 29012 18124 29013 18188
rect 28947 18123 29013 18124
rect 28950 17917 29010 18123
rect 28947 17916 29013 17917
rect 28947 17852 28948 17916
rect 29012 17852 29013 17916
rect 28947 17851 29013 17852
rect 28763 17372 28829 17373
rect 28763 17308 28764 17372
rect 28828 17308 28829 17372
rect 28763 17307 28829 17308
rect 28947 15332 29013 15333
rect 28947 15268 28948 15332
rect 29012 15268 29013 15332
rect 28947 15267 29013 15268
rect 28579 12476 28645 12477
rect 28579 12412 28580 12476
rect 28644 12412 28645 12476
rect 28579 12411 28645 12412
rect 28950 11661 29010 15267
rect 28947 11660 29013 11661
rect 28947 11596 28948 11660
rect 29012 11596 29013 11660
rect 28947 11595 29013 11596
rect 29134 10981 29194 18667
rect 29315 12340 29381 12341
rect 29315 12276 29316 12340
rect 29380 12276 29381 12340
rect 29315 12275 29381 12276
rect 29131 10980 29197 10981
rect 29131 10916 29132 10980
rect 29196 10916 29197 10980
rect 29131 10915 29197 10916
rect 28947 9892 29013 9893
rect 28947 9828 28948 9892
rect 29012 9828 29013 9892
rect 28947 9827 29013 9828
rect 28395 5540 28461 5541
rect 28395 5476 28396 5540
rect 28460 5476 28461 5540
rect 28395 5475 28461 5476
rect 28950 5133 29010 9827
rect 28947 5132 29013 5133
rect 28947 5068 28948 5132
rect 29012 5068 29013 5132
rect 28947 5067 29013 5068
rect 29318 4045 29378 12275
rect 30054 11797 30114 23427
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 31523 22540 31589 22541
rect 31523 22476 31524 22540
rect 31588 22476 31589 22540
rect 31523 22475 31589 22476
rect 30419 18188 30485 18189
rect 30419 18124 30420 18188
rect 30484 18124 30485 18188
rect 30419 18123 30485 18124
rect 30422 12450 30482 18123
rect 30787 13156 30853 13157
rect 30787 13092 30788 13156
rect 30852 13092 30853 13156
rect 30787 13091 30853 13092
rect 30422 12390 30666 12450
rect 30051 11796 30117 11797
rect 30051 11732 30052 11796
rect 30116 11732 30117 11796
rect 30051 11731 30117 11732
rect 30419 11660 30485 11661
rect 30419 11596 30420 11660
rect 30484 11596 30485 11660
rect 30419 11595 30485 11596
rect 30422 8533 30482 11595
rect 30606 9893 30666 12390
rect 30603 9892 30669 9893
rect 30603 9828 30604 9892
rect 30668 9828 30669 9892
rect 30603 9827 30669 9828
rect 30790 8941 30850 13091
rect 31526 12205 31586 22475
rect 34928 22336 35248 23360
rect 36859 23084 36925 23085
rect 36859 23020 36860 23084
rect 36924 23020 36925 23084
rect 36859 23019 36925 23020
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 32259 21860 32325 21861
rect 32259 21796 32260 21860
rect 32324 21796 32325 21860
rect 32259 21795 32325 21796
rect 31891 19412 31957 19413
rect 31891 19348 31892 19412
rect 31956 19348 31957 19412
rect 31891 19347 31957 19348
rect 32075 19412 32141 19413
rect 32075 19348 32076 19412
rect 32140 19348 32141 19412
rect 32075 19347 32141 19348
rect 31523 12204 31589 12205
rect 31523 12140 31524 12204
rect 31588 12140 31589 12204
rect 31523 12139 31589 12140
rect 31523 11660 31589 11661
rect 31523 11596 31524 11660
rect 31588 11596 31589 11660
rect 31523 11595 31589 11596
rect 30787 8940 30853 8941
rect 30787 8876 30788 8940
rect 30852 8876 30853 8940
rect 30787 8875 30853 8876
rect 30419 8532 30485 8533
rect 30419 8468 30420 8532
rect 30484 8468 30485 8532
rect 30419 8467 30485 8468
rect 30787 8532 30853 8533
rect 30787 8468 30788 8532
rect 30852 8468 30853 8532
rect 30787 8467 30853 8468
rect 30419 7988 30485 7989
rect 30419 7924 30420 7988
rect 30484 7924 30485 7988
rect 30419 7923 30485 7924
rect 30422 6901 30482 7923
rect 30419 6900 30485 6901
rect 30419 6836 30420 6900
rect 30484 6836 30485 6900
rect 30419 6835 30485 6836
rect 30790 6629 30850 8467
rect 31526 7037 31586 11595
rect 31523 7036 31589 7037
rect 31523 6972 31524 7036
rect 31588 6972 31589 7036
rect 31523 6971 31589 6972
rect 30787 6628 30853 6629
rect 30787 6564 30788 6628
rect 30852 6564 30853 6628
rect 30787 6563 30853 6564
rect 24715 4044 24781 4045
rect 24715 3980 24716 4044
rect 24780 3980 24781 4044
rect 24715 3979 24781 3980
rect 26555 4044 26621 4045
rect 26555 3980 26556 4044
rect 26620 3980 26621 4044
rect 26555 3979 26621 3980
rect 29315 4044 29381 4045
rect 29315 3980 29316 4044
rect 29380 3980 29381 4044
rect 29315 3979 29381 3980
rect 26558 3229 26618 3979
rect 26555 3228 26621 3229
rect 26555 3164 26556 3228
rect 26620 3164 26621 3228
rect 26555 3163 26621 3164
rect 31894 2790 31954 19347
rect 32078 15741 32138 19347
rect 32075 15740 32141 15741
rect 32075 15676 32076 15740
rect 32140 15676 32141 15740
rect 32075 15675 32141 15676
rect 32262 12613 32322 21795
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 32443 19820 32509 19821
rect 32443 19756 32444 19820
rect 32508 19756 32509 19820
rect 32443 19755 32509 19756
rect 32259 12612 32325 12613
rect 32259 12548 32260 12612
rect 32324 12548 32325 12612
rect 32259 12547 32325 12548
rect 32446 12477 32506 19755
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 32627 17372 32693 17373
rect 32627 17308 32628 17372
rect 32692 17308 32693 17372
rect 32627 17307 32693 17308
rect 32443 12476 32509 12477
rect 32443 12412 32444 12476
rect 32508 12412 32509 12476
rect 32443 12411 32509 12412
rect 32075 8940 32141 8941
rect 32075 8876 32076 8940
rect 32140 8876 32141 8940
rect 32075 8875 32141 8876
rect 32078 7717 32138 8875
rect 32075 7716 32141 7717
rect 32075 7652 32076 7716
rect 32140 7652 32141 7716
rect 32075 7651 32141 7652
rect 32630 3773 32690 17307
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 33179 16692 33245 16693
rect 33179 16628 33180 16692
rect 33244 16628 33245 16692
rect 33179 16627 33245 16628
rect 33182 14653 33242 16627
rect 33731 16556 33797 16557
rect 33731 16492 33732 16556
rect 33796 16492 33797 16556
rect 33731 16491 33797 16492
rect 33179 14652 33245 14653
rect 33179 14588 33180 14652
rect 33244 14588 33245 14652
rect 33179 14587 33245 14588
rect 33734 5541 33794 16491
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 35755 12884 35821 12885
rect 35755 12820 35756 12884
rect 35820 12820 35821 12884
rect 35755 12819 35821 12820
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 33731 5540 33797 5541
rect 33731 5476 33732 5540
rect 33796 5476 33797 5540
rect 33731 5475 33797 5476
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 35758 4045 35818 12819
rect 36123 11116 36189 11117
rect 36123 11052 36124 11116
rect 36188 11052 36189 11116
rect 36123 11051 36189 11052
rect 35755 4044 35821 4045
rect 35755 3980 35756 4044
rect 35820 3980 35821 4044
rect 35755 3979 35821 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 32627 3772 32693 3773
rect 32627 3708 32628 3772
rect 32692 3708 32693 3772
rect 32627 3707 32693 3708
rect 31710 2730 31954 2790
rect 34928 2752 35248 3776
rect 24531 2684 24597 2685
rect 24531 2620 24532 2684
rect 24596 2620 24597 2684
rect 24531 2619 24597 2620
rect 31710 2549 31770 2730
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 31707 2548 31773 2549
rect 31707 2484 31708 2548
rect 31772 2484 31773 2548
rect 31707 2483 31773 2484
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 36126 2413 36186 11051
rect 36862 5541 36922 23019
rect 36859 5540 36925 5541
rect 36859 5476 36860 5540
rect 36924 5476 36925 5540
rect 36859 5475 36925 5476
rect 36123 2412 36189 2413
rect 36123 2348 36124 2412
rect 36188 2348 36189 2412
rect 36123 2347 36189 2348
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 33488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 34132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 33488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1667941163
transform 1 0 35512 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1667941163
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1667941163
transform 1 0 17388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1667941163
transform 1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1667941163
transform 1 0 27600 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1667941163
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1667941163
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1667941163
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1667941163
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1667941163
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1667941163
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1667941163
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1667941163
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1667941163
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1667941163
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_196
timestamp 1667941163
transform 1 0 19136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1667941163
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1667941163
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1667941163
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1667941163
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1667941163
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_376
timestamp 1667941163
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_100
timestamp 1667941163
transform 1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1667941163
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1667941163
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1667941163
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_259
timestamp 1667941163
transform 1 0 24932 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_267
timestamp 1667941163
transform 1 0 25668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_291
timestamp 1667941163
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1667941163
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1667941163
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_318
timestamp 1667941163
transform 1 0 30360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_343
timestamp 1667941163
transform 1 0 32660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1667941163
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_380
timestamp 1667941163
transform 1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1667941163
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1667941163
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1667941163
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1667941163
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_153
timestamp 1667941163
transform 1 0 15180 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1667941163
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_180
timestamp 1667941163
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1667941163
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1667941163
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_240
timestamp 1667941163
transform 1 0 23184 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_246
timestamp 1667941163
transform 1 0 23736 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_270
timestamp 1667941163
transform 1 0 25944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1667941163
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_306
timestamp 1667941163
transform 1 0 29256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1667941163
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_357
timestamp 1667941163
transform 1 0 33948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_376
timestamp 1667941163
transform 1 0 35696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_380
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1667941163
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1667941163
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1667941163
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_100
timestamp 1667941163
transform 1 0 10304 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1667941163
transform 1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1667941163
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1667941163
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_214
timestamp 1667941163
transform 1 0 20792 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1667941163
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_266
timestamp 1667941163
transform 1 0 25576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_293
timestamp 1667941163
transform 1 0 28060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1667941163
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1667941163
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_355
timestamp 1667941163
transform 1 0 33764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1667941163
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_385
timestamp 1667941163
transform 1 0 36524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_391
timestamp 1667941163
transform 1 0 37076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_17
timestamp 1667941163
transform 1 0 2668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1667941163
transform 1 0 3220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1667941163
transform 1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 1667941163
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1667941163
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1667941163
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1667941163
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1667941163
transform 1 0 13800 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1667941163
transform 1 0 19228 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_247
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_251
timestamp 1667941163
transform 1 0 24196 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1667941163
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_306
timestamp 1667941163
transform 1 0 29256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_330
timestamp 1667941163
transform 1 0 31464 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_350
timestamp 1667941163
transform 1 0 33304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_354
timestamp 1667941163
transform 1 0 33672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_369
timestamp 1667941163
transform 1 0 35052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_376
timestamp 1667941163
transform 1 0 35696 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_384
timestamp 1667941163
transform 1 0 36432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1667941163
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_17
timestamp 1667941163
transform 1 0 2668 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1667941163
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_37
timestamp 1667941163
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1667941163
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1667941163
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_167
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1667941163
transform 1 0 19596 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1667941163
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1667941163
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_257
timestamp 1667941163
transform 1 0 24748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_268
timestamp 1667941163
transform 1 0 25760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1667941163
transform 1 0 28244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1667941163
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1667941163
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_348
timestamp 1667941163
transform 1 0 33120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1667941163
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1667941163
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_384
timestamp 1667941163
transform 1 0 36432 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_392
timestamp 1667941163
transform 1 0 37168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1667941163
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1667941163
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1667941163
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1667941163
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1667941163
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1667941163
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1667941163
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1667941163
transform 1 0 14996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1667941163
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_212
timestamp 1667941163
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1667941163
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1667941163
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_271
timestamp 1667941163
transform 1 0 26036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_303
timestamp 1667941163
transform 1 0 28980 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_327
timestamp 1667941163
transform 1 0 31188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1667941163
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_350
timestamp 1667941163
transform 1 0 33304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_354
timestamp 1667941163
transform 1 0 33672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_369
timestamp 1667941163
transform 1 0 35052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_376
timestamp 1667941163
transform 1 0 35696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_383
timestamp 1667941163
transform 1 0 36340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1667941163
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1667941163
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp 1667941163
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1667941163
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1667941163
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1667941163
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1667941163
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_89
timestamp 1667941163
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_104
timestamp 1667941163
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1667941163
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1667941163
transform 1 0 15272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1667941163
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_187
timestamp 1667941163
transform 1 0 18308 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_203
timestamp 1667941163
transform 1 0 19780 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_211
timestamp 1667941163
transform 1 0 20516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_236
timestamp 1667941163
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_296
timestamp 1667941163
transform 1 0 28336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1667941163
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1667941163
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_348
timestamp 1667941163
transform 1 0 33120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_355
timestamp 1667941163
transform 1 0 33764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1667941163
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_370
timestamp 1667941163
transform 1 0 35144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_384
timestamp 1667941163
transform 1 0 36432 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_391
timestamp 1667941163
transform 1 0 37076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_399
timestamp 1667941163
transform 1 0 37812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1667941163
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1667941163
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1667941163
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1667941163
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1667941163
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1667941163
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1667941163
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1667941163
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1667941163
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1667941163
transform 1 0 14444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1667941163
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1667941163
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_204
timestamp 1667941163
transform 1 0 19872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1667941163
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1667941163
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_247
timestamp 1667941163
transform 1 0 23828 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_271
timestamp 1667941163
transform 1 0 26036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_303
timestamp 1667941163
transform 1 0 28980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_327
timestamp 1667941163
transform 1 0 31188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1667941163
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_348
timestamp 1667941163
transform 1 0 33120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_355
timestamp 1667941163
transform 1 0 33764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_362
timestamp 1667941163
transform 1 0 34408 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_369
timestamp 1667941163
transform 1 0 35052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_376
timestamp 1667941163
transform 1 0 35696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_383
timestamp 1667941163
transform 1 0 36340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1667941163
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_398
timestamp 1667941163
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_9
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_19
timestamp 1667941163
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1667941163
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_111
timestamp 1667941163
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_146
timestamp 1667941163
transform 1 0 14536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1667941163
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_222
timestamp 1667941163
transform 1 0 21528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_226
timestamp 1667941163
transform 1 0 21896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1667941163
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_269
timestamp 1667941163
transform 1 0 25852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_296
timestamp 1667941163
transform 1 0 28336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1667941163
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_322
timestamp 1667941163
transform 1 0 30728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_341
timestamp 1667941163
transform 1 0 32476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_348
timestamp 1667941163
transform 1 0 33120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_355
timestamp 1667941163
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1667941163
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_370
timestamp 1667941163
transform 1 0 35144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_384
timestamp 1667941163
transform 1 0 36432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_391
timestamp 1667941163
transform 1 0 37076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_399
timestamp 1667941163
transform 1 0 37812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1667941163
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_17
timestamp 1667941163
transform 1 0 2668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1667941163
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_38
timestamp 1667941163
transform 1 0 4600 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_44
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1667941163
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1667941163
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1667941163
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1667941163
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_247
timestamp 1667941163
transform 1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_271
timestamp 1667941163
transform 1 0 26036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_303
timestamp 1667941163
transform 1 0 28980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp 1667941163
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_311
timestamp 1667941163
transform 1 0 29716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1667941163
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_342
timestamp 1667941163
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_356
timestamp 1667941163
transform 1 0 33856 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_363
timestamp 1667941163
transform 1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_370
timestamp 1667941163
transform 1 0 35144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_377
timestamp 1667941163
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1667941163
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1667941163
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1667941163
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1667941163
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1667941163
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1667941163
transform 1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1667941163
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1667941163
transform 1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1667941163
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1667941163
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1667941163
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1667941163
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1667941163
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_266
timestamp 1667941163
transform 1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_293
timestamp 1667941163
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1667941163
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1667941163
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_352
timestamp 1667941163
transform 1 0 33488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1667941163
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_370
timestamp 1667941163
transform 1 0 35144 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_379
timestamp 1667941163
transform 1 0 35972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_386
timestamp 1667941163
transform 1 0 36616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_393
timestamp 1667941163
transform 1 0 37260 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_8
timestamp 1667941163
transform 1 0 1840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1667941163
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_26
timestamp 1667941163
transform 1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1667941163
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1667941163
transform 1 0 4784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_47
timestamp 1667941163
transform 1 0 5428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_138
timestamp 1667941163
transform 1 0 13800 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1667941163
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_188
timestamp 1667941163
transform 1 0 18400 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_247
timestamp 1667941163
transform 1 0 23828 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_255
timestamp 1667941163
transform 1 0 24564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1667941163
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_303
timestamp 1667941163
transform 1 0 28980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_310
timestamp 1667941163
transform 1 0 29624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_314
timestamp 1667941163
transform 1 0 29992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_328
timestamp 1667941163
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_342
timestamp 1667941163
transform 1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_356
timestamp 1667941163
transform 1 0 33856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_363
timestamp 1667941163
transform 1 0 34500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_370
timestamp 1667941163
transform 1 0 35144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_374
timestamp 1667941163
transform 1 0 35512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_378
timestamp 1667941163
transform 1 0 35880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_398
timestamp 1667941163
transform 1 0 37720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1667941163
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1667941163
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_37
timestamp 1667941163
transform 1 0 4508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1667941163
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1667941163
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1667941163
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_166
timestamp 1667941163
transform 1 0 16376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_205
timestamp 1667941163
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1667941163
transform 1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1667941163
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1667941163
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1667941163
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_334
timestamp 1667941163
transform 1 0 31832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_341
timestamp 1667941163
transform 1 0 32476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_348
timestamp 1667941163
transform 1 0 33120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_355
timestamp 1667941163
transform 1 0 33764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1667941163
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1667941163
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_385
timestamp 1667941163
transform 1 0 36524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_390
timestamp 1667941163
transform 1 0 36984 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_397
timestamp 1667941163
transform 1 0 37628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1667941163
transform 1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_29
timestamp 1667941163
transform 1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1667941163
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1667941163
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_63
timestamp 1667941163
transform 1 0 6900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1667941163
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 1667941163
transform 1 0 9384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1667941163
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_122
timestamp 1667941163
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1667941163
transform 1 0 14536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1667941163
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_200
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_212
timestamp 1667941163
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1667941163
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1667941163
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_320
timestamp 1667941163
transform 1 0 30544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_327
timestamp 1667941163
transform 1 0 31188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1667941163
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_345
timestamp 1667941163
transform 1 0 32844 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_352
timestamp 1667941163
transform 1 0 33488 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_364
timestamp 1667941163
transform 1 0 34592 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_372
timestamp 1667941163
transform 1 0 35328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1667941163
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_383
timestamp 1667941163
transform 1 0 36340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1667941163
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_16
timestamp 1667941163
transform 1 0 2576 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_22
timestamp 1667941163
transform 1 0 3128 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_34
timestamp 1667941163
transform 1 0 4232 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_42
timestamp 1667941163
transform 1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1667941163
transform 1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_54
timestamp 1667941163
transform 1 0 6072 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1667941163
transform 1 0 6624 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1667941163
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1667941163
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114
timestamp 1667941163
transform 1 0 11592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1667941163
transform 1 0 14536 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1667941163
transform 1 0 15088 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_174
timestamp 1667941163
transform 1 0 17112 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1667941163
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_222
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_296
timestamp 1667941163
transform 1 0 28336 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_328
timestamp 1667941163
transform 1 0 31280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_335
timestamp 1667941163
transform 1 0 31924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_354
timestamp 1667941163
transform 1 0 33672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1667941163
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_384
timestamp 1667941163
transform 1 0 36432 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_392
timestamp 1667941163
transform 1 0 37168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1667941163
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1667941163
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_16
timestamp 1667941163
transform 1 0 2576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_28
timestamp 1667941163
transform 1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_34
timestamp 1667941163
transform 1 0 4232 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_42
timestamp 1667941163
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_66
timestamp 1667941163
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1667941163
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp 1667941163
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1667941163
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1667941163
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_210
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_263
timestamp 1667941163
transform 1 0 25300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1667941163
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1667941163
transform 1 0 29256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_314
timestamp 1667941163
transform 1 0 29992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_319
timestamp 1667941163
transform 1 0 30452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_326
timestamp 1667941163
transform 1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1667941163
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_344
timestamp 1667941163
transform 1 0 32752 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_356
timestamp 1667941163
transform 1 0 33856 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_368
timestamp 1667941163
transform 1 0 34960 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_383
timestamp 1667941163
transform 1 0 36340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_398
timestamp 1667941163
transform 1 0 37720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_45
timestamp 1667941163
transform 1 0 5244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_57
timestamp 1667941163
transform 1 0 6348 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_66
timestamp 1667941163
transform 1 0 7176 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1667941163
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_96
timestamp 1667941163
transform 1 0 9936 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1667941163
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_114
timestamp 1667941163
transform 1 0 11592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_230
timestamp 1667941163
transform 1 0 22264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1667941163
transform 1 0 23000 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1667941163
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_290
timestamp 1667941163
transform 1 0 27784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_335
timestamp 1667941163
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_347
timestamp 1667941163
transform 1 0 33028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_355
timestamp 1667941163
transform 1 0 33764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1667941163
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_370
timestamp 1667941163
transform 1 0 35144 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_382
timestamp 1667941163
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_394
timestamp 1667941163
transform 1 0 37352 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_405
timestamp 1667941163
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_32
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_40
timestamp 1667941163
transform 1 0 4784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_44
timestamp 1667941163
transform 1 0 5152 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_50
timestamp 1667941163
transform 1 0 5704 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1667941163
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 1667941163
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1667941163
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1667941163
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_122
timestamp 1667941163
transform 1 0 12328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1667941163
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 1667941163
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_201
timestamp 1667941163
transform 1 0 19596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_250
timestamp 1667941163
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1667941163
transform 1 0 24748 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_264
timestamp 1667941163
transform 1 0 25392 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1667941163
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_321
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1667941163
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_368
timestamp 1667941163
transform 1 0 34960 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_380
timestamp 1667941163
transform 1 0 36064 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_9
timestamp 1667941163
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1667941163
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_37
timestamp 1667941163
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_49
timestamp 1667941163
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1667941163
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_90
timestamp 1667941163
transform 1 0 9384 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1667941163
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_106
timestamp 1667941163
transform 1 0 10856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1667941163
transform 1 0 11592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1667941163
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1667941163
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_216
timestamp 1667941163
transform 1 0 20976 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1667941163
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1667941163
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_280
timestamp 1667941163
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_295
timestamp 1667941163
transform 1 0 28244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_351
timestamp 1667941163
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_64
timestamp 1667941163
transform 1 0 6992 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1667941163
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1667941163
transform 1 0 8280 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1667941163
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_102
timestamp 1667941163
transform 1 0 10488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_106
timestamp 1667941163
transform 1 0 10856 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_124
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_153
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1667941163
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_248
timestamp 1667941163
transform 1 0 23920 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_256
timestamp 1667941163
transform 1 0 24656 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_306
timestamp 1667941163
transform 1 0 29256 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_312
timestamp 1667941163
transform 1 0 29808 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1667941163
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_323
timestamp 1667941163
transform 1 0 30820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_13
timestamp 1667941163
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1667941163
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_60
timestamp 1667941163
transform 1 0 6624 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_68
timestamp 1667941163
transform 1 0 7360 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1667941163
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1667941163
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1667941163
transform 1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1667941163
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1667941163
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_170
timestamp 1667941163
transform 1 0 16744 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_242
timestamp 1667941163
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1667941163
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_264
timestamp 1667941163
transform 1 0 25392 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1667941163
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_295
timestamp 1667941163
transform 1 0 28244 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1667941163
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_313
timestamp 1667941163
transform 1 0 29900 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_323
timestamp 1667941163
transform 1 0 30820 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_330
timestamp 1667941163
transform 1 0 31464 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_342
timestamp 1667941163
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_354
timestamp 1667941163
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1667941163
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_393
timestamp 1667941163
transform 1 0 37260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_397
timestamp 1667941163
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_70
timestamp 1667941163
transform 1 0 7544 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_89
timestamp 1667941163
transform 1 0 9292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_95
timestamp 1667941163
transform 1 0 9844 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1667941163
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1667941163
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_148
timestamp 1667941163
transform 1 0 14720 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1667941163
transform 1 0 17480 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_185
timestamp 1667941163
transform 1 0 18124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_202
timestamp 1667941163
transform 1 0 19688 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_208
timestamp 1667941163
transform 1 0 20240 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1667941163
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1667941163
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_241
timestamp 1667941163
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1667941163
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_258
timestamp 1667941163
transform 1 0 24840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1667941163
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_300
timestamp 1667941163
transform 1 0 28704 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_307
timestamp 1667941163
transform 1 0 29348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_314
timestamp 1667941163
transform 1 0 29992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_318
timestamp 1667941163
transform 1 0 30360 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_328
timestamp 1667941163
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_342
timestamp 1667941163
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_354
timestamp 1667941163
transform 1 0 33672 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_366
timestamp 1667941163
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_378
timestamp 1667941163
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1667941163
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_402
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1667941163
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1667941163
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1667941163
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1667941163
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_60
timestamp 1667941163
transform 1 0 6624 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1667941163
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1667941163
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_105
timestamp 1667941163
transform 1 0 10764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_113
timestamp 1667941163
transform 1 0 11500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1667941163
transform 1 0 11868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1667941163
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_173
timestamp 1667941163
transform 1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1667941163
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1667941163
transform 1 0 18308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1667941163
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_211
timestamp 1667941163
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 1667941163
transform 1 0 23276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1667941163
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_261
timestamp 1667941163
transform 1 0 25116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_268
timestamp 1667941163
transform 1 0 25760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_275
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_282
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1667941163
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_328
timestamp 1667941163
transform 1 0 31280 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_335
timestamp 1667941163
transform 1 0 31924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_347
timestamp 1667941163
transform 1 0 33028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_73
timestamp 1667941163
transform 1 0 7820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_90
timestamp 1667941163
transform 1 0 9384 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_128
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_141
timestamp 1667941163
transform 1 0 14076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_155
timestamp 1667941163
transform 1 0 15364 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1667941163
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_190
timestamp 1667941163
transform 1 0 18584 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_204
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_211
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_252
timestamp 1667941163
transform 1 0 24288 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_259
timestamp 1667941163
transform 1 0 24932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_266
timestamp 1667941163
transform 1 0 25576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_313
timestamp 1667941163
transform 1 0 29900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_320
timestamp 1667941163
transform 1 0 30544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_327
timestamp 1667941163
transform 1 0 31188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1667941163
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_352
timestamp 1667941163
transform 1 0 33488 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_364
timestamp 1667941163
transform 1 0 34592 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_376
timestamp 1667941163
transform 1 0 35696 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1667941163
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_10
timestamp 1667941163
transform 1 0 2024 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1667941163
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1667941163
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_49
timestamp 1667941163
transform 1 0 5612 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_56
timestamp 1667941163
transform 1 0 6256 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1667941163
transform 1 0 6900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1667941163
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_100
timestamp 1667941163
transform 1 0 10304 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_106
timestamp 1667941163
transform 1 0 10856 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_110
timestamp 1667941163
transform 1 0 11224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1667941163
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1667941163
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1667941163
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1667941163
transform 1 0 14536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_166
timestamp 1667941163
transform 1 0 16376 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_172
timestamp 1667941163
transform 1 0 16928 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_176
timestamp 1667941163
transform 1 0 17296 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_218
timestamp 1667941163
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_235
timestamp 1667941163
transform 1 0 22724 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_258
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_272
timestamp 1667941163
transform 1 0 26128 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1667941163
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_314
timestamp 1667941163
transform 1 0 29992 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_322
timestamp 1667941163
transform 1 0 30728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_336
timestamp 1667941163
transform 1 0 32016 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1667941163
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1667941163
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_370
timestamp 1667941163
transform 1 0 35144 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_382
timestamp 1667941163
transform 1 0 36248 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_394
timestamp 1667941163
transform 1 0 37352 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1667941163
transform 1 0 38456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp 1667941163
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1667941163
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1667941163
transform 1 0 9200 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1667941163
transform 1 0 9568 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1667941163
transform 1 0 9936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1667941163
transform 1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_128
timestamp 1667941163
transform 1 0 12880 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_198
timestamp 1667941163
transform 1 0 19320 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_212
timestamp 1667941163
transform 1 0 20608 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_242
timestamp 1667941163
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1667941163
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1667941163
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_289
timestamp 1667941163
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1667941163
transform 1 0 29624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_327
timestamp 1667941163
transform 1 0 31188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1667941163
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_342
timestamp 1667941163
transform 1 0 32568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_356
timestamp 1667941163
transform 1 0 33856 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_368
timestamp 1667941163
transform 1 0 34960 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_380
timestamp 1667941163
transform 1 0 36064 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_401
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_57
timestamp 1667941163
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1667941163
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1667941163
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_96
timestamp 1667941163
transform 1 0 9936 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_104
timestamp 1667941163
transform 1 0 10672 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_108
timestamp 1667941163
transform 1 0 11040 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_115
timestamp 1667941163
transform 1 0 11684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1667941163
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_155
timestamp 1667941163
transform 1 0 15364 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1667941163
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1667941163
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_183
timestamp 1667941163
transform 1 0 17940 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_210
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_223
timestamp 1667941163
transform 1 0 21620 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1667941163
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1667941163
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_268
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_276
timestamp 1667941163
transform 1 0 26496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_287
timestamp 1667941163
transform 1 0 27508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1667941163
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_326
timestamp 1667941163
transform 1 0 31096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_339
timestamp 1667941163
transform 1 0 32292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_346
timestamp 1667941163
transform 1 0 32936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_353
timestamp 1667941163
transform 1 0 33580 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1667941163
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_370
timestamp 1667941163
transform 1 0 35144 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1667941163
transform 1 0 7728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_79
timestamp 1667941163
transform 1 0 8372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_85
timestamp 1667941163
transform 1 0 8924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1667941163
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1667941163
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1667941163
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1667941163
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_134
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_146
timestamp 1667941163
transform 1 0 14536 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_154
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1667941163
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1667941163
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1667941163
transform 1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_216
timestamp 1667941163
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp 1667941163
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_233
timestamp 1667941163
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_240
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_259
timestamp 1667941163
transform 1 0 24932 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_267
timestamp 1667941163
transform 1 0 25668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_292
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1667941163
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1667941163
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1667941163
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_355
timestamp 1667941163
transform 1 0 33764 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1667941163
transform 1 0 34408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_369
timestamp 1667941163
transform 1 0 35052 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_376
timestamp 1667941163
transform 1 0 35696 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1667941163
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_62
timestamp 1667941163
transform 1 0 6808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_74
timestamp 1667941163
transform 1 0 7912 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1667941163
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1667941163
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_127
timestamp 1667941163
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1667941163
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_164
timestamp 1667941163
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_175
timestamp 1667941163
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_187
timestamp 1667941163
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1667941163
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1667941163
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_215
timestamp 1667941163
transform 1 0 20884 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1667941163
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1667941163
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_258
timestamp 1667941163
transform 1 0 24840 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_266
timestamp 1667941163
transform 1 0 25576 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1667941163
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1667941163
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1667941163
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_320
timestamp 1667941163
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_341
timestamp 1667941163
transform 1 0 32476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1667941163
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_370
timestamp 1667941163
transform 1 0 35144 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_382
timestamp 1667941163
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_394
timestamp 1667941163
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1667941163
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1667941163
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_72
timestamp 1667941163
transform 1 0 7728 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_78
timestamp 1667941163
transform 1 0 8280 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1667941163
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1667941163
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_129
timestamp 1667941163
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_133
timestamp 1667941163
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_140
timestamp 1667941163
transform 1 0 13984 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_151
timestamp 1667941163
transform 1 0 14996 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_155
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1667941163
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1667941163
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_239
timestamp 1667941163
transform 1 0 23092 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_256
timestamp 1667941163
transform 1 0 24656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1667941163
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_303
timestamp 1667941163
transform 1 0 28980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_322
timestamp 1667941163
transform 1 0 30728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_330
timestamp 1667941163
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_342
timestamp 1667941163
transform 1 0 32568 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_359
timestamp 1667941163
transform 1 0 34132 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_366
timestamp 1667941163
transform 1 0 34776 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_381
timestamp 1667941163
transform 1 0 36156 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_401
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_122
timestamp 1667941163
transform 1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1667941163
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1667941163
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1667941163
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_232
timestamp 1667941163
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1667941163
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_268
timestamp 1667941163
transform 1 0 25760 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1667941163
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_279
timestamp 1667941163
transform 1 0 26772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1667941163
transform 1 0 28336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_303
timestamp 1667941163
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_320
timestamp 1667941163
transform 1 0 30544 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_335
timestamp 1667941163
transform 1 0 31924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_342
timestamp 1667941163
transform 1 0 32568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_349
timestamp 1667941163
transform 1 0 33212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1667941163
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_370
timestamp 1667941163
transform 1 0 35144 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_382
timestamp 1667941163
transform 1 0 36248 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_394
timestamp 1667941163
transform 1 0 37352 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_400
timestamp 1667941163
transform 1 0 37904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_10
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_22
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_34
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1667941163
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_65
timestamp 1667941163
transform 1 0 7084 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_77
timestamp 1667941163
transform 1 0 8188 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_89
timestamp 1667941163
transform 1 0 9292 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_101
timestamp 1667941163
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1667941163
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1667941163
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1667941163
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_132
timestamp 1667941163
transform 1 0 13248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1667941163
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_156
timestamp 1667941163
transform 1 0 15456 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_162
timestamp 1667941163
transform 1 0 16008 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_184
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_190
timestamp 1667941163
transform 1 0 18584 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_204
timestamp 1667941163
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1667941163
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1667941163
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_240
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_268
timestamp 1667941163
transform 1 0 25760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1667941163
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_296
timestamp 1667941163
transform 1 0 28336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_313
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_319
timestamp 1667941163
transform 1 0 30452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1667941163
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1667941163
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_355
timestamp 1667941163
transform 1 0 33764 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_362
timestamp 1667941163
transform 1 0 34408 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_369
timestamp 1667941163
transform 1 0 35052 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_381
timestamp 1667941163
transform 1 0 36156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1667941163
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1667941163
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1667941163
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_122
timestamp 1667941163
transform 1 0 12328 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1667941163
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1667941163
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1667941163
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1667941163
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_216
timestamp 1667941163
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_220
timestamp 1667941163
transform 1 0 21344 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1667941163
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_241
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_258
timestamp 1667941163
transform 1 0 24840 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_264
timestamp 1667941163
transform 1 0 25392 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_286
timestamp 1667941163
transform 1 0 27416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_290
timestamp 1667941163
transform 1 0 27784 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1667941163
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_327
timestamp 1667941163
transform 1 0 31188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1667941163
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_349
timestamp 1667941163
transform 1 0 33212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_356
timestamp 1667941163
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_99
timestamp 1667941163
transform 1 0 10212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_118
timestamp 1667941163
transform 1 0 11960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1667941163
transform 1 0 13248 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_145
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_157
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1667941163
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_186
timestamp 1667941163
transform 1 0 18216 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_190
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_197
timestamp 1667941163
transform 1 0 19228 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1667941163
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1667941163
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1667941163
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1667941163
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1667941163
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1667941163
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_312
timestamp 1667941163
transform 1 0 29808 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_320
timestamp 1667941163
transform 1 0 30544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1667941163
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_342
timestamp 1667941163
transform 1 0 32568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_356
timestamp 1667941163
transform 1 0 33856 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_363
timestamp 1667941163
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_375
timestamp 1667941163
transform 1 0 35604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1667941163
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1667941163
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_71
timestamp 1667941163
transform 1 0 7636 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1667941163
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1667941163
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_127
timestamp 1667941163
transform 1 0 12788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_147
timestamp 1667941163
transform 1 0 14628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_173
timestamp 1667941163
transform 1 0 17020 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_179
timestamp 1667941163
transform 1 0 17572 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1667941163
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_218
timestamp 1667941163
transform 1 0 21160 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1667941163
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_237
timestamp 1667941163
transform 1 0 22908 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1667941163
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_259
timestamp 1667941163
transform 1 0 24932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_273
timestamp 1667941163
transform 1 0 26220 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1667941163
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1667941163
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_314
timestamp 1667941163
transform 1 0 29992 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_335
timestamp 1667941163
transform 1 0 31924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_342
timestamp 1667941163
transform 1 0 32568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_346
timestamp 1667941163
transform 1 0 32936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_350
timestamp 1667941163
transform 1 0 33304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_371
timestamp 1667941163
transform 1 0 35236 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_383
timestamp 1667941163
transform 1 0 36340 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_395
timestamp 1667941163
transform 1 0 37444 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_91
timestamp 1667941163
transform 1 0 9476 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_120
timestamp 1667941163
transform 1 0 12144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_127
timestamp 1667941163
transform 1 0 12788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_144
timestamp 1667941163
transform 1 0 14352 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_150
timestamp 1667941163
transform 1 0 14904 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1667941163
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_178
timestamp 1667941163
transform 1 0 17480 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_186
timestamp 1667941163
transform 1 0 18216 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_190
timestamp 1667941163
transform 1 0 18584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_198
timestamp 1667941163
transform 1 0 19320 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_210
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_229
timestamp 1667941163
transform 1 0 22172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_243
timestamp 1667941163
transform 1 0 23460 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1667941163
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_269
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1667941163
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1667941163
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_309
timestamp 1667941163
transform 1 0 29532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_313
timestamp 1667941163
transform 1 0 29900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_327
timestamp 1667941163
transform 1 0 31188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1667941163
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_342
timestamp 1667941163
transform 1 0 32568 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_370
timestamp 1667941163
transform 1 0 35144 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_382
timestamp 1667941163
transform 1 0 36248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1667941163
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_69
timestamp 1667941163
transform 1 0 7452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1667941163
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_90
timestamp 1667941163
transform 1 0 9384 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_102
timestamp 1667941163
transform 1 0 10488 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1667941163
transform 1 0 10856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_113
timestamp 1667941163
transform 1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1667941163
transform 1 0 13064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_134
timestamp 1667941163
transform 1 0 13432 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_152
timestamp 1667941163
transform 1 0 15088 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_158
timestamp 1667941163
transform 1 0 15640 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1667941163
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_202
timestamp 1667941163
transform 1 0 19688 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_214
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1667941163
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1667941163
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_268
timestamp 1667941163
transform 1 0 25760 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_275
timestamp 1667941163
transform 1 0 26404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_281
timestamp 1667941163
transform 1 0 26956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_285
timestamp 1667941163
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_292
timestamp 1667941163
transform 1 0 27968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_299
timestamp 1667941163
transform 1 0 28612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1667941163
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_324
timestamp 1667941163
transform 1 0 30912 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_331
timestamp 1667941163
transform 1 0 31556 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_348
timestamp 1667941163
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1667941163
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_372
timestamp 1667941163
transform 1 0 35328 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_384
timestamp 1667941163
transform 1 0 36432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_396
timestamp 1667941163
transform 1 0 37536 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_404
timestamp 1667941163
transform 1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_10
timestamp 1667941163
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_17
timestamp 1667941163
transform 1 0 2668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1667941163
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 1667941163
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1667941163
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_99
timestamp 1667941163
transform 1 0 10212 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_119
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_127
timestamp 1667941163
transform 1 0 12788 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_135
timestamp 1667941163
transform 1 0 13524 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1667941163
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_201
timestamp 1667941163
transform 1 0 19596 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1667941163
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1667941163
transform 1 0 23184 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1667941163
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1667941163
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_268
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_274
timestamp 1667941163
transform 1 0 26312 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_296
timestamp 1667941163
transform 1 0 28336 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_313
timestamp 1667941163
transform 1 0 29900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_320
timestamp 1667941163
transform 1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_327
timestamp 1667941163
transform 1 0 31188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1667941163
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_344
timestamp 1667941163
transform 1 0 32752 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_352
timestamp 1667941163
transform 1 0 33488 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_357
timestamp 1667941163
transform 1 0 33948 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_369
timestamp 1667941163
transform 1 0 35052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_381
timestamp 1667941163
transform 1 0 36156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1667941163
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_402
timestamp 1667941163
transform 1 0 38088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1667941163
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1667941163
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1667941163
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1667941163
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1667941163
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_93
timestamp 1667941163
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_110
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_116
timestamp 1667941163
transform 1 0 11776 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1667941163
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1667941163
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_146
timestamp 1667941163
transform 1 0 14536 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_156
timestamp 1667941163
transform 1 0 15456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_206
timestamp 1667941163
transform 1 0 20056 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_214
timestamp 1667941163
transform 1 0 20792 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_229
timestamp 1667941163
transform 1 0 22172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_258
timestamp 1667941163
transform 1 0 24840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1667941163
transform 1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_279
timestamp 1667941163
transform 1 0 26772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_285
timestamp 1667941163
transform 1 0 27324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_326
timestamp 1667941163
transform 1 0 31096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_334
timestamp 1667941163
transform 1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_349
timestamp 1667941163
transform 1 0 33212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1667941163
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1667941163
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_102
timestamp 1667941163
transform 1 0 10488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_106
timestamp 1667941163
transform 1 0 10856 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_122
timestamp 1667941163
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_129
timestamp 1667941163
transform 1 0 12972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_136
timestamp 1667941163
transform 1 0 13616 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_144
timestamp 1667941163
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_156
timestamp 1667941163
transform 1 0 15456 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_162
timestamp 1667941163
transform 1 0 16008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_184
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1667941163
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_195
timestamp 1667941163
transform 1 0 19044 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_199
timestamp 1667941163
transform 1 0 19412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_231
timestamp 1667941163
transform 1 0 22356 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_245
timestamp 1667941163
transform 1 0 23644 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1667941163
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_269
timestamp 1667941163
transform 1 0 25852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1667941163
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_304
timestamp 1667941163
transform 1 0 29072 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_311
timestamp 1667941163
transform 1 0 29716 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_324
timestamp 1667941163
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_345
timestamp 1667941163
transform 1 0 32844 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_9
timestamp 1667941163
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1667941163
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_94
timestamp 1667941163
transform 1 0 9752 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1667941163
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_108
timestamp 1667941163
transform 1 0 11040 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_120
timestamp 1667941163
transform 1 0 12144 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_128
timestamp 1667941163
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_156
timestamp 1667941163
transform 1 0 15456 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_162
timestamp 1667941163
transform 1 0 16008 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_166
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_183
timestamp 1667941163
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_215
timestamp 1667941163
transform 1 0 20884 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_228
timestamp 1667941163
transform 1 0 22080 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1667941163
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1667941163
transform 1 0 24932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_276
timestamp 1667941163
transform 1 0 26496 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_293
timestamp 1667941163
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1667941163
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_324
timestamp 1667941163
transform 1 0 30912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_328
timestamp 1667941163
transform 1 0 31280 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_342
timestamp 1667941163
transform 1 0 32568 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_350
timestamp 1667941163
transform 1 0 33304 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_98
timestamp 1667941163
transform 1 0 10120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_129
timestamp 1667941163
transform 1 0 12972 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_133
timestamp 1667941163
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1667941163
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1667941163
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_174
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_189
timestamp 1667941163
transform 1 0 18492 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_204
timestamp 1667941163
transform 1 0 19872 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_216
timestamp 1667941163
transform 1 0 20976 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_231
timestamp 1667941163
transform 1 0 22356 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_250
timestamp 1667941163
transform 1 0 24104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_263
timestamp 1667941163
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_270
timestamp 1667941163
transform 1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1667941163
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_297
timestamp 1667941163
transform 1 0 28428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1667941163
transform 1 0 28796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_318
timestamp 1667941163
transform 1 0 30360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_325
timestamp 1667941163
transform 1 0 31004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1667941163
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_357
timestamp 1667941163
transform 1 0 33948 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_362
timestamp 1667941163
transform 1 0 34408 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_374
timestamp 1667941163
transform 1 0 35512 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1667941163
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_100
timestamp 1667941163
transform 1 0 10304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1667941163
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_151
timestamp 1667941163
transform 1 0 14996 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_159
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_169
timestamp 1667941163
transform 1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_173
timestamp 1667941163
transform 1 0 17020 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_187
timestamp 1667941163
transform 1 0 18308 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_212
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_231
timestamp 1667941163
transform 1 0 22356 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1667941163
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_264
timestamp 1667941163
transform 1 0 25392 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_285
timestamp 1667941163
transform 1 0 27324 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_292
timestamp 1667941163
transform 1 0 27968 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_299
timestamp 1667941163
transform 1 0 28612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_324
timestamp 1667941163
transform 1 0 30912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_331
timestamp 1667941163
transform 1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_338
timestamp 1667941163
transform 1 0 32200 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_8
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1667941163
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1667941163
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_96
timestamp 1667941163
transform 1 0 9936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_123
timestamp 1667941163
transform 1 0 12420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_140
timestamp 1667941163
transform 1 0 13984 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1667941163
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_186
timestamp 1667941163
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_199
timestamp 1667941163
transform 1 0 19412 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_207
timestamp 1667941163
transform 1 0 20148 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1667941163
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_230
timestamp 1667941163
transform 1 0 22264 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_247
timestamp 1667941163
transform 1 0 23828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_253
timestamp 1667941163
transform 1 0 24380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1667941163
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1667941163
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_287
timestamp 1667941163
transform 1 0 27508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_291
timestamp 1667941163
transform 1 0 27876 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_312
timestamp 1667941163
transform 1 0 29808 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_324
timestamp 1667941163
transform 1 0 30912 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_344
timestamp 1667941163
transform 1 0 32752 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_352
timestamp 1667941163
transform 1 0 33488 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_364
timestamp 1667941163
transform 1 0 34592 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_376
timestamp 1667941163
transform 1 0 35696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1667941163
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_401
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1667941163
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1667941163
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1667941163
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_100
timestamp 1667941163
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_113
timestamp 1667941163
transform 1 0 11500 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1667941163
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1667941163
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_156
timestamp 1667941163
transform 1 0 15456 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_169
timestamp 1667941163
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1667941163
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_215
timestamp 1667941163
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_223
timestamp 1667941163
transform 1 0 21620 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_240
timestamp 1667941163
transform 1 0 23184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1667941163
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_268
timestamp 1667941163
transform 1 0 25760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1667941163
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1667941163
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_314
timestamp 1667941163
transform 1 0 29992 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_63
timestamp 1667941163
transform 1 0 6900 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_70
timestamp 1667941163
transform 1 0 7544 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_88
timestamp 1667941163
transform 1 0 9200 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_100
timestamp 1667941163
transform 1 0 10304 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1667941163
transform 1 0 12328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_129
timestamp 1667941163
transform 1 0 12972 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_141
timestamp 1667941163
transform 1 0 14076 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_153
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_174
timestamp 1667941163
transform 1 0 17112 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_200
timestamp 1667941163
transform 1 0 19504 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_206
timestamp 1667941163
transform 1 0 20056 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_210
timestamp 1667941163
transform 1 0 20424 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_218
timestamp 1667941163
transform 1 0 21160 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_231
timestamp 1667941163
transform 1 0 22356 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1667941163
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_269
timestamp 1667941163
transform 1 0 25852 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1667941163
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_286
timestamp 1667941163
transform 1 0 27416 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_310
timestamp 1667941163
transform 1 0 29624 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_323
timestamp 1667941163
transform 1 0 30820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_49
timestamp 1667941163
transform 1 0 5612 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_60
timestamp 1667941163
transform 1 0 6624 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_66
timestamp 1667941163
transform 1 0 7176 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_70
timestamp 1667941163
transform 1 0 7544 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1667941163
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_124
timestamp 1667941163
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_131
timestamp 1667941163
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1667941163
transform 1 0 14536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_166
timestamp 1667941163
transform 1 0 16376 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_173
timestamp 1667941163
transform 1 0 17020 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_185
timestamp 1667941163
transform 1 0 18124 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1667941163
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_212
timestamp 1667941163
transform 1 0 20608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_216
timestamp 1667941163
transform 1 0 20976 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1667941163
transform 1 0 22264 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1667941163
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_258
timestamp 1667941163
transform 1 0 24840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_282
timestamp 1667941163
transform 1 0 27048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_294
timestamp 1667941163
transform 1 0 28152 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_298
timestamp 1667941163
transform 1 0 28520 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_302
timestamp 1667941163
transform 1 0 28888 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1667941163
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_317
timestamp 1667941163
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_323
timestamp 1667941163
transform 1 0 30820 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_335
timestamp 1667941163
transform 1 0 31924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_347
timestamp 1667941163
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1667941163
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1667941163
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_87
timestamp 1667941163
transform 1 0 9108 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_91
timestamp 1667941163
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_103
timestamp 1667941163
transform 1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_132
timestamp 1667941163
transform 1 0 13248 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_145
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_157
timestamp 1667941163
transform 1 0 15548 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_213
timestamp 1667941163
transform 1 0 20700 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1667941163
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_230
timestamp 1667941163
transform 1 0 22264 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_236
timestamp 1667941163
transform 1 0 22816 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1667941163
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_257
timestamp 1667941163
transform 1 0 24748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_265
timestamp 1667941163
transform 1 0 25484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1667941163
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_286
timestamp 1667941163
transform 1 0 27416 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_298
timestamp 1667941163
transform 1 0 28520 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_310
timestamp 1667941163
transform 1 0 29624 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_322
timestamp 1667941163
transform 1 0 30728 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1667941163
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1667941163
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_59
timestamp 1667941163
transform 1 0 6532 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_63
timestamp 1667941163
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_75
timestamp 1667941163
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_95
timestamp 1667941163
transform 1 0 9844 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_106
timestamp 1667941163
transform 1 0 10856 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_118
timestamp 1667941163
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_130
timestamp 1667941163
transform 1 0 13064 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1667941163
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_150
timestamp 1667941163
transform 1 0 14904 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_157
timestamp 1667941163
transform 1 0 15548 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_164
timestamp 1667941163
transform 1 0 16192 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1667941163
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_176
timestamp 1667941163
transform 1 0 17296 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_187
timestamp 1667941163
transform 1 0 18308 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1667941163
transform 1 0 22080 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_236
timestamp 1667941163
transform 1 0 22816 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_241
timestamp 1667941163
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1667941163
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_274
timestamp 1667941163
transform 1 0 26312 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_281
timestamp 1667941163
transform 1 0 26956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_293
timestamp 1667941163
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1667941163
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_122
timestamp 1667941163
transform 1 0 12328 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_133
timestamp 1667941163
transform 1 0 13340 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_140
timestamp 1667941163
transform 1 0 13984 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_157
timestamp 1667941163
transform 1 0 15548 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_180
timestamp 1667941163
transform 1 0 17664 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_192
timestamp 1667941163
transform 1 0 18768 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_204
timestamp 1667941163
transform 1 0 19872 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1667941163
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_240
timestamp 1667941163
transform 1 0 23184 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_247
timestamp 1667941163
transform 1 0 23828 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_254
timestamp 1667941163
transform 1 0 24472 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_264
timestamp 1667941163
transform 1 0 25392 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_272
timestamp 1667941163
transform 1 0 26128 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_301
timestamp 1667941163
transform 1 0 28796 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_312
timestamp 1667941163
transform 1 0 29808 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_324
timestamp 1667941163
transform 1 0 30912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1667941163
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_33
timestamp 1667941163
transform 1 0 4140 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_37
timestamp 1667941163
transform 1 0 4508 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_49
timestamp 1667941163
transform 1 0 5612 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_61
timestamp 1667941163
transform 1 0 6716 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_73
timestamp 1667941163
transform 1 0 7820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1667941163
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_105
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_119
timestamp 1667941163
transform 1 0 12052 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_127
timestamp 1667941163
transform 1 0 12788 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1667941163
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_157
timestamp 1667941163
transform 1 0 15548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_169
timestamp 1667941163
transform 1 0 16652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_181
timestamp 1667941163
transform 1 0 17756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1667941163
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1667941163
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1667941163
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_258
timestamp 1667941163
transform 1 0 24840 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_270
timestamp 1667941163
transform 1 0 25944 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_282
timestamp 1667941163
transform 1 0 27048 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_294
timestamp 1667941163
transform 1 0 28152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1667941163
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_73
timestamp 1667941163
transform 1 0 7820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_85
timestamp 1667941163
transform 1 0 8924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_97
timestamp 1667941163
transform 1 0 10028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_109
timestamp 1667941163
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_153
timestamp 1667941163
transform 1 0 15180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1667941163
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_175
timestamp 1667941163
transform 1 0 17204 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_187
timestamp 1667941163
transform 1 0 18308 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_199
timestamp 1667941163
transform 1 0 19412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1667941163
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_268
timestamp 1667941163
transform 1 0 25760 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_398
timestamp 1667941163
transform 1 0 37720 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1667941163
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_49
timestamp 1667941163
transform 1 0 5612 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_90
timestamp 1667941163
transform 1 0 9384 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_102
timestamp 1667941163
transform 1 0 10488 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_114
timestamp 1667941163
transform 1 0 11592 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_122
timestamp 1667941163
transform 1 0 12328 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_127
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1667941163
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_210
timestamp 1667941163
transform 1 0 20424 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1667941163
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_324
timestamp 1667941163
transform 1 0 30912 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_202
timestamp 1667941163
transform 1 0 19688 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_214
timestamp 1667941163
transform 1 0 20792 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_226
timestamp 1667941163
transform 1 0 21896 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_238
timestamp 1667941163
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_274
timestamp 1667941163
transform 1 0 26312 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_286
timestamp 1667941163
transform 1 0 27416 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1667941163
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1667941163
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1667941163
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1667941163
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_45
timestamp 1667941163
transform 1 0 5244 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_286
timestamp 1667941163
transform 1 0 27416 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_290
timestamp 1667941163
transform 1 0 27784 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_302
timestamp 1667941163
transform 1 0 28888 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_314
timestamp 1667941163
transform 1 0 29992 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_326
timestamp 1667941163
transform 1 0 31096 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1667941163
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_380
timestamp 1667941163
transform 1 0 36064 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1667941163
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_20
timestamp 1667941163
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_32
timestamp 1667941163
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_44
timestamp 1667941163
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_395
timestamp 1667941163
transform 1 0 37444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_399
timestamp 1667941163
transform 1 0 37812 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_16
timestamp 1667941163
transform 1 0 2576 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_28
timestamp 1667941163
transform 1 0 3680 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_40
timestamp 1667941163
transform 1 0 4784 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1667941163
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_230
timestamp 1667941163
transform 1 0 22264 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_238
timestamp 1667941163
transform 1 0 23000 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_244
timestamp 1667941163
transform 1 0 23552 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_256
timestamp 1667941163
transform 1 0 24656 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_268
timestamp 1667941163
transform 1 0 25760 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_17
timestamp 1667941163
transform 1 0 2668 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1667941163
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_69
timestamp 1667941163
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1667941163
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_17
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_25
timestamp 1667941163
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_37
timestamp 1667941163
transform 1 0 4508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 1667941163
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_61
timestamp 1667941163
transform 1 0 6716 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_65
timestamp 1667941163
transform 1 0 7084 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_73
timestamp 1667941163
transform 1 0 7820 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_77
timestamp 1667941163
transform 1 0 8188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_85
timestamp 1667941163
transform 1 0 8924 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_90
timestamp 1667941163
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1667941163
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_119
timestamp 1667941163
transform 1 0 12052 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_131
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_153
timestamp 1667941163
transform 1 0 15180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1667941163
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_174
timestamp 1667941163
transform 1 0 17112 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_186
timestamp 1667941163
transform 1 0 18216 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_192
timestamp 1667941163
transform 1 0 18768 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_196
timestamp 1667941163
transform 1 0 19136 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1667941163
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_207
timestamp 1667941163
transform 1 0 20148 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_211
timestamp 1667941163
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_231
timestamp 1667941163
transform 1 0 22356 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_235
timestamp 1667941163
transform 1 0 22724 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_241
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1667941163
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_252
timestamp 1667941163
transform 1 0 24288 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_264
timestamp 1667941163
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1667941163
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_343
timestamp 1667941163
transform 1 0 32660 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_355
timestamp 1667941163
transform 1 0 33764 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_367
timestamp 1667941163
transform 1 0 34868 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_372
timestamp 1667941163
transform 1 0 35328 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_376
timestamp 1667941163
transform 1 0 35696 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_382
timestamp 1667941163
transform 1 0 36248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_96
timestamp 1667941163
transform 1 0 9936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_155
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_186
timestamp 1667941163
transform 1 0 18216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_217
timestamp 1667941163
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1667941163
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1667941163
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_246
timestamp 1667941163
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_275
timestamp 1667941163
transform 1 0 26404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_302
timestamp 1667941163
transform 1 0 28888 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_349
timestamp 1667941163
transform 1 0 33212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_387
timestamp 1667941163
transform 1 0 36708 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0493_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 16744 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 16100 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 15272 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 10304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 12052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 28520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 28428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 16100 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 32936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 27048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 36156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 19596 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 19688 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 20976 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 12144 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 12512 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 9200 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 10948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 14352 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 14628 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 12972 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 16100 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 9844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 26128 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 7820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 26128 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 20884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 28336 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 31648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 29532 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 30912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 26128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 36064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 31464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 30360 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 32936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 34776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 32936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 32476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 34500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 22632 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 28704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 22264 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 7360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 17112 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 6716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 3220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 33304 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 32292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 32936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 29532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 33488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 26772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 32936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 32292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 23276 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 6716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 17204 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 11316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 25208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 27784 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 28980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 25208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 19136 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 20148 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 34776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 21528 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 12052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 11224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 25484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 36064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 6808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 36708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 26312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 33488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 32292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 29900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 34132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 32292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 22908 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 31280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 31556 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 22632 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 13156 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 17296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 25208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 25208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 17480 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 21804 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 28980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 28980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 24196 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 32292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 31556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 32292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 18124 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 15088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 14536 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 30544 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 33580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 33580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 6164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 14444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 8004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 17204 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 31004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 32660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 20148 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 19504 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 15916 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 20884 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 18952 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 12052 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 20240 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 31280 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 28336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 13616 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 19228 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 26036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 16652 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 36064 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 18308 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 25576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 23276 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 27416 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 12696 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 34132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 24656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 18400 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 12328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 33212 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 30912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 34132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 6624 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 13432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 5336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 25576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 36156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 36156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 31556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 25208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 19780 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 30912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 32292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 31556 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 15180 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 37352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0799_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 6624 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 5704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 33672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 23276 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0807_
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 5704 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 30636 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 7268 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 26036 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 35052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 13156 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 26312 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 7360 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 32476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 32292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 34776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 33488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 28244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 37444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 17020 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 34132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 36708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 8280 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 7268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 4508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 33580 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 23552 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 12880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0852_
timestamp 1667941163
transform 1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 31924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 34040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 25668 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 28520 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 27140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 10580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1667941163
transform 1 0 23000 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 7544 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 32568 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 26496 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 32936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 37444 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 25484 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1667941163
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1667941163
transform 1 0 35696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1667941163
transform 1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1667941163
transform 1 0 34224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1667941163
transform 1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1667941163
transform 1 0 7176 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1667941163
transform 1 0 34132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1667941163
transform 1 0 25576 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1667941163
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1667941163
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1667941163
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1667941163
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1667941163
transform 1 0 10580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1667941163
transform 1 0 33580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1667941163
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1667941163
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1667941163
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1667941163
transform 1 0 8924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1667941163
transform 1 0 26312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1667941163
transform 1 0 11776 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1667941163
transform 1 0 33028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1667941163
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1667941163
transform 1 0 8280 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1667941163
transform 1 0 12512 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0909_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0910_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0911_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20976 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1667941163
transform 1 0 37444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1667941163
transform 1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1667941163
transform 1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1667941163
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1667941163
transform 1 0 31556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1667941163
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1667941163
transform 1 0 34224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1667941163
transform 1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1667941163
transform 1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0922_
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1667941163
transform 1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1667941163
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1667941163
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1667941163
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1667941163
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1667941163
transform 1 0 34132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1667941163
transform 1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1667941163
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0933_
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1667941163
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1667941163
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1667941163
transform 1 0 16744 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1667941163
transform 1 0 13432 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1667941163
transform 1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1667941163
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1667941163
transform 1 0 24564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1667941163
transform 1 0 23736 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0944_
timestamp 1667941163
transform 1 0 21804 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1667941163
transform 1 0 29072 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1667941163
transform 1 0 28612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1667941163
transform 1 0 14260 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0955_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21620 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1667941163
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1667941163
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1667941163
transform 1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1667941163
transform 1 0 32568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0966_
timestamp 1667941163
transform 1 0 23644 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1667941163
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1667941163
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1667941163
transform 1 0 17848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1667941163
transform 1 0 15824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1667941163
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1667941163
transform 1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1667941163
transform 1 0 17204 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1667941163
transform 1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0977_
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1667941163
transform 1 0 18032 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1667941163
transform 1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1667941163
transform 1 0 29624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1667941163
transform 1 0 27784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1667941163
transform 1 0 28428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1667941163
transform 1 0 27968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1667941163
transform 1 0 26128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1667941163
transform 1 0 30728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1667941163
transform 1 0 36800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1667941163
transform 1 0 33580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1667941163
transform 1 0 20976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1667941163
transform 1 0 14720 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1667941163
transform 1 0 35512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0999_
timestamp 1667941163
transform 1 0 25944 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1667941163
transform 1 0 36064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1667941163
transform 1 0 36156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1667941163
transform 1 0 35512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1667941163
transform 1 0 20332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1667941163
transform 1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1667941163
transform 1 0 34132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1667941163
transform 1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1010_
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1667941163
transform 1 0 20056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1667941163
transform 1 0 33580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1667941163
transform 1 0 30176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1667941163
transform 1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1667941163
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1021_
timestamp 1667941163
transform 1 0 28704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1667941163
transform 1 0 33488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1667941163
transform 1 0 35512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1667941163
transform 1 0 31648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1667941163
transform 1 0 33488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1667941163
transform 1 0 30544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1667941163
transform 1 0 37352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1032_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1667941163
transform 1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1667941163
transform 1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1667941163
transform 1 0 32936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1667941163
transform 1 0 33856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1667941163
transform 1 0 35512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1667941163
transform 1 0 29716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1667941163
transform 1 0 24472 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1667941163
transform 1 0 31188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1043_
timestamp 1667941163
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1667941163
transform 1 0 13064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1667941163
transform 1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1667941163
transform 1 0 12972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1667941163
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1667941163
transform 1 0 29348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1667941163
transform 1 0 30360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1667941163
transform 1 0 36156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1667941163
transform 1 0 15824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1054_
timestamp 1667941163
transform 1 0 22724 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1667941163
transform 1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1667941163
transform 1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1667941163
transform 1 0 12880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1065_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1667941163
transform 1 0 36800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1667941163
transform 1 0 36708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1667941163
transform 1 0 19412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1667941163
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1667941163
transform 1 0 19044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1078_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1079_
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 1667941163
transform 1 0 29716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 1667941163
transform 1 0 24196 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1082_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1083_
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1084_
timestamp 1667941163
transform 1 0 25760 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1085_
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1086_
timestamp 1667941163
transform 1 0 4600 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 1667941163
transform 1 0 7084 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1089_
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1090_
timestamp 1667941163
transform 1 0 11776 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1091_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1092_
timestamp 1667941163
transform 1 0 11040 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1093_
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1667941163
transform 1 0 29624 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1667941163
transform 1 0 14168 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1098_
timestamp 1667941163
transform 1 0 11684 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1099_
timestamp 1667941163
transform 1 0 16836 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1100_
timestamp 1667941163
transform 1 0 18032 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1101_
timestamp 1667941163
transform 1 0 11224 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1667941163
transform 1 0 9384 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1667941163
transform 1 0 12328 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1667941163
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1106_
timestamp 1667941163
transform 1 0 17388 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1107_
timestamp 1667941163
transform 1 0 20148 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1108_
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1109_
timestamp 1667941163
transform 1 0 25944 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1667941163
transform 1 0 9384 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1114_
timestamp 1667941163
transform 1 0 12236 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1115_
timestamp 1667941163
transform 1 0 19044 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1116_
timestamp 1667941163
transform 1 0 13064 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1117_
timestamp 1667941163
transform 1 0 16468 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1667941163
transform 1 0 6716 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1667941163
transform 1 0 4232 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1667941163
transform 1 0 4600 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1667941163
transform 1 0 6808 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1122_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1123_
timestamp 1667941163
transform 1 0 13064 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1124_
timestamp 1667941163
transform 1 0 11040 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1125_
timestamp 1667941163
transform 1 0 15456 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1667941163
transform 1 0 24196 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1667941163
transform 1 0 27140 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1130_
timestamp 1667941163
transform 1 0 18308 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1131_
timestamp 1667941163
transform 1 0 12236 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1132_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1133_
timestamp 1667941163
transform 1 0 18952 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1667941163
transform 1 0 14628 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1667941163
transform 1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1667941163
transform 1 0 9476 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1138_
timestamp 1667941163
transform 1 0 10948 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1139_
timestamp 1667941163
transform 1 0 20792 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1141_
timestamp 1667941163
transform 1 0 25944 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1667941163
transform 1 0 23460 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1143_
timestamp 1667941163
transform 1 0 22080 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1667941163
transform 1 0 22264 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1146_
timestamp 1667941163
transform 1 0 20792 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1147_
timestamp 1667941163
transform 1 0 25668 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1148_
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1149_
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1154_
timestamp 1667941163
transform 1 0 14260 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1155_
timestamp 1667941163
transform 1 0 16836 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1156_
timestamp 1667941163
transform 1 0 16836 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1157_
timestamp 1667941163
transform 1 0 20424 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1667941163
transform 1 0 24196 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1162_
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1163_
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1164_
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1165_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1667941163
transform 1 0 14628 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1667941163
transform 1 0 17112 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1667941163
transform 1 0 14536 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1170_
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1171_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1172_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1173_
timestamp 1667941163
transform 1 0 26220 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1667941163
transform 1 0 24840 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1178_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1179_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1180_
timestamp 1667941163
transform 1 0 19412 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1181_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1667941163
transform 1 0 21988 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1667941163
transform 1 0 14904 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1186_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1187_
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1188_
timestamp 1667941163
transform 1 0 14536 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1189_
timestamp 1667941163
transform 1 0 20700 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1667941163
transform 1 0 29624 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1667941163
transform 1 0 29348 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1667941163
transform 1 0 29348 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1194_
timestamp 1667941163
transform 1 0 26220 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1195_
timestamp 1667941163
transform 1 0 24748 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1196_
timestamp 1667941163
transform 1 0 24196 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1197_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1667941163
transform 1 0 7176 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1667941163
transform 1 0 9476 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1667941163
transform 1 0 6808 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1667941163
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1202_
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1203_
timestamp 1667941163
transform 1 0 24288 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1204_
timestamp 1667941163
transform 1 0 20884 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1205_
timestamp 1667941163
transform 1 0 26128 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1667941163
transform 1 0 9752 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1667941163
transform 1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1209_
timestamp 1667941163
transform 1 0 11684 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1210_
timestamp 1667941163
transform 1 0 12420 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1211_
timestamp 1667941163
transform 1 0 12420 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1667941163
transform 1 0 24196 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1667941163
transform 1 0 14536 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1215_
timestamp 1667941163
transform 1 0 16836 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1216_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1217_
timestamp 1667941163
transform 1 0 11684 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1221_
timestamp 1667941163
transform 1 0 18492 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1222_
timestamp 1667941163
transform 1 0 16744 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1223_
timestamp 1667941163
transform 1 0 11684 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1224_
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1667941163
transform 1 0 11960 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1226_
timestamp 1667941163
transform 1 0 12328 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1227_
timestamp 1667941163
transform 1 0 11684 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1228_
timestamp 1667941163
transform 1 0 16192 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1229_
timestamp 1667941163
transform 1 0 12328 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_2  _1250_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1251_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1667941163
transform 1 0 19504 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1254_
timestamp 1667941163
transform 1 0 37812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1255_
timestamp 1667941163
transform 1 0 12420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1667941163
transform 1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1667941163
transform 1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1667941163
transform 1 0 7912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1667941163
transform 1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1260_
timestamp 1667941163
transform 1 0 36248 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1667941163
transform 1 0 23368 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1667941163
transform 1 0 2300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1667941163
transform 1 0 20240 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1667941163
transform 1 0 38088 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1667941163
transform 1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1267_
timestamp 1667941163
transform 1 0 36248 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1268_
timestamp 1667941163
transform 1 0 35788 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1269_
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1667941163
transform 1 0 6808 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1272_
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1667941163
transform 1 0 11868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1274_
timestamp 1667941163
transform 1 0 33672 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1667941163
transform 1 0 6624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1276_
timestamp 1667941163
transform 1 0 32476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1667941163
transform 1 0 37812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1667941163
transform 1 0 35512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1280_
timestamp 1667941163
transform 1 0 20148 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1281_
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1282_
timestamp 1667941163
transform 1 0 33120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1667941163
transform 1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1285_
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1286_
timestamp 1667941163
transform 1 0 25024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1288_
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1289_
timestamp 1667941163
transform 1 0 33120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1290_
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1291_
timestamp 1667941163
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1667941163
transform 1 0 31556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1293_
timestamp 1667941163
transform 1 0 27784 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1667941163
transform 1 0 3772 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1667941163
transform 1 0 22448 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1667941163
transform 1 0 21988 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1297_
timestamp 1667941163
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1667941163
transform 1 0 36340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1667941163
transform 1 0 37352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1300_
timestamp 1667941163
transform 1 0 12972 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1667941163
transform 1 0 35052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1667941163
transform 1 0 38088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1303_
timestamp 1667941163
transform 1 0 27140 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1667941163
transform 1 0 18032 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1306_
timestamp 1667941163
transform 1 0 37168 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1667941163
transform 1 0 22632 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1308_
timestamp 1667941163
transform 1 0 31096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1309_
timestamp 1667941163
transform 1 0 4232 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1310_
timestamp 1667941163
transform 1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1667941163
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1667941163
transform 1 0 6348 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1314_
timestamp 1667941163
transform 1 0 9108 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1315_
timestamp 1667941163
transform 1 0 34960 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1316_
timestamp 1667941163
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1667941163
transform 1 0 34684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1318_
timestamp 1667941163
transform 1 0 16836 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1320_
timestamp 1667941163
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 1667941163
transform 1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1322_
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1667941163
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1324_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1667941163
transform 1 0 35604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1326_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29348 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1327_
timestamp 1667941163
transform 1 0 29808 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1328__172 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1328_
timestamp 1667941163
transform 1 0 31924 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1329_
timestamp 1667941163
transform 1 0 30084 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1330_
timestamp 1667941163
transform 1 0 20148 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1331_
timestamp 1667941163
transform 1 0 18400 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1332_
timestamp 1667941163
transform 1 0 25668 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1333_
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1334_
timestamp 1667941163
transform 1 0 12052 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1335_
timestamp 1667941163
transform 1 0 29992 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1336_
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1337_
timestamp 1667941163
transform 1 0 33856 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1338_
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1339_
timestamp 1667941163
transform 1 0 27140 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1340_
timestamp 1667941163
transform 1 0 30728 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1341_
timestamp 1667941163
transform 1 0 33028 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1342_
timestamp 1667941163
transform 1 0 7452 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1343_
timestamp 1667941163
transform 1 0 7820 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1344_
timestamp 1667941163
transform 1 0 7820 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1344__173
timestamp 1667941163
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1345_
timestamp 1667941163
transform 1 0 14168 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1346_
timestamp 1667941163
transform 1 0 7360 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1347_
timestamp 1667941163
transform 1 0 7268 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1348_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5796 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1349_
timestamp 1667941163
transform 1 0 6624 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1350_
timestamp 1667941163
transform 1 0 6716 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1351_
timestamp 1667941163
transform 1 0 6992 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1352_
timestamp 1667941163
transform 1 0 6624 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1353_
timestamp 1667941163
transform 1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1354_
timestamp 1667941163
transform 1 0 4876 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1355_
timestamp 1667941163
transform 1 0 5428 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1356_
timestamp 1667941163
transform 1 0 7360 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1357_
timestamp 1667941163
transform 1 0 5244 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1358_
timestamp 1667941163
transform 1 0 30728 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1359_
timestamp 1667941163
transform 1 0 22172 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1360_
timestamp 1667941163
transform 1 0 32476 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1360__174
timestamp 1667941163
transform 1 0 32568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1361_
timestamp 1667941163
transform 1 0 11592 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1362_
timestamp 1667941163
transform 1 0 10028 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1363_
timestamp 1667941163
transform 1 0 16744 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1364_
timestamp 1667941163
transform 1 0 30820 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1365_
timestamp 1667941163
transform 1 0 30544 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1366_
timestamp 1667941163
transform 1 0 28428 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1367_
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1368_
timestamp 1667941163
transform 1 0 14904 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1369_
timestamp 1667941163
transform 1 0 28060 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1370_
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1371_
timestamp 1667941163
transform 1 0 15824 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1372_
timestamp 1667941163
transform 1 0 21252 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1373_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1374_
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1375_
timestamp 1667941163
transform 1 0 18676 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1376__175
timestamp 1667941163
transform 1 0 12696 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1376_
timestamp 1667941163
transform 1 0 12604 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1377_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1378_
timestamp 1667941163
transform 1 0 18584 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1379_
timestamp 1667941163
transform 1 0 18124 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1380_
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1381_
timestamp 1667941163
transform 1 0 18676 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1382_
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1383_
timestamp 1667941163
transform 1 0 26128 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1384_
timestamp 1667941163
transform 1 0 29716 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1385_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1386_
timestamp 1667941163
transform 1 0 19780 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1387_
timestamp 1667941163
transform 1 0 24472 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1388_
timestamp 1667941163
transform 1 0 34500 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1389_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1390_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1391_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1392__176
timestamp 1667941163
transform 1 0 19412 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1392_
timestamp 1667941163
transform 1 0 19228 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1393_
timestamp 1667941163
transform 1 0 21068 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1394_
timestamp 1667941163
transform 1 0 20976 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1395_
timestamp 1667941163
transform 1 0 14996 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1396_
timestamp 1667941163
transform 1 0 22632 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1397_
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1398_
timestamp 1667941163
transform 1 0 11684 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1399_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1400_
timestamp 1667941163
transform 1 0 29900 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1401_
timestamp 1667941163
transform 1 0 7544 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1402_
timestamp 1667941163
transform 1 0 17664 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1403_
timestamp 1667941163
transform 1 0 14352 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1404_
timestamp 1667941163
transform 1 0 10856 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1405_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _1406_
timestamp 1667941163
transform 1 0 6624 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1407_
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1408_
timestamp 1667941163
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1408__177
timestamp 1667941163
transform 1 0 5796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1409_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1410_
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1411_
timestamp 1667941163
transform 1 0 9200 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1412_
timestamp 1667941163
transform 1 0 8096 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1413_
timestamp 1667941163
transform 1 0 5888 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1414_
timestamp 1667941163
transform 1 0 34868 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1415_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1416_
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1417_
timestamp 1667941163
transform 1 0 36432 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1418_
timestamp 1667941163
transform 1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1419_
timestamp 1667941163
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1420_
timestamp 1667941163
transform 1 0 6532 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1421_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1422_
timestamp 1667941163
transform 1 0 30820 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1423_
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1424__178
timestamp 1667941163
transform 1 0 35144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1424_
timestamp 1667941163
transform 1 0 33304 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1425_
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1426_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1427_
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1428_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1429_
timestamp 1667941163
transform 1 0 28980 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1430_
timestamp 1667941163
transform 1 0 30360 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1431_
timestamp 1667941163
transform 1 0 17664 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1432_
timestamp 1667941163
transform 1 0 23552 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1433_
timestamp 1667941163
transform 1 0 28336 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1434_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1435_
timestamp 1667941163
transform 1 0 28704 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1436_
timestamp 1667941163
transform 1 0 30820 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1437_
timestamp 1667941163
transform 1 0 28428 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1438_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1439_
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1440_
timestamp 1667941163
transform 1 0 9292 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1440__179
timestamp 1667941163
transform 1 0 9384 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1441_
timestamp 1667941163
transform 1 0 24656 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1442_
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1443_
timestamp 1667941163
transform 1 0 17112 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1444_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1445_
timestamp 1667941163
transform 1 0 22264 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1446_
timestamp 1667941163
transform 1 0 17296 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1447_
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1448_
timestamp 1667941163
transform 1 0 9936 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1449_
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1450_
timestamp 1667941163
transform 1 0 15732 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1451_
timestamp 1667941163
transform 1 0 25024 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1452_
timestamp 1667941163
transform 1 0 25116 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1453_
timestamp 1667941163
transform 1 0 23920 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1454_
timestamp 1667941163
transform 1 0 26772 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1455_
timestamp 1667941163
transform 1 0 22632 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1456__180
timestamp 1667941163
transform 1 0 30728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1456_
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1457_
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1458_
timestamp 1667941163
transform 1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1459_
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1460_
timestamp 1667941163
transform 1 0 32016 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1461_
timestamp 1667941163
transform 1 0 31372 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1462_
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1463_
timestamp 1667941163
transform 1 0 32292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1464_
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1465_
timestamp 1667941163
transform 1 0 30912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1466_
timestamp 1667941163
transform 1 0 31924 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1467_
timestamp 1667941163
transform 1 0 21712 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1468_
timestamp 1667941163
transform 1 0 25852 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1469_
timestamp 1667941163
transform 1 0 30084 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1470_
timestamp 1667941163
transform 1 0 33488 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1471_
timestamp 1667941163
transform 1 0 31372 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1472_
timestamp 1667941163
transform 1 0 32292 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1472__181
timestamp 1667941163
transform 1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1473_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1474_
timestamp 1667941163
transform 1 0 18676 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1475_
timestamp 1667941163
transform 1 0 7452 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1476_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1477_
timestamp 1667941163
transform 1 0 7820 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1478_
timestamp 1667941163
transform 1 0 34500 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1479_
timestamp 1667941163
transform 1 0 9844 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1480_
timestamp 1667941163
transform 1 0 22448 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1481_
timestamp 1667941163
transform 1 0 8188 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1482_
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1483_
timestamp 1667941163
transform 1 0 8188 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1484_
timestamp 1667941163
transform 1 0 16928 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1485_
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1486_
timestamp 1667941163
transform 1 0 25300 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1487_
timestamp 1667941163
transform 1 0 21712 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1488__182
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1488_
timestamp 1667941163
transform 1 0 31924 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1489_
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1490_
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1491_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1492_
timestamp 1667941163
transform 1 0 14352 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1493_
timestamp 1667941163
transform 1 0 22816 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1494_
timestamp 1667941163
transform 1 0 7360 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1495_
timestamp 1667941163
transform 1 0 20332 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1496_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1497_
timestamp 1667941163
transform 1 0 19780 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1498_
timestamp 1667941163
transform 1 0 23736 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1499_
timestamp 1667941163
transform 1 0 15732 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1500_
timestamp 1667941163
transform 1 0 9476 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1501_
timestamp 1667941163
transform 1 0 25300 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1502_
timestamp 1667941163
transform 1 0 19964 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1503_
timestamp 1667941163
transform 1 0 18124 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1504__183
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1504_
timestamp 1667941163
transform 1 0 6624 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1505_
timestamp 1667941163
transform 1 0 22908 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1506_
timestamp 1667941163
transform 1 0 17020 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1507_
timestamp 1667941163
transform 1 0 12788 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1508_
timestamp 1667941163
transform 1 0 29716 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1509_
timestamp 1667941163
transform 1 0 22724 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1510_
timestamp 1667941163
transform 1 0 29900 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1511_
timestamp 1667941163
transform 1 0 23092 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1512_
timestamp 1667941163
transform 1 0 11868 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1513_
timestamp 1667941163
transform 1 0 11316 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1514_
timestamp 1667941163
transform 1 0 17020 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1515_
timestamp 1667941163
transform 1 0 24472 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1516_
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1517_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1518_
timestamp 1667941163
transform 1 0 27232 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1519_
timestamp 1667941163
transform 1 0 23736 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1520__184
timestamp 1667941163
transform 1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1520_
timestamp 1667941163
transform 1 0 29900 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1521_
timestamp 1667941163
transform 1 0 9752 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1522_
timestamp 1667941163
transform 1 0 9384 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1523_
timestamp 1667941163
transform 1 0 3312 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1524_
timestamp 1667941163
transform 1 0 26864 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1525_
timestamp 1667941163
transform 1 0 32292 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1526_
timestamp 1667941163
transform 1 0 26680 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1527_
timestamp 1667941163
transform 1 0 28336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1528_
timestamp 1667941163
transform 1 0 31464 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1529_
timestamp 1667941163
transform 1 0 30452 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1530_
timestamp 1667941163
transform 1 0 29532 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1531_
timestamp 1667941163
transform 1 0 15088 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1532_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1533_
timestamp 1667941163
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1534_
timestamp 1667941163
transform 1 0 18492 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1535_
timestamp 1667941163
transform 1 0 21528 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1536__185
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1536_
timestamp 1667941163
transform 1 0 27876 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1537_
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1538_
timestamp 1667941163
transform 1 0 7176 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1539_
timestamp 1667941163
transform 1 0 7452 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1540_
timestamp 1667941163
transform 1 0 4876 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1541_
timestamp 1667941163
transform 1 0 7452 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1542_
timestamp 1667941163
transform 1 0 7452 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1543_
timestamp 1667941163
transform 1 0 5244 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1544_
timestamp 1667941163
transform 1 0 2668 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1545_
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1546_
timestamp 1667941163
transform 1 0 17756 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1547_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1548_
timestamp 1667941163
transform 1 0 8188 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1549_
timestamp 1667941163
transform 1 0 9568 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1550_
timestamp 1667941163
transform 1 0 33212 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1551_
timestamp 1667941163
transform 1 0 32292 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1552_
timestamp 1667941163
transform 1 0 31280 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1552__186
timestamp 1667941163
transform 1 0 34132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1553_
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1554_
timestamp 1667941163
transform 1 0 31096 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1555_
timestamp 1667941163
transform 1 0 33580 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1556_
timestamp 1667941163
transform 1 0 21160 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1557_
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1558_
timestamp 1667941163
transform 1 0 32660 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1559_
timestamp 1667941163
transform 1 0 26128 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1560_
timestamp 1667941163
transform 1 0 25024 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1561_
timestamp 1667941163
transform 1 0 29992 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1562_
timestamp 1667941163
transform 1 0 32384 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1563_
timestamp 1667941163
transform 1 0 29992 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1564_
timestamp 1667941163
transform 1 0 22448 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1565_
timestamp 1667941163
transform 1 0 27968 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1566_
timestamp 1667941163
transform 1 0 17848 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1567_
timestamp 1667941163
transform 1 0 10028 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1568__187
timestamp 1667941163
transform 1 0 8096 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1568_
timestamp 1667941163
transform 1 0 8004 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1667941163
transform 1 0 30728 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1667941163
transform 1 0 8924 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1572_
timestamp 1667941163
transform 1 0 28704 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1573_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1574_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1575_
timestamp 1667941163
transform 1 0 23460 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1576_
timestamp 1667941163
transform 1 0 9752 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1577_
timestamp 1667941163
transform 1 0 10028 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1578_
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1667941163
transform 1 0 7544 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1580_
timestamp 1667941163
transform 1 0 26864 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1581_
timestamp 1667941163
transform 1 0 23460 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1582_
timestamp 1667941163
transform 1 0 11776 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1583_
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1584_
timestamp 1667941163
transform 1 0 15824 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1585__188
timestamp 1667941163
transform 1 0 12328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1585_
timestamp 1667941163
transform 1 0 13616 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1586_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1587_
timestamp 1667941163
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1588_
timestamp 1667941163
transform 1 0 10212 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1589_
timestamp 1667941163
transform 1 0 9568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1590_
timestamp 1667941163
transform 1 0 10672 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1591_
timestamp 1667941163
transform 1 0 14904 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1592_
timestamp 1667941163
transform 1 0 10488 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1593_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1594_
timestamp 1667941163
transform 1 0 20148 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1595_
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1596_
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1597_
timestamp 1667941163
transform 1 0 16192 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1597__189
timestamp 1667941163
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1598_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1599_
timestamp 1667941163
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1600_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1601_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1602_
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1603_
timestamp 1667941163
transform 1 0 14996 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1604_
timestamp 1667941163
transform 1 0 11500 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1605_
timestamp 1667941163
transform 1 0 13616 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1606_
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1607_
timestamp 1667941163
transform 1 0 26864 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1608_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1609_
timestamp 1667941163
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1609__190
timestamp 1667941163
transform 1 0 28704 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1610_
timestamp 1667941163
transform 1 0 33856 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1611_
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1612_
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1613_
timestamp 1667941163
transform 1 0 17940 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1614_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1615_
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1616_
timestamp 1667941163
transform 1 0 16376 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1617_
timestamp 1667941163
transform 1 0 17204 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1618_
timestamp 1667941163
transform 1 0 15824 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1619_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1620_
timestamp 1667941163
transform 1 0 14444 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1621__191
timestamp 1667941163
transform 1 0 15548 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1621_
timestamp 1667941163
transform 1 0 14812 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1622_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1623_
timestamp 1667941163
transform 1 0 11408 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1624_
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1625_
timestamp 1667941163
transform 1 0 14444 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1626_
timestamp 1667941163
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1627_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1628_
timestamp 1667941163
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1629_
timestamp 1667941163
transform 1 0 13340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 11684 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 15364 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 17940 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 28244 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 29716 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 20516 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 27968 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 27232 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 36984 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 37444 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 20516 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform 1 0 14260 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 23368 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 38088 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform 1 0 26036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 38088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1667941163
transform 1 0 37444 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 28612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 5336 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 35604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1667941163
transform 1 0 15456 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1667941163
transform 1 0 10304 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1667941163
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 36708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1667941163
transform 1 0 37444 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1667941163
transform 1 0 37444 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 36708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1667941163
transform 1 0 36064 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1667941163
transform 1 0 37444 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1667941163
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1667941163
transform 1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1667941163
transform 1 0 34868 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1667941163
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 38088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1667941163
transform 1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1667941163
transform 1 0 1564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1667941163
transform 1 0 38088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1667941163
transform 1 0 28980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1667941163
transform 1 0 3036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1667941163
transform 1 0 7176 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1667941163
transform 1 0 28704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1667941163
transform 1 0 38088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 36708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 36340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 35880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 3036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1667941163
transform 1 0 36616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1667941163
transform 1 0 2300 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1667941163
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1667941163
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1667941163
transform 1 0 37260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1667941163
transform 1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1667941163
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1667941163
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1667941163
transform 1 0 18584 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1667941163
transform 1 0 2300 0 1 5440
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 2 nsew signal input
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 3 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 ccff_head
port 4 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal3 s 39200 31288 39800 31408 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 82 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 83 nsew signal input
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 84 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_bottom_in[12]
port 85 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 86 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 87 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 88 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 89 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 90 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chany_bottom_in[18]
port 91 nsew signal input
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 92 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 93 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 94 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 95 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 96 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 97 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 98 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 99 nsew signal input
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 100 nsew signal input
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 101 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 102 nsew signal tristate
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 103 nsew signal tristate
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 104 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 105 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 106 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 107 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 108 nsew signal tristate
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 109 nsew signal tristate
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 110 nsew signal tristate
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 111 nsew signal tristate
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 112 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 113 nsew signal tristate
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 114 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 115 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 116 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 117 nsew signal tristate
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 118 nsew signal tristate
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 119 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chany_top_in[0]
port 120 nsew signal input
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 121 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 122 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_top_in[12]
port 123 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 124 nsew signal input
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chany_top_in[14]
port 125 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_in[15]
port 126 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 127 nsew signal input
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 128 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 129 nsew signal input
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chany_top_in[1]
port 130 nsew signal input
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_in[2]
port 131 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chany_top_in[3]
port 132 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 133 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_top_in[5]
port 134 nsew signal input
flabel metal3 s 39200 12928 39800 13048 0 FreeSans 480 0 0 0 chany_top_in[6]
port 135 nsew signal input
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chany_top_in[7]
port 136 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_top_in[8]
port 137 nsew signal input
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_top_in[9]
port 138 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_out[0]
port 139 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 140 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_top_out[11]
port 141 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chany_top_out[12]
port 142 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 143 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 144 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_top_out[15]
port 145 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[16]
port 146 nsew signal tristate
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 147 nsew signal tristate
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 148 nsew signal tristate
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chany_top_out[1]
port 149 nsew signal tristate
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 150 nsew signal tristate
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 151 nsew signal tristate
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_top_out[4]
port 152 nsew signal tristate
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 153 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 154 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 155 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_top_out[8]
port 156 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_top_out[9]
port 157 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 158 nsew signal input
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 159 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 160 nsew signal input
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 161 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 pReset
port 162 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 prog_clk
port 163 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 164 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 165 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 166 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 167 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 168 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 169 nsew signal input
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 170 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 171 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 172 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 172 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 173 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 38272 11594 38272 11594 0 _0000_
rlabel metal1 33541 4590 33541 4590 0 _0001_
rlabel metal1 32752 10234 32752 10234 0 _0002_
rlabel metal2 26818 10846 26818 10846 0 _0003_
rlabel metal1 20608 7174 20608 7174 0 _0004_
rlabel metal2 25070 7208 25070 7208 0 _0005_
rlabel metal1 32522 3468 32522 3468 0 _0006_
rlabel metal2 34362 9248 34362 9248 0 _0007_
rlabel metal1 6217 3434 6217 3434 0 _0008_
rlabel metal1 5612 6630 5612 6630 0 _0009_
rlabel metal2 7866 3213 7866 3213 0 _0010_
rlabel metal1 7038 2312 7038 2312 0 _0011_
rlabel metal2 10902 3366 10902 3366 0 _0012_
rlabel metal2 8878 5321 8878 5321 0 _0013_
rlabel metal2 2070 5032 2070 5032 0 _0014_
rlabel metal2 17618 2108 17618 2108 0 _0015_
rlabel metal1 29571 3094 29571 3094 0 _0016_
rlabel metal1 16790 2482 16790 2482 0 _0017_
rlabel metal1 23644 9010 23644 9010 0 _0018_
rlabel metal1 21620 15878 21620 15878 0 _0019_
rlabel via1 12466 12155 12466 12155 0 _0020_
rlabel metal3 19527 12444 19527 12444 0 _0021_
rlabel metal1 17112 15334 17112 15334 0 _0022_
rlabel metal1 13202 15878 13202 15878 0 _0023_
rlabel metal1 11040 16422 11040 16422 0 _0024_
rlabel metal1 13011 8534 13011 8534 0 _0025_
rlabel metal1 15081 11798 15081 11798 0 _0026_
rlabel metal1 18538 10139 18538 10139 0 _0027_
rlabel metal1 19879 10710 19879 10710 0 _0028_
rlabel metal1 22133 12206 22133 12206 0 _0029_
rlabel metal1 28336 14858 28336 14858 0 _0030_
rlabel metal1 25852 15674 25852 15674 0 _0031_
rlabel via2 19366 13957 19366 13957 0 _0032_
rlabel metal2 19366 15266 19366 15266 0 _0033_
rlabel metal2 17710 14824 17710 14824 0 _0034_
rlabel metal2 13662 16320 13662 16320 0 _0035_
rlabel metal3 15157 16660 15157 16660 0 _0036_
rlabel metal1 21167 8534 21167 8534 0 _0037_
rlabel metal2 13846 14654 13846 14654 0 _0038_
rlabel metal1 16422 14858 16422 14858 0 _0039_
rlabel metal1 7307 4182 7307 4182 0 _0040_
rlabel metal2 3726 6256 3726 6256 0 _0041_
rlabel metal1 2254 4590 2254 4590 0 _0042_
rlabel metal1 2898 8874 2898 8874 0 _0043_
rlabel metal1 14766 11118 14766 11118 0 _0044_
rlabel metal1 15962 9350 15962 9350 0 _0045_
rlabel metal2 11960 9588 11960 9588 0 _0046_
rlabel metal1 13662 15538 13662 15538 0 _0047_
rlabel metal1 31648 7514 31648 7514 0 _0048_
rlabel metal2 31694 8602 31694 8602 0 _0049_
rlabel metal1 25346 15878 25346 15878 0 _0050_
rlabel metal1 28566 9513 28566 9513 0 _0051_
rlabel metal1 18538 14790 18538 14790 0 _0052_
rlabel metal1 15686 13498 15686 13498 0 _0053_
rlabel metal2 23966 13022 23966 13022 0 _0054_
rlabel via3 20355 10676 20355 10676 0 _0055_
rlabel metal3 16652 13668 16652 13668 0 _0056_
rlabel metal1 14996 15334 14996 15334 0 _0057_
rlabel metal2 15318 14144 15318 14144 0 _0058_
rlabel via3 10557 9588 10557 9588 0 _0059_
rlabel metal2 13938 11441 13938 11441 0 _0060_
rlabel metal1 24840 15334 24840 15334 0 _0061_
rlabel metal1 23927 13226 23927 13226 0 _0062_
rlabel metal1 27554 11798 27554 11798 0 _0063_
rlabel metal1 26680 14790 26680 14790 0 _0064_
rlabel metal1 27830 14790 27830 14790 0 _0065_
rlabel metal1 28520 14790 28520 14790 0 _0066_
rlabel metal1 24157 11118 24157 11118 0 _0067_
rlabel metal1 26036 15334 26036 15334 0 _0068_
rlabel metal1 24702 12070 24702 12070 0 _0069_
rlabel metal1 27055 14382 27055 14382 0 _0070_
rlabel metal1 28366 11050 28366 11050 0 _0071_
rlabel metal1 33396 10438 33396 10438 0 _0072_
rlabel metal1 35604 7990 35604 7990 0 _0073_
rlabel metal1 29309 2346 29309 2346 0 _0074_
rlabel metal1 23782 2346 23782 2346 0 _0075_
rlabel metal1 14943 3094 14943 3094 0 _0076_
rlabel metal2 18262 4845 18262 4845 0 _0077_
rlabel metal1 15686 7480 15686 7480 0 _0078_
rlabel metal2 31786 5950 31786 5950 0 _0079_
rlabel metal1 30038 6392 30038 6392 0 _0080_
rlabel metal2 35742 7565 35742 7565 0 _0081_
rlabel metal2 35650 8228 35650 8228 0 _0082_
rlabel metal1 19734 14926 19734 14926 0 _0083_
rlabel metal2 15318 11628 15318 11628 0 _0084_
rlabel metal2 18354 13974 18354 13974 0 _0085_
rlabel metal3 17204 13260 17204 13260 0 _0086_
rlabel metal2 34270 5729 34270 5729 0 _0087_
rlabel metal2 14398 17289 14398 17289 0 _0088_
rlabel metal2 17894 13668 17894 13668 0 _0089_
rlabel metal1 19550 7956 19550 7956 0 _0090_
rlabel metal1 16291 9554 16291 9554 0 _0091_
rlabel metal1 13110 13335 13110 13335 0 _0092_
rlabel metal1 20378 13158 20378 13158 0 _0093_
rlabel metal1 26634 12954 26634 12954 0 _0094_
rlabel metal1 29033 6698 29033 6698 0 _0095_
rlabel metal1 31425 6766 31425 6766 0 _0096_
rlabel metal1 30222 11526 30222 11526 0 _0097_
rlabel metal1 30038 8330 30038 8330 0 _0098_
rlabel metal2 23138 7480 23138 7480 0 _0099_
rlabel metal1 21167 2346 21167 2346 0 _0100_
rlabel metal1 27416 9894 27416 9894 0 _0101_
rlabel metal2 32982 7939 32982 7939 0 _0102_
rlabel metal2 31786 10200 31786 10200 0 _0103_
rlabel via2 33626 7803 33626 7803 0 _0104_
rlabel metal1 29302 13770 29302 13770 0 _0105_
rlabel metal2 16330 7973 16330 7973 0 _0106_
rlabel metal1 11093 2346 11093 2346 0 _0107_
rlabel metal1 17335 3094 17335 3094 0 _0108_
rlabel metal2 12558 5440 12558 5440 0 _0109_
rlabel metal2 15870 6851 15870 6851 0 _0110_
rlabel metal1 23736 15334 23736 15334 0 _0111_
rlabel metal2 31878 5321 31878 5321 0 _0112_
rlabel metal2 35006 8840 35006 8840 0 _0113_
rlabel metal1 32660 9350 32660 9350 0 _0114_
rlabel metal1 33580 8874 33580 8874 0 _0115_
rlabel metal2 27646 9010 27646 9010 0 _0116_
rlabel metal1 27147 13294 27147 13294 0 _0117_
rlabel metal1 24794 12614 24794 12614 0 _0118_
rlabel metal1 31004 14246 31004 14246 0 _0119_
rlabel metal2 13202 19720 13202 19720 0 _0120_
rlabel via2 15502 19771 15502 19771 0 _0121_
rlabel metal2 13294 18683 13294 18683 0 _0122_
rlabel metal1 9890 20298 9890 20298 0 _0123_
rlabel metal2 20102 4097 20102 4097 0 _0124_
rlabel metal2 29486 9214 29486 9214 0 _0125_
rlabel metal1 22310 4631 22310 4631 0 _0126_
rlabel metal2 35742 6545 35742 6545 0 _0127_
rlabel metal1 12834 14518 12834 14518 0 _0128_
rlabel metal1 15916 14246 15916 14246 0 _0129_
rlabel metal2 14674 12070 14674 12070 0 _0130_
rlabel metal2 12558 10081 12558 10081 0 _0131_
rlabel metal2 14030 13600 14030 13600 0 _0132_
rlabel metal2 13938 13435 13938 13435 0 _0133_
rlabel metal1 22586 18598 22586 18598 0 _0134_
rlabel metal2 20746 18377 20746 18377 0 _0135_
rlabel metal3 15985 16660 15985 16660 0 _0136_
rlabel metal1 16514 15878 16514 15878 0 _0137_
rlabel via3 12627 6868 12627 6868 0 _0138_
rlabel metal1 12880 16422 12880 16422 0 _0139_
rlabel metal1 36439 2346 36439 2346 0 _0140_
rlabel metal1 34277 2346 34277 2346 0 _0141_
rlabel metal1 31287 2346 31287 2346 0 _0142_
rlabel metal3 20286 12444 20286 12444 0 _0143_
rlabel via3 16261 15300 16261 15300 0 _0144_
rlabel metal2 12696 12172 12696 12172 0 _0145_
rlabel metal1 15180 11050 15180 11050 0 _0146_
rlabel metal1 12328 15334 12328 15334 0 _0147_
rlabel metal1 11914 15334 11914 15334 0 _0148_
rlabel metal2 12972 13260 12972 13260 0 _0149_
rlabel metal1 19780 13158 19780 13158 0 _0150_
rlabel metal2 19320 12988 19320 12988 0 _0151_
rlabel metal1 27508 17170 27508 17170 0 _0152_
rlabel metal1 20884 15470 20884 15470 0 _0153_
rlabel metal1 20240 7378 20240 7378 0 _0154_
rlabel metal1 2070 6766 2070 6766 0 _0155_
rlabel metal2 23782 14688 23782 14688 0 _0156_
rlabel metal2 29026 15232 29026 15232 0 _0157_
rlabel metal2 2622 9520 2622 9520 0 _0158_
rlabel metal1 17848 14994 17848 14994 0 _0159_
rlabel metal2 29670 15504 29670 15504 0 _0160_
rlabel metal1 20700 6290 20700 6290 0 _0161_
rlabel metal1 20378 15028 20378 15028 0 _0162_
rlabel metal1 20194 13294 20194 13294 0 _0163_
rlabel metal1 16054 10642 16054 10642 0 _0164_
rlabel metal1 33028 9554 33028 9554 0 _0165_
rlabel metal1 15962 14382 15962 14382 0 _0166_
rlabel metal1 20654 18700 20654 18700 0 _0167_
rlabel metal2 22034 17748 22034 17748 0 _0168_
rlabel metal2 32430 9690 32430 9690 0 _0169_
rlabel metal1 33488 7174 33488 7174 0 _0170_
rlabel metal2 26542 6086 26542 6086 0 _0171_
rlabel metal1 30682 10506 30682 10506 0 _0172_
rlabel metal1 20558 23766 20558 23766 0 _0173_
rlabel metal2 18630 19176 18630 19176 0 _0174_
rlabel metal1 28474 17714 28474 17714 0 _0175_
rlabel metal1 14904 20502 14904 20502 0 _0176_
rlabel metal2 13018 18632 13018 18632 0 _0177_
rlabel metal1 31510 16218 31510 16218 0 _0178_
rlabel metal1 24610 22678 24610 22678 0 _0179_
rlabel metal1 34592 5270 34592 5270 0 _0180_
rlabel metal2 31786 7667 31786 7667 0 _0181_
rlabel metal1 26956 23766 26956 23766 0 _0182_
rlabel metal1 31326 22406 31326 22406 0 _0183_
rlabel metal1 36432 11050 36432 11050 0 _0184_
rlabel metal1 4738 6970 4738 6970 0 _0185_
rlabel metal2 4738 8330 4738 8330 0 _0186_
rlabel metal1 6072 7990 6072 7990 0 _0187_
rlabel metal1 13984 16150 13984 16150 0 _0188_
rlabel metal1 7452 12886 7452 12886 0 _0189_
rlabel metal1 7130 16490 7130 16490 0 _0190_
rlabel metal1 6026 15368 6026 15368 0 _0191_
rlabel metal2 6854 10608 6854 10608 0 _0192_
rlabel metal2 6946 15742 6946 15742 0 _0193_
rlabel metal2 7222 11118 7222 11118 0 _0194_
rlabel metal2 4830 7140 4830 7140 0 _0195_
rlabel metal1 4922 9894 4922 9894 0 _0196_
rlabel metal1 5152 5270 5152 5270 0 _0197_
rlabel metal2 5934 14178 5934 14178 0 _0198_
rlabel metal2 7590 11560 7590 11560 0 _0199_
rlabel via1 5470 8534 5470 8534 0 _0200_
rlabel metal1 33442 8942 33442 8942 0 _0201_
rlabel metal1 24150 16150 24150 16150 0 _0202_
rlabel metal1 34178 7718 34178 7718 0 _0203_
rlabel metal2 11822 21794 11822 21794 0 _0204_
rlabel metal1 11040 19414 11040 19414 0 _0205_
rlabel metal1 18446 24718 18446 24718 0 _0206_
rlabel metal2 33166 16728 33166 16728 0 _0207_
rlabel metal1 31970 20434 31970 20434 0 _0208_
rlabel metal1 30590 16218 30590 16218 0 _0209_
rlabel metal2 13386 23630 13386 23630 0 _0210_
rlabel metal1 13984 24650 13984 24650 0 _0211_
rlabel viali 28286 24106 28286 24106 0 _0212_
rlabel metal2 22586 16830 22586 16830 0 _0213_
rlabel metal2 16054 24616 16054 24616 0 _0214_
rlabel metal2 21482 19992 21482 19992 0 _0215_
rlabel metal2 14490 27914 14490 27914 0 _0216_
rlabel metal1 19780 19414 19780 19414 0 _0217_
rlabel metal1 20194 21658 20194 21658 0 _0218_
rlabel metal1 13294 20570 13294 20570 0 _0219_
rlabel metal2 24794 26520 24794 26520 0 _0220_
rlabel metal2 18814 26792 18814 26792 0 _0221_
rlabel metal1 18354 27336 18354 27336 0 _0222_
rlabel metal1 23000 22678 23000 22678 0 _0223_
rlabel metal2 18906 20910 18906 20910 0 _0224_
rlabel metal1 25944 21930 25944 21930 0 _0225_
rlabel metal1 26772 26282 26772 26282 0 _0226_
rlabel metal2 29946 25466 29946 25466 0 _0227_
rlabel metal2 24794 27880 24794 27880 0 _0228_
rlabel metal1 20194 20570 20194 20570 0 _0229_
rlabel via1 26358 24803 26358 24803 0 _0230_
rlabel metal1 35098 4182 35098 4182 0 _0231_
rlabel metal1 29946 22984 29946 22984 0 _0232_
rlabel metal2 19366 21777 19366 21777 0 _0233_
rlabel metal1 19550 22746 19550 22746 0 _0234_
rlabel metal1 19734 32470 19734 32470 0 _0235_
rlabel metal2 21298 28696 21298 28696 0 _0236_
rlabel metal2 21206 24616 21206 24616 0 _0237_
rlabel metal1 15456 22678 15456 22678 0 _0238_
rlabel metal2 22862 28016 22862 28016 0 _0239_
rlabel metal2 11086 23936 11086 23936 0 _0240_
rlabel metal1 11408 17238 11408 17238 0 _0241_
rlabel metal1 30728 18054 30728 18054 0 _0242_
rlabel metal1 30636 10098 30636 10098 0 _0243_
rlabel metal1 7728 5118 7728 5118 0 _0244_
rlabel metal1 17618 22406 17618 22406 0 _0245_
rlabel metal2 16054 30056 16054 30056 0 _0246_
rlabel metal1 11638 30362 11638 30362 0 _0247_
rlabel metal2 24334 24208 24334 24208 0 _0248_
rlabel metal1 7176 11662 7176 11662 0 _0249_
rlabel metal2 5750 10472 5750 10472 0 _0250_
rlabel metal2 6302 11016 6302 11016 0 _0251_
rlabel metal2 9338 17816 9338 17816 0 _0252_
rlabel metal1 15778 16456 15778 16456 0 _0253_
rlabel metal1 8464 14246 8464 14246 0 _0254_
rlabel metal1 8234 14042 8234 14042 0 _0255_
rlabel metal1 5382 7514 5382 7514 0 _0256_
rlabel metal1 33442 3944 33442 3944 0 _0257_
rlabel metal1 25806 16762 25806 16762 0 _0258_
rlabel metal2 9338 3298 9338 3298 0 _0259_
rlabel metal2 30130 5389 30130 5389 0 _0260_
rlabel metal1 9338 9044 9338 9044 0 _0261_
rlabel metal2 7038 17374 7038 17374 0 _0262_
rlabel metal1 6670 17850 6670 17850 0 _0263_
rlabel metal1 9338 16456 9338 16456 0 _0264_
rlabel metal1 29946 18258 29946 18258 0 _0265_
rlabel metal1 31004 17306 31004 17306 0 _0266_
rlabel metal1 32936 15130 32936 15130 0 _0267_
rlabel metal1 15042 23766 15042 23766 0 _0268_
rlabel metal2 17066 20638 17066 20638 0 _0269_
rlabel metal2 18262 23970 18262 23970 0 _0270_
rlabel metal2 29946 19278 29946 19278 0 _0271_
rlabel metal2 26818 30056 26818 30056 0 _0272_
rlabel metal1 32706 20808 32706 20808 0 _0273_
rlabel metal1 17756 27642 17756 27642 0 _0274_
rlabel metal2 23782 29614 23782 29614 0 _0275_
rlabel metal2 28566 22814 28566 22814 0 _0276_
rlabel metal1 29762 16490 29762 16490 0 _0277_
rlabel metal2 30406 20910 30406 20910 0 _0278_
rlabel metal1 30866 28662 30866 28662 0 _0279_
rlabel metal2 28658 28254 28658 28254 0 _0280_
rlabel metal1 16376 21590 16376 21590 0 _0281_
rlabel metal1 17480 20026 17480 20026 0 _0282_
rlabel metal1 11500 18598 11500 18598 0 _0283_
rlabel metal2 24886 28254 24886 28254 0 _0284_
rlabel metal1 24472 24378 24472 24378 0 _0285_
rlabel metal1 17158 26010 17158 26010 0 _0286_
rlabel metal2 21942 30056 21942 30056 0 _0287_
rlabel metal1 22862 23018 22862 23018 0 _0288_
rlabel metal2 17526 23256 17526 23256 0 _0289_
rlabel metal2 23138 27166 23138 27166 0 _0290_
rlabel metal1 10442 13498 10442 13498 0 _0291_
rlabel metal1 11914 21114 11914 21114 0 _0292_
rlabel metal1 16054 20026 16054 20026 0 _0293_
rlabel metal1 25438 23494 25438 23494 0 _0294_
rlabel metal2 25346 29410 25346 29410 0 _0295_
rlabel metal1 24150 20536 24150 20536 0 _0296_
rlabel metal1 28704 21046 28704 21046 0 _0297_
rlabel metal1 23230 25194 23230 25194 0 _0298_
rlabel metal1 32062 19380 32062 19380 0 _0299_
rlabel metal2 21482 25432 21482 25432 0 _0300_
rlabel metal1 21206 27404 21206 27404 0 _0301_
rlabel metal2 19550 23392 19550 23392 0 _0302_
rlabel metal2 32246 23970 32246 23970 0 _0303_
rlabel metal2 31602 25704 31602 25704 0 _0304_
rlabel metal2 13846 23902 13846 23902 0 _0305_
rlabel metal1 33396 18326 33396 18326 0 _0306_
rlabel metal1 30130 14042 30130 14042 0 _0307_
rlabel metal1 32384 17306 32384 17306 0 _0308_
rlabel metal1 33074 22950 33074 22950 0 _0309_
rlabel metal1 21942 27336 21942 27336 0 _0310_
rlabel metal1 26220 28458 26220 28458 0 _0311_
rlabel metal1 30360 23834 30360 23834 0 _0312_
rlabel metal1 34546 5610 34546 5610 0 _0313_
rlabel metal1 34868 5814 34868 5814 0 _0314_
rlabel metal1 32568 7446 32568 7446 0 _0315_
rlabel metal1 28980 15674 28980 15674 0 _0316_
rlabel metal1 18538 16150 18538 16150 0 _0317_
rlabel metal1 7682 13192 7682 13192 0 _0318_
rlabel metal1 24610 3162 24610 3162 0 _0319_
rlabel metal1 8234 7446 8234 7446 0 _0320_
rlabel metal1 34730 3128 34730 3128 0 _0321_
rlabel metal1 10074 5304 10074 5304 0 _0322_
rlabel metal1 13386 2074 13386 2074 0 _0323_
rlabel metal1 8372 10710 8372 10710 0 _0324_
rlabel metal2 31878 4386 31878 4386 0 _0325_
rlabel metal1 8602 14042 8602 14042 0 _0326_
rlabel metal1 16882 6358 16882 6358 0 _0327_
rlabel metal1 9798 13498 9798 13498 0 _0328_
rlabel metal2 25530 17289 25530 17289 0 _0329_
rlabel metal2 21942 18088 21942 18088 0 _0330_
rlabel metal1 32522 6698 32522 6698 0 _0331_
rlabel metal1 12098 22984 12098 22984 0 _0332_
rlabel metal2 11178 19720 11178 19720 0 _0333_
rlabel metal2 14490 25466 14490 25466 0 _0334_
rlabel metal2 14582 26792 14582 26792 0 _0335_
rlabel metal2 23046 19992 23046 19992 0 _0336_
rlabel metal1 8878 26554 8878 26554 0 _0337_
rlabel metal1 20516 27030 20516 27030 0 _0338_
rlabel metal1 23000 19414 23000 19414 0 _0339_
rlabel metal1 19872 24854 19872 24854 0 _0340_
rlabel metal2 25346 17442 25346 17442 0 _0341_
rlabel metal2 15916 23018 15916 23018 0 _0342_
rlabel metal2 9706 6919 9706 6919 0 _0343_
rlabel metal1 25760 24378 25760 24378 0 _0344_
rlabel metal2 19458 16269 19458 16269 0 _0345_
rlabel metal2 18354 17646 18354 17646 0 _0346_
rlabel metal2 6854 15096 6854 15096 0 _0347_
rlabel metal1 23138 24072 23138 24072 0 _0348_
rlabel metal2 17618 26520 17618 26520 0 _0349_
rlabel metal1 11914 26486 11914 26486 0 _0350_
rlabel metal1 29946 26248 29946 26248 0 _0351_
rlabel metal2 22954 26010 22954 26010 0 _0352_
rlabel metal2 30498 16575 30498 16575 0 _0353_
rlabel metal2 23322 28254 23322 28254 0 _0354_
rlabel metal2 12098 24327 12098 24327 0 _0355_
rlabel metal2 11546 28696 11546 28696 0 _0356_
rlabel metal1 17296 16150 17296 16150 0 _0357_
rlabel metal1 26266 26554 26266 26554 0 _0358_
rlabel metal2 27922 27608 27922 27608 0 _0359_
rlabel metal1 24472 18938 24472 18938 0 _0360_
rlabel metal1 27186 15674 27186 15674 0 _0361_
rlabel metal2 23966 17374 23966 17374 0 _0362_
rlabel metal1 33028 24038 33028 24038 0 _0363_
rlabel metal1 10304 12614 10304 12614 0 _0364_
rlabel metal2 9614 9656 9614 9656 0 _0365_
rlabel metal2 3542 6222 3542 6222 0 _0366_
rlabel metal1 27186 19754 27186 19754 0 _0367_
rlabel metal1 34224 20026 34224 20026 0 _0368_
rlabel metal2 32430 18462 32430 18462 0 _0369_
rlabel metal1 29302 21590 29302 21590 0 _0370_
rlabel metal2 33074 17408 33074 17408 0 _0371_
rlabel metal2 30682 15198 30682 15198 0 _0372_
rlabel metal1 32614 17646 32614 17646 0 _0373_
rlabel metal1 15272 17238 15272 17238 0 _0374_
rlabel metal1 30038 19754 30038 19754 0 _0375_
rlabel metal2 32430 21726 32430 21726 0 _0376_
rlabel metal1 17986 14586 17986 14586 0 _0377_
rlabel metal2 22218 17272 22218 17272 0 _0378_
rlabel metal1 28474 19482 28474 19482 0 _0379_
rlabel metal1 9338 4488 9338 4488 0 _0380_
rlabel metal1 7452 14042 7452 14042 0 _0381_
rlabel via2 5382 8075 5382 8075 0 _0382_
rlabel metal1 4232 6358 4232 6358 0 _0383_
rlabel via2 7682 9979 7682 9979 0 _0384_
rlabel metal1 7636 14314 7636 14314 0 _0385_
rlabel metal2 5474 5882 5474 5882 0 _0386_
rlabel metal2 2714 8585 2714 8585 0 _0387_
rlabel metal2 2622 5100 2622 5100 0 _0388_
rlabel metal2 17940 14314 17940 14314 0 _0389_
rlabel metal1 22172 21658 22172 21658 0 _0390_
rlabel metal2 8418 11934 8418 11934 0 _0391_
rlabel metal2 9798 16184 9798 16184 0 _0392_
rlabel metal1 33028 15334 33028 15334 0 _0393_
rlabel metal1 31694 16116 31694 16116 0 _0394_
rlabel metal1 35742 7446 35742 7446 0 _0395_
rlabel metal1 32522 20026 32522 20026 0 _0396_
rlabel metal2 31326 19907 31326 19907 0 _0397_
rlabel metal1 33442 24786 33442 24786 0 _0398_
rlabel metal2 21390 26520 21390 26520 0 _0399_
rlabel metal2 22310 21080 22310 21080 0 _0400_
rlabel metal1 33488 18666 33488 18666 0 _0401_
rlabel metal1 26404 27370 26404 27370 0 _0402_
rlabel metal1 25760 19414 25760 19414 0 _0403_
rlabel metal1 30636 22678 30636 22678 0 _0404_
rlabel metal1 32200 15674 32200 15674 0 _0405_
rlabel metal2 30498 27846 30498 27846 0 _0406_
rlabel metal2 23966 24038 23966 24038 0 _0407_
rlabel metal1 28934 27030 28934 27030 0 _0408_
rlabel metal1 17526 17306 17526 17306 0 _0409_
rlabel metal1 10488 12410 10488 12410 0 _0410_
rlabel metal2 8234 17374 8234 17374 0 _0411_
rlabel metal2 30912 4182 30912 4182 0 _0412_
rlabel metal1 25990 20978 25990 20978 0 _0413_
rlabel metal1 9154 4012 9154 4012 0 _0414_
rlabel metal1 28704 23290 28704 23290 0 _0415_
rlabel metal1 24748 21114 24748 21114 0 _0416_
rlabel metal2 22218 20910 22218 20910 0 _0417_
rlabel via1 23686 19414 23686 19414 0 _0418_
rlabel metal1 9975 11832 9975 11832 0 _0419_
rlabel metal1 10350 21658 10350 21658 0 _0420_
rlabel metal1 11500 14042 11500 14042 0 _0421_
rlabel metal2 7774 22814 7774 22814 0 _0422_
rlabel metal2 27830 24242 27830 24242 0 _0423_
rlabel metal2 23966 21352 23966 21352 0 _0424_
rlabel metal2 12650 22474 12650 22474 0 _0425_
rlabel metal1 14398 19482 14398 19482 0 _0426_
rlabel via1 16050 26282 16050 26282 0 _0427_
rlabel metal1 13478 29206 13478 29206 0 _0428_
rlabel metal1 13202 25840 13202 25840 0 _0429_
rlabel metal2 13294 24990 13294 24990 0 _0430_
rlabel metal2 11086 27812 11086 27812 0 _0431_
rlabel metal2 9798 27268 9798 27268 0 _0432_
rlabel metal1 12420 18394 12420 18394 0 _0433_
rlabel metal2 15134 28968 15134 28968 0 _0434_
rlabel metal1 10350 25874 10350 25874 0 _0435_
rlabel metal2 9338 29444 9338 29444 0 _0436_
rlabel metal2 21114 18088 21114 18088 0 _0437_
rlabel metal2 20930 16745 20930 16745 0 _0438_
rlabel metal1 20194 21930 20194 21930 0 _0439_
rlabel metal1 16606 21930 16606 21930 0 _0440_
rlabel metal1 19642 19720 19642 19720 0 _0441_
rlabel metal2 12190 20366 12190 20366 0 _0442_
rlabel metal1 19504 18666 19504 18666 0 _0443_
rlabel metal1 13754 21862 13754 21862 0 _0444_
rlabel metal1 19826 17544 19826 17544 0 _0445_
rlabel metal1 15226 21896 15226 21896 0 _0446_
rlabel metal2 11730 19992 11730 19992 0 _0447_
rlabel metal1 13478 21590 13478 21590 0 _0448_
rlabel metal1 33994 5882 33994 5882 0 _0449_
rlabel metal1 28198 9146 28198 9146 0 _0450_
rlabel metal2 27370 22814 27370 22814 0 _0451_
rlabel metal1 28750 21624 28750 21624 0 _0452_
rlabel metal1 33936 6358 33936 6358 0 _0453_
rlabel metal1 30038 8534 30038 8534 0 _0454_
rlabel metal2 23000 18666 23000 18666 0 _0455_
rlabel metal1 18308 22406 18308 22406 0 _0456_
rlabel metal1 28290 19346 28290 19346 0 _0457_
rlabel metal1 16744 20570 16744 20570 0 _0458_
rlabel metal1 16606 17544 16606 17544 0 _0459_
rlabel metal1 17250 18938 17250 18938 0 _0460_
rlabel metal1 14996 21114 14996 21114 0 _0461_
rlabel metal1 16652 30294 16652 30294 0 _0462_
rlabel metal1 13524 30294 13524 30294 0 _0463_
rlabel metal2 15410 30260 15410 30260 0 _0464_
rlabel metal1 12052 26962 12052 26962 0 _0465_
rlabel metal1 10626 25330 10626 25330 0 _0466_
rlabel metal2 15042 29580 15042 29580 0 _0467_
rlabel metal1 15042 28050 15042 28050 0 _0468_
rlabel metal1 13800 23290 13800 23290 0 _0469_
rlabel metal1 14444 26418 14444 26418 0 _0470_
rlabel metal1 10580 27098 10580 27098 0 _0471_
rlabel metal2 13570 27778 13570 27778 0 _0472_
rlabel metal3 1234 30668 1234 30668 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 37214 8908 37214 8908 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 1234 22508 1234 22508 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25162 823 25162 823 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 29026 4784 29026 4784 0 ccff_head
rlabel metal1 2944 37094 2944 37094 0 ccff_tail
rlabel metal1 37766 37298 37766 37298 0 chanx_left_in[0]
rlabel metal1 33902 2890 33902 2890 0 chanx_left_in[10]
rlabel metal1 16928 36754 16928 36754 0 chanx_left_in[11]
rlabel metal2 32430 4828 32430 4828 0 chanx_left_in[12]
rlabel metal2 17710 3366 17710 3366 0 chanx_left_in[13]
rlabel metal1 8004 5270 8004 5270 0 chanx_left_in[14]
rlabel metal3 1234 17748 1234 17748 0 chanx_left_in[15]
rlabel metal1 14260 36754 14260 36754 0 chanx_left_in[16]
rlabel metal2 16146 38226 16146 38226 0 chanx_left_in[17]
rlabel metal1 3726 37230 3726 37230 0 chanx_left_in[18]
rlabel metal3 1280 748 1280 748 0 chanx_left_in[1]
rlabel metal1 23368 37230 23368 37230 0 chanx_left_in[2]
rlabel metal1 38364 10030 38364 10030 0 chanx_left_in[3]
rlabel metal1 25990 37230 25990 37230 0 chanx_left_in[4]
rlabel metal3 1188 2788 1188 2788 0 chanx_left_in[5]
rlabel metal1 18032 37230 18032 37230 0 chanx_left_in[6]
rlabel metal1 9798 37230 9798 37230 0 chanx_left_in[7]
rlabel metal2 38318 17119 38318 17119 0 chanx_left_in[8]
rlabel metal1 2714 3094 2714 3094 0 chanx_left_in[9]
rlabel metal3 38786 36788 38786 36788 0 chanx_left_out[0]
rlabel metal1 4738 37094 4738 37094 0 chanx_left_out[10]
rlabel metal1 30268 3366 30268 3366 0 chanx_left_out[11]
rlabel metal3 1234 20468 1234 20468 0 chanx_left_out[12]
rlabel metal1 36386 4454 36386 4454 0 chanx_left_out[13]
rlabel metal2 38226 25177 38226 25177 0 chanx_left_out[14]
rlabel via2 38226 33371 38226 33371 0 chanx_left_out[15]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[16]
rlabel metal1 25346 37094 25346 37094 0 chanx_left_out[17]
rlabel metal3 1234 14348 1234 14348 0 chanx_left_out[18]
rlabel metal1 36340 37094 36340 37094 0 chanx_left_out[1]
rlabel metal1 1564 36890 1564 36890 0 chanx_left_out[2]
rlabel metal3 1234 19108 1234 19108 0 chanx_left_out[3]
rlabel metal2 38226 31637 38226 31637 0 chanx_left_out[4]
rlabel metal1 7912 37094 7912 37094 0 chanx_left_out[5]
rlabel metal1 2714 36890 2714 36890 0 chanx_left_out[6]
rlabel metal1 32384 36890 32384 36890 0 chanx_left_out[7]
rlabel metal1 38272 6630 38272 6630 0 chanx_left_out[8]
rlabel metal2 10350 1384 10350 1384 0 chanx_left_out[9]
rlabel metal1 38088 4046 38088 4046 0 chanx_right_in[0]
rlabel metal2 38134 30107 38134 30107 0 chanx_right_in[10]
rlabel metal2 23874 1231 23874 1231 0 chanx_right_in[11]
rlabel metal3 1142 36788 1142 36788 0 chanx_right_in[12]
rlabel metal2 38318 20689 38318 20689 0 chanx_right_in[13]
rlabel metal3 1142 12988 1142 12988 0 chanx_right_in[14]
rlabel metal2 38318 21913 38318 21913 0 chanx_right_in[15]
rlabel metal2 18078 1761 18078 1761 0 chanx_right_in[16]
rlabel metal1 37168 36822 37168 36822 0 chanx_right_in[17]
rlabel metal2 14858 1761 14858 1761 0 chanx_right_in[18]
rlabel metal3 1188 5508 1188 5508 0 chanx_right_in[1]
rlabel metal3 1234 24548 1234 24548 0 chanx_right_in[2]
rlabel metal1 5382 37230 5382 37230 0 chanx_right_in[3]
rlabel metal1 35374 37230 35374 37230 0 chanx_right_in[4]
rlabel metal3 1142 32028 1142 32028 0 chanx_right_in[5]
rlabel metal2 15502 38260 15502 38260 0 chanx_right_in[6]
rlabel metal2 16790 1761 16790 1761 0 chanx_right_in[7]
rlabel metal3 38694 12308 38694 12308 0 chanx_right_in[8]
rlabel metal2 10350 38260 10350 38260 0 chanx_right_in[9]
rlabel metal1 24702 37094 24702 37094 0 chanx_right_out[0]
rlabel metal1 11776 36890 11776 36890 0 chanx_right_out[10]
rlabel via2 38226 24565 38226 24565 0 chanx_right_out[11]
rlabel metal3 1234 28628 1234 28628 0 chanx_right_out[12]
rlabel metal1 34822 37094 34822 37094 0 chanx_right_out[13]
rlabel metal3 1234 21828 1234 21828 0 chanx_right_out[14]
rlabel metal2 38226 34833 38226 34833 0 chanx_right_out[15]
rlabel metal2 38226 14297 38226 14297 0 chanx_right_out[16]
rlabel metal1 3220 36890 3220 36890 0 chanx_right_out[17]
rlabel metal2 1334 2880 1334 2880 0 chanx_right_out[18]
rlabel metal1 5635 2550 5635 2550 0 chanx_right_out[1]
rlabel metal3 1234 31348 1234 31348 0 chanx_right_out[2]
rlabel metal3 1234 15708 1234 15708 0 chanx_right_out[3]
rlabel metal3 1234 10948 1234 10948 0 chanx_right_out[4]
rlabel metal1 36248 3910 36248 3910 0 chanx_right_out[5]
rlabel metal1 36156 36890 36156 36890 0 chanx_right_out[6]
rlabel metal2 21298 823 21298 823 0 chanx_right_out[7]
rlabel metal2 38226 15793 38226 15793 0 chanx_right_out[8]
rlabel metal2 38226 8857 38226 8857 0 chanx_right_out[9]
rlabel metal1 37260 36074 37260 36074 0 chany_bottom_in[0]
rlabel metal2 18722 1503 18722 1503 0 chany_bottom_in[10]
rlabel metal2 29670 1180 29670 1180 0 chany_bottom_in[11]
rlabel metal2 37490 32181 37490 32181 0 chany_bottom_in[12]
rlabel metal2 13570 2608 13570 2608 0 chany_bottom_in[13]
rlabel metal3 1188 36108 1188 36108 0 chany_bottom_in[14]
rlabel metal1 9200 36754 9200 36754 0 chany_bottom_in[15]
rlabel metal1 38410 4658 38410 4658 0 chany_bottom_in[16]
rlabel metal2 38134 10455 38134 10455 0 chany_bottom_in[17]
rlabel metal1 2438 10608 2438 10608 0 chany_bottom_in[18]
rlabel metal2 38134 18003 38134 18003 0 chany_bottom_in[1]
rlabel metal2 36754 1761 36754 1761 0 chany_bottom_in[2]
rlabel metal1 30544 37230 30544 37230 0 chany_bottom_in[3]
rlabel via2 38134 19771 38134 19771 0 chany_bottom_in[4]
rlabel metal3 1142 17068 1142 17068 0 chany_bottom_in[5]
rlabel metal3 1188 12308 1188 12308 0 chany_bottom_in[6]
rlabel metal1 21758 37230 21758 37230 0 chany_bottom_in[7]
rlabel metal1 26726 3094 26726 3094 0 chany_bottom_in[8]
rlabel metal1 35144 2890 35144 2890 0 chany_bottom_in[9]
rlabel metal2 38226 36057 38226 36057 0 chany_bottom_out[0]
rlabel metal3 1234 35428 1234 35428 0 chany_bottom_out[10]
rlabel metal1 22724 37094 22724 37094 0 chany_bottom_out[11]
rlabel metal3 1234 7548 1234 7548 0 chany_bottom_out[12]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[13]
rlabel metal2 690 2370 690 2370 0 chany_bottom_out[14]
rlabel metal2 5842 1622 5842 1622 0 chany_bottom_out[15]
rlabel metal2 36846 4573 36846 4573 0 chany_bottom_out[16]
rlabel metal1 1610 36346 1610 36346 0 chany_bottom_out[17]
rlabel metal2 38226 29393 38226 29393 0 chany_bottom_out[18]
rlabel metal1 12512 37094 12512 37094 0 chany_bottom_out[1]
rlabel metal1 29808 37094 29808 37094 0 chany_bottom_out[2]
rlabel metal2 4554 1690 4554 1690 0 chany_bottom_out[3]
rlabel metal2 38226 8279 38226 8279 0 chany_bottom_out[4]
rlabel via2 38226 22491 38226 22491 0 chany_bottom_out[5]
rlabel metal1 14030 37094 14030 37094 0 chany_bottom_out[6]
rlabel metal2 38226 15181 38226 15181 0 chany_bottom_out[7]
rlabel metal3 38418 748 38418 748 0 chany_bottom_out[8]
rlabel metal2 20654 1761 20654 1761 0 chany_bottom_out[9]
rlabel metal1 37352 29070 37352 29070 0 chany_top_in[0]
rlabel metal1 31970 37298 31970 37298 0 chany_top_in[10]
rlabel metal2 9706 1761 9706 1761 0 chany_top_in[11]
rlabel metal2 38134 10999 38134 10999 0 chany_top_in[12]
rlabel metal2 28566 7514 28566 7514 0 chany_top_in[13]
rlabel metal3 37498 1428 37498 1428 0 chany_top_in[14]
rlabel metal3 1234 23868 1234 23868 0 chany_top_in[15]
rlabel metal2 33534 823 33534 823 0 chany_top_in[16]
rlabel metal1 4324 3162 4324 3162 0 chany_top_in[17]
rlabel metal2 16192 5100 16192 5100 0 chany_top_in[18]
rlabel metal3 1188 15028 1188 15028 0 chany_top_in[1]
rlabel metal1 37352 34510 37352 34510 0 chany_top_in[2]
rlabel metal2 38318 24021 38318 24021 0 chany_top_in[3]
rlabel metal1 36156 2822 36156 2822 0 chany_top_in[4]
rlabel metal3 1142 19788 1142 19788 0 chany_top_in[5]
rlabel metal2 38318 13141 38318 13141 0 chany_top_in[6]
rlabel metal3 1234 26588 1234 26588 0 chany_top_in[7]
rlabel metal3 1234 9588 1234 9588 0 chany_top_in[8]
rlabel metal1 36800 36754 36800 36754 0 chany_top_in[9]
rlabel metal1 38134 5542 38134 5542 0 chany_top_out[0]
rlabel metal1 37720 36346 37720 36346 0 chany_top_out[10]
rlabel metal3 1234 27268 1234 27268 0 chany_top_out[11]
rlabel metal3 1234 29308 1234 29308 0 chany_top_out[12]
rlabel metal1 24012 3366 24012 3366 0 chany_top_out[13]
rlabel metal2 46 1044 46 1044 0 chany_top_out[14]
rlabel metal3 1234 3468 1234 3468 0 chany_top_out[15]
rlabel metal3 1234 33388 1234 33388 0 chany_top_out[16]
rlabel metal1 6302 37094 6302 37094 0 chany_top_out[17]
rlabel metal1 20838 37094 20838 37094 0 chany_top_out[18]
rlabel metal3 1234 25228 1234 25228 0 chany_top_out[1]
rlabel metal2 7130 1571 7130 1571 0 chany_top_out[2]
rlabel metal2 2622 2064 2622 2064 0 chany_top_out[3]
rlabel metal3 1234 6188 1234 6188 0 chany_top_out[4]
rlabel metal1 18768 37094 18768 37094 0 chany_top_out[5]
rlabel metal1 19504 6630 19504 6630 0 chany_top_out[6]
rlabel metal1 33672 37094 33672 37094 0 chany_top_out[7]
rlabel metal2 38226 7633 38226 7633 0 chany_top_out[8]
rlabel metal3 1096 1428 1096 1428 0 chany_top_out[9]
rlabel metal1 19734 4590 19734 4590 0 clknet_0_prog_clk
rlabel metal1 6808 2482 6808 2482 0 clknet_4_0_0_prog_clk
rlabel metal1 33626 2482 33626 2482 0 clknet_4_10_0_prog_clk
rlabel metal2 29394 7616 29394 7616 0 clknet_4_11_0_prog_clk
rlabel metal2 20838 9520 20838 9520 0 clknet_4_12_0_prog_clk
rlabel metal1 21252 12750 21252 12750 0 clknet_4_13_0_prog_clk
rlabel metal2 27186 9792 27186 9792 0 clknet_4_14_0_prog_clk
rlabel metal1 27002 13838 27002 13838 0 clknet_4_15_0_prog_clk
rlabel metal1 7038 6290 7038 6290 0 clknet_4_1_0_prog_clk
rlabel metal1 19826 2482 19826 2482 0 clknet_4_2_0_prog_clk
rlabel metal1 17020 4658 17020 4658 0 clknet_4_3_0_prog_clk
rlabel metal1 14444 10098 14444 10098 0 clknet_4_4_0_prog_clk
rlabel metal2 13110 13396 13110 13396 0 clknet_4_5_0_prog_clk
rlabel metal1 17020 10030 17020 10030 0 clknet_4_6_0_prog_clk
rlabel metal2 16882 14178 16882 14178 0 clknet_4_7_0_prog_clk
rlabel metal1 21482 2482 21482 2482 0 clknet_4_8_0_prog_clk
rlabel metal2 22034 4080 22034 4080 0 clknet_4_9_0_prog_clk
rlabel metal2 38318 27353 38318 27353 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 7774 1761 7774 1761 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 14214 1571 14214 1571 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal3 1050 8228 1050 8228 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 24610 14489 24610 14489 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal1 29670 14858 29670 14858 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal2 31878 24684 31878 24684 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 21114 10438 21114 10438 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 20516 19652 20516 19652 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 33534 18734 33534 18734 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 26680 13838 26680 13838 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal1 23920 14042 23920 14042 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal2 21390 9146 21390 9146 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal1 35098 4250 35098 4250 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal2 21022 7684 21022 7684 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 17940 13158 17940 13158 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 21850 20162 21850 20162 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal1 16376 10098 16376 10098 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal1 20378 8364 20378 8364 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal3 27347 18156 27347 18156 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal2 21666 15589 21666 15589 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal2 28934 6868 28934 6868 0 mem_bottom_track_17.DFFR_7_.Q
rlabel metal1 24564 18734 24564 18734 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 19734 11356 19734 11356 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 21620 13770 21620 13770 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal2 21114 15572 21114 15572 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal1 16606 16626 16606 16626 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal1 18308 13498 18308 13498 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal1 17434 18258 17434 18258 0 mem_bottom_track_25.DFFR_6_.Q
rlabel metal1 6900 13906 6900 13906 0 mem_bottom_track_25.DFFR_7_.Q
rlabel metal1 16974 18768 16974 18768 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal2 18768 6222 18768 6222 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal4 32292 17204 32292 17204 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal1 29946 2278 29946 2278 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal1 35374 2482 35374 2482 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal2 36662 2176 36662 2176 0 mem_bottom_track_33.DFFR_5_.Q
rlabel metal1 14122 7854 14122 7854 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal1 17066 3570 17066 3570 0 mem_bottom_track_9.DFFR_1_.Q
rlabel via3 18653 16660 18653 16660 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal1 24518 2346 24518 2346 0 mem_bottom_track_9.DFFR_3_.Q
rlabel via2 27462 2363 27462 2363 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal1 29210 2618 29210 2618 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal1 33442 4046 33442 4046 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal1 15134 19414 15134 19414 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 19734 7752 19734 7752 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 20240 2278 20240 2278 0 mem_left_track_1.DFFR_2_.Q
rlabel metal1 21896 2346 21896 2346 0 mem_left_track_1.DFFR_3_.Q
rlabel metal2 33350 15249 33350 15249 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 26726 15470 26726 15470 0 mem_left_track_1.DFFR_5_.Q
rlabel metal2 28520 15028 28520 15028 0 mem_left_track_1.DFFR_6_.Q
rlabel metal1 33626 20434 33626 20434 0 mem_left_track_1.DFFR_7_.Q
rlabel metal1 27830 19142 27830 19142 0 mem_left_track_17.DFFR_0_.D
rlabel metal2 29210 11220 29210 11220 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 32982 20009 32982 20009 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 34822 20502 34822 20502 0 mem_left_track_17.DFFR_2_.Q
rlabel metal1 32936 24786 32936 24786 0 mem_left_track_17.DFFR_3_.Q
rlabel metal1 31648 15470 31648 15470 0 mem_left_track_17.DFFR_4_.Q
rlabel metal1 32131 11730 32131 11730 0 mem_left_track_17.DFFR_5_.Q
rlabel metal1 31464 5542 31464 5542 0 mem_left_track_17.DFFR_6_.Q
rlabel metal2 26726 5304 26726 5304 0 mem_left_track_17.DFFR_7_.Q
rlabel metal2 7866 22780 7866 22780 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 26174 19465 26174 19465 0 mem_left_track_25.DFFR_1_.Q
rlabel via2 21850 3179 21850 3179 0 mem_left_track_25.DFFR_2_.Q
rlabel metal2 20930 21471 20930 21471 0 mem_left_track_25.DFFR_3_.Q
rlabel metal1 8694 13804 8694 13804 0 mem_left_track_25.DFFR_4_.Q
rlabel metal1 9200 4794 9200 4794 0 mem_left_track_25.DFFR_5_.Q
rlabel metal1 11362 5814 11362 5814 0 mem_left_track_25.DFFR_6_.Q
rlabel metal1 8602 17646 8602 17646 0 mem_left_track_25.DFFR_7_.Q
rlabel metal2 14536 17612 14536 17612 0 mem_left_track_33.DFFR_0_.Q
rlabel metal1 18124 6698 18124 6698 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 15088 29614 15088 29614 0 mem_left_track_33.DFFR_2_.Q
rlabel metal2 14168 20876 14168 20876 0 mem_left_track_33.DFFR_3_.Q
rlabel metal1 14260 20774 14260 20774 0 mem_left_track_33.DFFR_4_.Q
rlabel via3 22011 20740 22011 20740 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 2484 6290 2484 6290 0 mem_left_track_9.DFFR_1_.Q
rlabel metal1 2622 9588 2622 9588 0 mem_left_track_9.DFFR_2_.Q
rlabel metal1 2622 7888 2622 7888 0 mem_left_track_9.DFFR_3_.Q
rlabel metal1 11500 2550 11500 2550 0 mem_left_track_9.DFFR_4_.Q
rlabel metal2 17158 13401 17158 13401 0 mem_left_track_9.DFFR_5_.Q
rlabel metal2 23276 15300 23276 15300 0 mem_left_track_9.DFFR_6_.Q
rlabel metal1 14582 19346 14582 19346 0 mem_right_track_0.DFFR_0_.D
rlabel metal1 18262 13362 18262 13362 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 14996 13838 14996 13838 0 mem_right_track_0.DFFR_1_.Q
rlabel metal3 20677 13668 20677 13668 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 12742 18088 12742 18088 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 17296 13974 17296 13974 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 19504 14314 19504 14314 0 mem_right_track_0.DFFR_5_.Q
rlabel metal1 20608 14246 20608 14246 0 mem_right_track_0.DFFR_6_.Q
rlabel metal1 20792 22610 20792 22610 0 mem_right_track_0.DFFR_7_.Q
rlabel metal2 16146 9537 16146 9537 0 mem_right_track_16.DFFR_0_.D
rlabel metal1 32476 21522 32476 21522 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 12735 14790 12735 14790 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 14720 14926 14720 14926 0 mem_right_track_16.DFFR_2_.Q
rlabel metal1 33442 20910 33442 20910 0 mem_right_track_16.DFFR_3_.Q
rlabel metal1 29256 16626 29256 16626 0 mem_right_track_16.DFFR_4_.Q
rlabel metal1 28060 14450 28060 14450 0 mem_right_track_16.DFFR_5_.Q
rlabel metal1 30866 17102 30866 17102 0 mem_right_track_16.DFFR_6_.Q
rlabel metal1 32039 14994 32039 14994 0 mem_right_track_16.DFFR_7_.Q
rlabel metal1 21666 13192 21666 13192 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 23046 13362 23046 13362 0 mem_right_track_24.DFFR_1_.Q
rlabel via2 13202 8789 13202 8789 0 mem_right_track_24.DFFR_2_.Q
rlabel metal1 13524 20910 13524 20910 0 mem_right_track_24.DFFR_3_.Q
rlabel metal1 11178 7990 11178 7990 0 mem_right_track_24.DFFR_4_.Q
rlabel metal1 14766 8874 14766 8874 0 mem_right_track_24.DFFR_5_.Q
rlabel metal1 17434 19822 17434 19822 0 mem_right_track_24.DFFR_6_.Q
rlabel metal2 15640 15572 15640 15572 0 mem_right_track_24.DFFR_7_.Q
rlabel metal2 13110 18462 13110 18462 0 mem_right_track_32.DFFR_0_.Q
rlabel metal2 19642 21148 19642 21148 0 mem_right_track_32.DFFR_1_.Q
rlabel metal2 13616 18836 13616 18836 0 mem_right_track_32.DFFR_2_.Q
rlabel metal3 17595 16796 17595 16796 0 mem_right_track_32.DFFR_3_.Q
rlabel metal2 21574 15844 21574 15844 0 mem_right_track_32.DFFR_4_.Q
rlabel metal1 7452 17646 7452 17646 0 mem_right_track_8.DFFR_0_.Q
rlabel metal4 13524 16184 13524 16184 0 mem_right_track_8.DFFR_1_.Q
rlabel metal3 14559 16660 14559 16660 0 mem_right_track_8.DFFR_2_.Q
rlabel metal1 16790 3434 16790 3434 0 mem_right_track_8.DFFR_3_.Q
rlabel metal2 13478 6562 13478 6562 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 6348 9724 6348 9724 0 mem_right_track_8.DFFR_5_.Q
rlabel metal2 6026 6460 6026 6460 0 mem_right_track_8.DFFR_6_.Q
rlabel metal2 29210 5270 29210 5270 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 31372 16082 31372 16082 0 mem_top_track_0.DFFR_1_.Q
rlabel metal2 20286 3740 20286 3740 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 18814 18734 18814 18734 0 mem_top_track_0.DFFR_3_.Q
rlabel metal2 25990 5406 25990 5406 0 mem_top_track_0.DFFR_4_.Q
rlabel metal1 32384 4522 32384 4522 0 mem_top_track_0.DFFR_5_.Q
rlabel metal1 33672 4454 33672 4454 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 17250 2142 17250 2142 0 mem_top_track_0.DFFR_7_.Q
rlabel metal2 11546 4794 11546 4794 0 mem_top_track_16.DFFR_0_.D
rlabel metal2 20930 20383 20930 20383 0 mem_top_track_16.DFFR_0_.Q
rlabel metal3 13455 20740 13455 20740 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 34270 16524 34270 16524 0 mem_top_track_16.DFFR_2_.Q
rlabel metal3 16077 12308 16077 12308 0 mem_top_track_16.DFFR_3_.Q
rlabel metal1 22954 2482 22954 2482 0 mem_top_track_16.DFFR_4_.Q
rlabel metal2 23782 1938 23782 1938 0 mem_top_track_16.DFFR_5_.Q
rlabel via2 16698 2635 16698 2635 0 mem_top_track_16.DFFR_6_.Q
rlabel metal1 26404 4522 26404 4522 0 mem_top_track_16.DFFR_7_.Q
rlabel metal2 35650 10319 35650 10319 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 20470 12002 20470 12002 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 18906 20774 18906 20774 0 mem_top_track_24.DFFR_2_.Q
rlabel metal2 18814 15708 18814 15708 0 mem_top_track_24.DFFR_3_.Q
rlabel metal1 18492 13770 18492 13770 0 mem_top_track_24.DFFR_4_.Q
rlabel metal1 16100 11526 16100 11526 0 mem_top_track_24.DFFR_5_.Q
rlabel metal3 19849 16524 19849 16524 0 mem_top_track_24.DFFR_6_.Q
rlabel metal2 13248 13940 13248 13940 0 mem_top_track_24.DFFR_7_.Q
rlabel metal1 14674 29682 14674 29682 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 16146 28628 16146 28628 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 13708 9622 13708 9622 0 mem_top_track_32.DFFR_2_.Q
rlabel metal1 13202 18224 13202 18224 0 mem_top_track_32.DFFR_3_.Q
rlabel metal1 12489 18734 12489 18734 0 mem_top_track_32.DFFR_4_.Q
rlabel metal2 18906 2006 18906 2006 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 13478 17238 13478 17238 0 mem_top_track_8.DFFR_1_.Q
rlabel via2 2622 6749 2622 6749 0 mem_top_track_8.DFFR_2_.Q
rlabel metal1 7176 2482 7176 2482 0 mem_top_track_8.DFFR_3_.Q
rlabel metal3 5796 10132 5796 10132 0 mem_top_track_8.DFFR_4_.Q
rlabel metal1 4692 3094 4692 3094 0 mem_top_track_8.DFFR_5_.Q
rlabel metal2 4922 5644 4922 5644 0 mem_top_track_8.DFFR_6_.Q
rlabel metal1 27462 24676 27462 24676 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 14030 31790 14030 31790 0 mux_bottom_track_1.INVTX1_10_.out
rlabel metal2 15134 23392 15134 23392 0 mux_bottom_track_1.INVTX1_11_.out
rlabel via1 31786 16235 31786 16235 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 33718 6766 33718 6766 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal2 34914 18632 34914 18632 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 26036 19890 26036 19890 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 32384 22406 32384 22406 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal2 30590 24038 30590 24038 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal2 9982 22848 9982 22848 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal2 21850 27880 21850 27880 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal1 20746 25194 20746 25194 0 mux_bottom_track_1.INVTX1_9_.out
rlabel metal2 32062 23868 32062 23868 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 31786 25075 31786 25075 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 22034 24378 22034 24378 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 33074 23154 33074 23154 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 37398 35836 37398 35836 0 mux_bottom_track_1.out
rlabel metal2 28106 26010 28106 26010 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal2 10166 19176 10166 19176 0 mux_bottom_track_17.INVTX1_10_.out
rlabel metal1 14306 25194 14306 25194 0 mux_bottom_track_17.INVTX1_11_.out
rlabel metal2 23690 29546 23690 29546 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 28612 20230 28612 20230 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 13754 22542 13754 22542 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 33258 5270 33258 5270 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 13754 29478 13754 29478 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal1 22080 20842 22080 20842 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal2 7498 27948 7498 27948 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal2 15962 24412 15962 24412 0 mux_bottom_track_17.INVTX1_8_.out
rlabel metal1 14398 20264 14398 20264 0 mux_bottom_track_17.INVTX1_9_.out
rlabel metal2 20930 25874 20930 25874 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 16100 26894 16100 26894 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 18722 17850 18722 17850 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 26450 16932 26450 16932 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 36708 6426 36708 6426 0 mux_bottom_track_17.out
rlabel metal2 33166 22304 33166 22304 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 17066 27030 17066 27030 0 mux_bottom_track_25.INVTX1_10_.out
rlabel metal1 7544 31110 7544 31110 0 mux_bottom_track_25.INVTX1_11_.out
rlabel metal1 23414 19312 23414 19312 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal1 10994 23290 10994 23290 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal1 9200 31926 9200 31926 0 mux_bottom_track_25.INVTX1_3_.out
rlabel metal1 27554 27506 27554 27506 0 mux_bottom_track_25.INVTX1_4_.out
rlabel metal1 28750 25670 28750 25670 0 mux_bottom_track_25.INVTX1_5_.out
rlabel metal2 25806 24446 25806 24446 0 mux_bottom_track_25.INVTX1_6_.out
rlabel metal1 32614 12410 32614 12410 0 mux_bottom_track_25.INVTX1_7_.out
rlabel metal1 25576 27982 25576 27982 0 mux_bottom_track_25.INVTX1_8_.out
rlabel metal1 24610 26282 24610 26282 0 mux_bottom_track_25.INVTX1_9_.out
rlabel metal2 17802 20128 17802 20128 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 30774 17578 30774 17578 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 18354 17102 18354 17102 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 17986 15810 17986 15810 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 4002 12988 4002 12988 0 mux_bottom_track_25.out
rlabel metal1 17250 19278 17250 19278 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal1 17710 27948 17710 27948 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal2 15042 19550 15042 19550 0 mux_bottom_track_33.INVTX1_2_.out
rlabel metal1 15732 17714 15732 17714 0 mux_bottom_track_33.INVTX1_3_.out
rlabel metal2 33534 6579 33534 6579 0 mux_bottom_track_33.INVTX1_4_.out
rlabel metal1 30222 9452 30222 9452 0 mux_bottom_track_33.INVTX1_5_.out
rlabel metal1 15180 22066 15180 22066 0 mux_bottom_track_33.INVTX1_6_.out
rlabel metal1 17526 22066 17526 22066 0 mux_bottom_track_33.INVTX1_7_.out
rlabel metal1 18814 19754 18814 19754 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 32246 6188 32246 6188 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 29026 21352 29026 21352 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 28152 16490 28152 16490 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 38318 9452 38318 9452 0 mux_bottom_track_33.out
rlabel metal1 9476 15538 9476 15538 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal2 18814 19047 18814 19047 0 mux_bottom_track_9.INVTX1_10_.out
rlabel metal1 9292 13498 9292 13498 0 mux_bottom_track_9.INVTX1_11_.out
rlabel metal1 4784 5610 4784 5610 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal2 19642 9248 19642 9248 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 6532 12682 6532 12682 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal2 17066 6528 17066 6528 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal2 18814 3536 18814 3536 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal2 7590 8772 7590 8772 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal2 34638 6494 34638 6494 0 mux_bottom_track_9.INVTX1_7_.out
rlabel metal1 8464 16014 8464 16014 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal2 15686 16354 15686 16354 0 mux_bottom_track_9.INVTX1_9_.out
rlabel metal2 28106 4114 28106 4114 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 17250 6222 17250 6222 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 8694 15198 8694 15198 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 33994 5814 33994 5814 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 37950 9554 37950 9554 0 mux_bottom_track_9.out
rlabel metal1 10534 18190 10534 18190 0 mux_left_track_1.INVTX1_10_.out
rlabel metal2 3450 7786 3450 7786 0 mux_left_track_1.INVTX1_11_.out
rlabel metal1 28382 21930 28382 21930 0 mux_left_track_1.INVTX1_1_.out
rlabel metal2 26634 25704 26634 25704 0 mux_left_track_1.INVTX1_7_.out
rlabel metal1 14628 20366 14628 20366 0 mux_left_track_1.INVTX1_8_.out
rlabel metal2 11822 16813 11822 16813 0 mux_left_track_1.INVTX1_9_.out
rlabel metal1 32062 17578 32062 17578 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 27462 20094 27462 20094 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 15686 17017 15686 17017 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 32614 26384 32614 26384 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 33672 26554 33672 26554 0 mux_left_track_1.out
rlabel metal1 34730 18938 34730 18938 0 mux_left_track_17.INVTX1_10_.out
rlabel metal2 33718 25500 33718 25500 0 mux_left_track_17.INVTX1_11_.out
rlabel metal2 24058 21998 24058 21998 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 34868 8058 34868 8058 0 mux_left_track_17.INVTX1_7_.out
rlabel metal2 29118 30362 29118 30362 0 mux_left_track_17.INVTX1_8_.out
rlabel metal1 33120 20978 33120 20978 0 mux_left_track_17.INVTX1_9_.out
rlabel metal2 31786 18071 31786 18071 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 33166 19040 33166 19040 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 34362 25160 34362 25160 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 35052 15402 35052 15402 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 36156 9146 36156 9146 0 mux_left_track_17.out
rlabel metal2 25162 21216 25162 21216 0 mux_left_track_25.INVTX1_10_.out
rlabel via2 8970 4131 8970 4131 0 mux_left_track_25.INVTX1_11_.out
rlabel metal3 6785 6596 6785 6596 0 mux_left_track_25.INVTX1_2_.out
rlabel metal1 22264 20366 22264 20366 0 mux_left_track_25.INVTX1_7_.out
rlabel metal1 18538 20366 18538 20366 0 mux_left_track_25.INVTX1_8_.out
rlabel metal1 35006 3400 35006 3400 0 mux_left_track_25.INVTX1_9_.out
rlabel metal1 11316 16150 11316 16150 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 20930 19550 20930 19550 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 32614 3655 32614 3655 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 8648 19414 8648 19414 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 7590 19958 7590 19958 0 mux_left_track_25.out
rlabel metal2 14858 28832 14858 28832 0 mux_left_track_33.INVTX1_1_.out
rlabel metal1 11316 19754 11316 19754 0 mux_left_track_33.INVTX1_5_.out
rlabel metal1 20654 19924 20654 19924 0 mux_left_track_33.INVTX1_6_.out
rlabel metal1 13570 31926 13570 31926 0 mux_left_track_33.INVTX1_7_.out
rlabel metal1 14444 27846 14444 27846 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 15962 27098 15962 27098 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 14950 28832 14950 28832 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 18262 30294 18262 30294 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19366 36754 19366 36754 0 mux_left_track_33.out
rlabel metal1 6440 17102 6440 17102 0 mux_left_track_9.INVTX1_10_.out
rlabel metal2 4002 8194 4002 8194 0 mux_left_track_9.INVTX1_11_.out
rlabel metal1 5612 2618 5612 2618 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 5612 15402 5612 15402 0 mux_left_track_9.INVTX1_7_.out
rlabel metal1 23874 31110 23874 31110 0 mux_left_track_9.INVTX1_8_.out
rlabel metal1 4600 6222 4600 6222 0 mux_left_track_9.INVTX1_9_.out
rlabel metal1 6210 2482 6210 2482 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 15594 15028 15594 15028 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 21574 16490 21574 16490 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 36478 31314 36478 31314 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 37950 31314 37950 31314 0 mux_left_track_9.out
rlabel metal1 7452 33286 7452 33286 0 mux_right_track_0.INVTX1_4_.out
rlabel metal1 17802 21896 17802 21896 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 12420 30770 12420 30770 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 21344 24242 21344 24242 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 20378 34102 20378 34102 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 23828 35802 23828 35802 0 mux_right_track_0.out
rlabel metal1 30866 29206 30866 29206 0 mux_right_track_16.INVTX1_4_.out
rlabel metal1 28980 18938 28980 18938 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 31096 21046 31096 21046 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 17894 19397 17894 19397 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 34914 17680 34914 17680 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 35374 17646 35374 17646 0 mux_right_track_16.out
rlabel metal1 25714 32742 25714 32742 0 mux_right_track_24.INVTX1_4_.out
rlabel metal1 15870 21012 15870 21012 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 17066 24718 17066 24718 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 17756 20978 17756 20978 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 18446 20808 18446 20808 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 6854 28016 6854 28016 0 mux_right_track_24.out
rlabel metal1 14536 21590 14536 21590 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20102 18326 20102 18326 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 21206 21930 21206 21930 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 21390 17000 21390 17000 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 34684 17306 34684 17306 0 mux_right_track_32.out
rlabel metal1 5980 31790 5980 31790 0 mux_right_track_8.INVTX1_4_.out
rlabel metal2 15410 17085 15410 17085 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 35282 3519 35282 3519 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 7590 17272 7590 17272 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 7038 8670 7038 8670 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 5106 12614 5106 12614 0 mux_right_track_8.out
rlabel metal1 33764 3570 33764 3570 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 32430 12070 32430 12070 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 15226 20009 15226 20009 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 20148 19210 20148 19210 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 33074 5576 33074 5576 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 35834 9758 35834 9758 0 mux_top_track_0.out
rlabel metal2 13662 28526 13662 28526 0 mux_top_track_16.INVTX1_0_.out
rlabel metal1 14766 22542 14766 22542 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 31924 16490 31924 16490 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 17940 16762 17940 16762 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 33396 12274 33396 12274 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 34868 12818 34868 12818 0 mux_top_track_16.out
rlabel metal2 33810 22610 33810 22610 0 mux_top_track_24.INVTX1_0_.out
rlabel metal2 19918 21148 19918 21148 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 20102 19822 20102 19822 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 19274 26656 19274 26656 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 21022 20842 21022 20842 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 6210 28526 6210 28526 0 mux_top_track_24.out
rlabel metal1 10212 28730 10212 28730 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13754 25568 13754 25568 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15686 28424 15686 28424 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 12834 27438 12834 27438 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 10718 30260 10718 30260 0 mux_top_track_32.out
rlabel metal1 4922 8398 4922 8398 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 7544 10710 7544 10710 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 7682 14926 7682 14926 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 14582 15844 14582 15844 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 4968 5134 4968 5134 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 2162 8738 2162 8738 0 mux_top_track_8.out
rlabel metal2 6762 29546 6762 29546 0 net1
rlabel metal3 20539 13260 20539 13260 0 net10
rlabel metal2 16514 23307 16514 23307 0 net100
rlabel metal1 37950 23834 37950 23834 0 net101
rlabel metal1 38042 33422 38042 33422 0 net102
rlabel metal1 19780 36890 19780 36890 0 net103
rlabel metal1 23736 37094 23736 37094 0 net104
rlabel metal1 2300 14586 2300 14586 0 net105
rlabel metal1 36340 37230 36340 37230 0 net106
rlabel metal1 2024 36686 2024 36686 0 net107
rlabel metal1 1702 19346 1702 19346 0 net108
rlabel metal1 38088 31450 38088 31450 0 net109
rlabel via2 9154 13277 9154 13277 0 net11
rlabel metal1 20286 36856 20286 36856 0 net110
rlabel metal2 2346 36278 2346 36278 0 net111
rlabel metal1 32338 36686 32338 36686 0 net112
rlabel metal1 37766 6766 37766 6766 0 net113
rlabel metal2 3174 2074 3174 2074 0 net114
rlabel metal2 24058 37060 24058 37060 0 net115
rlabel metal1 11040 36754 11040 36754 0 net116
rlabel metal1 36708 24786 36708 24786 0 net117
rlabel metal2 6670 28662 6670 28662 0 net118
rlabel metal1 34270 23834 34270 23834 0 net119
rlabel metal2 8326 18564 8326 18564 0 net12
rlabel metal1 1610 22032 1610 22032 0 net120
rlabel metal1 37582 34918 37582 34918 0 net121
rlabel metal1 37996 14382 37996 14382 0 net122
rlabel metal1 4968 36754 4968 36754 0 net123
rlabel metal1 1380 5202 1380 5202 0 net124
rlabel metal3 4531 2516 4531 2516 0 net125
rlabel metal1 1748 23834 1748 23834 0 net126
rlabel metal1 1610 16014 1610 16014 0 net127
rlabel metal1 1610 11084 1610 11084 0 net128
rlabel metal1 36110 4114 36110 4114 0 net129
rlabel metal1 9982 36686 9982 36686 0 net13
rlabel metal2 35558 36652 35558 36652 0 net130
rlabel metal1 20240 9894 20240 9894 0 net131
rlabel metal1 37628 16082 37628 16082 0 net132
rlabel metal1 37950 8942 37950 8942 0 net133
rlabel metal1 37628 36142 37628 36142 0 net134
rlabel metal1 1610 35700 1610 35700 0 net135
rlabel metal2 22494 37060 22494 37060 0 net136
rlabel metal1 1610 7922 1610 7922 0 net137
rlabel metal1 27370 37230 27370 37230 0 net138
rlabel metal2 3082 4641 3082 4641 0 net139
rlabel metal1 17020 37298 17020 37298 0 net14
rlabel metal2 2438 6154 2438 6154 0 net140
rlabel metal1 37398 5202 37398 5202 0 net141
rlabel metal1 2530 36142 2530 36142 0 net142
rlabel metal2 38042 27812 38042 27812 0 net143
rlabel metal1 12282 37230 12282 37230 0 net144
rlabel metal1 24150 29614 24150 29614 0 net145
rlabel metal2 2346 2601 2346 2601 0 net146
rlabel metal2 38042 8908 38042 8908 0 net147
rlabel metal2 38042 22780 38042 22780 0 net148
rlabel metal1 13662 37230 13662 37230 0 net149
rlabel metal2 4002 36890 4002 36890 0 net15
rlabel metal1 37720 14586 37720 14586 0 net150
rlabel metal2 37306 7378 37306 7378 0 net151
rlabel metal1 2668 7174 2668 7174 0 net152
rlabel metal1 37720 5678 37720 5678 0 net153
rlabel metal1 35788 21862 35788 21862 0 net154
rlabel metal1 6624 23290 6624 23290 0 net155
rlabel metal2 6394 29172 6394 29172 0 net156
rlabel metal3 24104 20740 24104 20740 0 net157
rlabel metal2 2346 8364 2346 8364 0 net158
rlabel metal1 1518 4114 1518 4114 0 net159
rlabel metal1 2392 4794 2392 4794 0 net16
rlabel metal1 3128 33490 3128 33490 0 net160
rlabel metal1 17250 19176 17250 19176 0 net161
rlabel metal1 20976 37230 20976 37230 0 net162
rlabel metal1 17986 25262 17986 25262 0 net163
rlabel metal1 1702 11254 1702 11254 0 net164
rlabel metal2 1978 3553 1978 3553 0 net165
rlabel metal1 1564 6290 1564 6290 0 net166
rlabel metal1 18676 29818 18676 29818 0 net167
rlabel metal1 9522 6120 9522 6120 0 net168
rlabel metal1 25392 33830 25392 33830 0 net169
rlabel metal1 23782 37298 23782 37298 0 net17
rlabel metal1 36386 12614 36386 12614 0 net170
rlabel metal1 1840 5678 1840 5678 0 net171
rlabel metal1 33764 5746 33764 5746 0 net172
rlabel metal1 4370 9044 4370 9044 0 net173
rlabel metal2 32614 10914 32614 10914 0 net174
rlabel metal2 12742 27200 12742 27200 0 net175
rlabel metal2 19366 32606 19366 32606 0 net176
rlabel metal2 5842 11424 5842 11424 0 net177
rlabel metal1 33442 19448 33442 19448 0 net178
rlabel metal2 9430 24480 9430 24480 0 net179
rlabel metal1 32338 9588 32338 9588 0 net18
rlabel metal1 29302 25976 29302 25976 0 net180
rlabel metal1 34822 6834 34822 6834 0 net181
rlabel metal1 32154 6834 32154 6834 0 net182
rlabel metal1 6302 16014 6302 16014 0 net183
rlabel metal2 30038 24480 30038 24480 0 net184
rlabel metal2 28014 21420 28014 21420 0 net185
rlabel metal1 34132 7514 34132 7514 0 net186
rlabel metal2 8142 17714 8142 17714 0 net187
rlabel metal1 13064 29070 13064 29070 0 net188
rlabel metal1 15824 21658 15824 21658 0 net189
rlabel metal2 33810 23868 33810 23868 0 net19
rlabel metal2 28750 20655 28750 20655 0 net190
rlabel metal2 14858 31008 14858 31008 0 net191
rlabel metal2 37030 10642 37030 10642 0 net2
rlabel metal1 1334 4794 1334 4794 0 net20
rlabel metal1 18814 37298 18814 37298 0 net21
rlabel metal1 10350 37094 10350 37094 0 net22
rlabel metal2 38134 16796 38134 16796 0 net23
rlabel metal2 2254 3315 2254 3315 0 net24
rlabel metal1 36478 19312 36478 19312 0 net25
rlabel metal2 38272 28084 38272 28084 0 net26
rlabel metal1 29854 5780 29854 5780 0 net27
rlabel metal1 1886 37196 1886 37196 0 net28
rlabel metal1 37996 23698 37996 23698 0 net29
rlabel metal1 6486 21998 6486 21998 0 net3
rlabel metal2 2070 23426 2070 23426 0 net30
rlabel metal1 33534 23630 33534 23630 0 net31
rlabel metal3 19113 21148 19113 21148 0 net32
rlabel metal2 37674 30974 37674 30974 0 net33
rlabel metal2 3266 10540 3266 10540 0 net34
rlabel metal2 1886 5865 1886 5865 0 net35
rlabel metal1 1748 24582 1748 24582 0 net36
rlabel metal2 5382 36822 5382 36822 0 net37
rlabel metal1 20470 36788 20470 36788 0 net38
rlabel metal2 1886 30226 1886 30226 0 net39
rlabel metal2 34178 9860 34178 9860 0 net4
rlabel metal2 23598 36550 23598 36550 0 net40
rlabel metal2 6946 10132 6946 10132 0 net41
rlabel metal2 38226 12665 38226 12665 0 net42
rlabel metal1 10672 37230 10672 37230 0 net43
rlabel metal2 37490 25299 37490 25299 0 net44
rlabel metal3 15985 3876 15985 3876 0 net45
rlabel metal1 26910 6664 26910 6664 0 net46
rlabel metal2 33166 30532 33166 30532 0 net47
rlabel metal1 2530 11696 2530 11696 0 net48
rlabel metal1 2070 36074 2070 36074 0 net49
rlabel metal1 26956 5270 26956 5270 0 net5
rlabel metal1 9292 36550 9292 36550 0 net50
rlabel metal1 36892 18734 36892 18734 0 net51
rlabel metal1 36708 19890 36708 19890 0 net52
rlabel metal1 5750 7378 5750 7378 0 net53
rlabel metal2 37306 16779 37306 16779 0 net54
rlabel metal1 37444 9894 37444 9894 0 net55
rlabel metal1 28014 31314 28014 31314 0 net56
rlabel metal1 20194 29614 20194 29614 0 net57
rlabel metal2 5474 18258 5474 18258 0 net58
rlabel metal1 1932 12886 1932 12886 0 net59
rlabel metal1 36018 37128 36018 37128 0 net6
rlabel metal1 23230 37162 23230 37162 0 net60
rlabel metal1 14766 6120 14766 6120 0 net61
rlabel metal1 35788 21998 35788 21998 0 net62
rlabel metal2 37766 28832 37766 28832 0 net63
rlabel metal1 22678 36720 22678 36720 0 net64
rlabel metal2 3266 7004 3266 7004 0 net65
rlabel metal2 34454 25466 34454 25466 0 net66
rlabel metal1 31878 6290 31878 6290 0 net67
rlabel metal2 21482 7905 21482 7905 0 net68
rlabel metal2 5566 23562 5566 23562 0 net69
rlabel metal1 36202 24242 36202 24242 0 net7
rlabel metal1 33442 26962 33442 26962 0 net70
rlabel metal2 966 12920 966 12920 0 net71
rlabel metal1 1978 9010 1978 9010 0 net72
rlabel metal2 1886 14603 1886 14603 0 net73
rlabel metal2 31786 31042 31786 31042 0 net74
rlabel metal2 38134 23358 38134 23358 0 net75
rlabel metal1 37720 2482 37720 2482 0 net76
rlabel metal1 6762 19890 6762 19890 0 net77
rlabel metal2 37582 15538 37582 15538 0 net78
rlabel metal2 8326 27574 8326 27574 0 net79
rlabel metal1 16974 36550 16974 36550 0 net8
rlabel metal2 2990 8806 2990 8806 0 net80
rlabel metal2 36846 36414 36846 36414 0 net81
rlabel metal1 34362 25874 34362 25874 0 net82
rlabel metal1 3082 6290 3082 6290 0 net83
rlabel metal1 13685 10438 13685 10438 0 net84
rlabel metal2 3910 8398 3910 8398 0 net85
rlabel metal1 37720 26758 37720 26758 0 net86
rlabel metal1 29854 32402 29854 32402 0 net87
rlabel metal2 26082 35020 26082 35020 0 net88
rlabel metal1 4462 36006 4462 36006 0 net89
rlabel metal1 34914 20842 34914 20842 0 net9
rlabel metal1 6118 31858 6118 31858 0 net90
rlabel metal2 29854 7667 29854 7667 0 net91
rlabel metal1 3634 8398 3634 8398 0 net92
rlabel metal2 2622 32198 2622 32198 0 net93
rlabel metal1 38088 19482 38088 19482 0 net94
rlabel metal1 4278 36822 4278 36822 0 net95
rlabel metal2 36754 34646 36754 34646 0 net96
rlabel metal2 5106 36924 5106 36924 0 net97
rlabel metal1 29900 3502 29900 3502 0 net98
rlabel metal2 6854 20740 6854 20740 0 net99
rlabel metal2 38318 26775 38318 26775 0 pReset
rlabel metal2 21942 5814 21942 5814 0 prog_clk
rlabel metal1 29118 37230 29118 37230 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal1 27922 37230 27922 37230 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 3128 36142 3128 36142 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 7268 36142 7268 36142 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 27738 1761 27738 1761 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal3 1234 10268 1234 10268 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 1234 34068 1234 34068 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 38318 19227 38318 19227 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
