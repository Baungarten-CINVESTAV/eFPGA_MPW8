magic
tech sky130A
magscale 1 2
timestamp 1672417828
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 20626 39200 20682 39800
rect 22558 39200 22614 39800
rect 23846 39200 23902 39800
rect 25778 39200 25834 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 13542 200 13598 800
rect 15474 200 15530 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
rect 38658 200 38714 800
<< obsm2 >>
rect 18 39144 606 39545
rect 774 39144 1894 39545
rect 2062 39144 3826 39545
rect 3994 39144 5114 39545
rect 5282 39144 7046 39545
rect 7214 39144 8334 39545
rect 8502 39144 10266 39545
rect 10434 39144 11554 39545
rect 11722 39144 12842 39545
rect 13010 39144 14774 39545
rect 14942 39144 16062 39545
rect 16230 39144 17994 39545
rect 18162 39144 19282 39545
rect 19450 39144 20570 39545
rect 20738 39144 22502 39545
rect 22670 39144 23790 39545
rect 23958 39144 25722 39545
rect 25890 39144 27010 39545
rect 27178 39144 28942 39545
rect 29110 39144 30230 39545
rect 30398 39144 31518 39545
rect 31686 39144 33450 39545
rect 33618 39144 34738 39545
rect 34906 39144 36670 39545
rect 36838 39144 37958 39545
rect 38126 39144 39246 39545
rect 18 856 39356 39144
rect 130 144 1250 856
rect 1418 144 2538 856
rect 2706 144 4470 856
rect 4638 144 5758 856
rect 5926 144 7690 856
rect 7858 144 8978 856
rect 9146 144 10266 856
rect 10434 144 12198 856
rect 12366 144 13486 856
rect 13654 144 15418 856
rect 15586 144 16706 856
rect 16874 144 18638 856
rect 18806 144 19926 856
rect 20094 144 21214 856
rect 21382 144 23146 856
rect 23314 144 24434 856
rect 24602 144 26366 856
rect 26534 144 27654 856
rect 27822 144 28942 856
rect 29110 144 30874 856
rect 31042 144 32162 856
rect 32330 144 34094 856
rect 34262 144 35382 856
rect 35550 144 37314 856
rect 37482 144 38602 856
rect 38770 144 39356 856
rect 18 31 39356 144
<< metal3 >>
rect 200 39448 800 39568
rect 39200 38088 39800 38208
rect 200 37408 800 37528
rect 39200 36728 39800 36848
rect 200 36048 800 36168
rect 39200 34688 39800 34808
rect 200 34008 800 34128
rect 39200 33328 39800 33448
rect 200 32648 800 32768
rect 39200 31288 39800 31408
rect 200 30608 800 30728
rect 39200 29928 39800 30048
rect 200 29248 800 29368
rect 39200 28568 39800 28688
rect 200 27888 800 28008
rect 39200 26528 39800 26648
rect 200 25848 800 25968
rect 39200 25168 39800 25288
rect 200 24488 800 24608
rect 39200 23128 39800 23248
rect 200 22448 800 22568
rect 39200 21768 39800 21888
rect 200 21088 800 21208
rect 200 19728 800 19848
rect 39200 19728 39800 19848
rect 39200 18368 39800 18488
rect 200 17688 800 17808
rect 39200 17008 39800 17128
rect 200 16328 800 16448
rect 39200 14968 39800 15088
rect 200 14288 800 14408
rect 39200 13608 39800 13728
rect 200 12928 800 13048
rect 39200 11568 39800 11688
rect 200 10888 800 11008
rect 39200 10208 39800 10328
rect 200 9528 800 9648
rect 39200 8848 39800 8968
rect 200 8168 800 8288
rect 39200 6808 39800 6928
rect 200 6128 800 6248
rect 39200 5448 39800 5568
rect 200 4768 800 4888
rect 39200 3408 39800 3528
rect 200 2728 800 2848
rect 39200 2048 39800 2168
rect 200 1368 800 1488
rect 39200 8 39800 128
<< obsm3 >>
rect 13 39368 120 39541
rect 880 39368 39200 39541
rect 13 38288 39200 39368
rect 13 38008 39120 38288
rect 13 37608 39200 38008
rect 13 37328 120 37608
rect 880 37328 39200 37608
rect 13 36928 39200 37328
rect 13 36648 39120 36928
rect 13 36248 39200 36648
rect 13 35968 120 36248
rect 880 35968 39200 36248
rect 13 34888 39200 35968
rect 13 34608 39120 34888
rect 13 34208 39200 34608
rect 13 33928 120 34208
rect 880 33928 39200 34208
rect 13 33528 39200 33928
rect 13 33248 39120 33528
rect 13 32848 39200 33248
rect 13 32568 120 32848
rect 880 32568 39200 32848
rect 13 31488 39200 32568
rect 13 31208 39120 31488
rect 13 30808 39200 31208
rect 13 30528 120 30808
rect 880 30528 39200 30808
rect 13 30128 39200 30528
rect 13 29848 39120 30128
rect 13 29448 39200 29848
rect 13 29168 120 29448
rect 880 29168 39200 29448
rect 13 28768 39200 29168
rect 13 28488 39120 28768
rect 13 28088 39200 28488
rect 13 27808 120 28088
rect 880 27808 39200 28088
rect 13 26728 39200 27808
rect 13 26448 39120 26728
rect 13 26048 39200 26448
rect 13 25768 120 26048
rect 880 25768 39200 26048
rect 13 25368 39200 25768
rect 13 25088 39120 25368
rect 13 24688 39200 25088
rect 13 24408 120 24688
rect 880 24408 39200 24688
rect 13 23328 39200 24408
rect 13 23048 39120 23328
rect 13 22648 39200 23048
rect 13 22368 120 22648
rect 880 22368 39200 22648
rect 13 21968 39200 22368
rect 13 21688 39120 21968
rect 13 21288 39200 21688
rect 13 21008 120 21288
rect 880 21008 39200 21288
rect 13 19928 39200 21008
rect 13 19648 120 19928
rect 880 19648 39120 19928
rect 13 18568 39200 19648
rect 13 18288 39120 18568
rect 13 17888 39200 18288
rect 13 17778 120 17888
rect 13 17776 200 17778
rect 13 17720 120 17776
rect 13 17718 200 17720
rect 13 17608 120 17718
rect 880 17608 39200 17888
rect 13 17208 39200 17608
rect 13 16928 39120 17208
rect 13 16528 39200 16928
rect 13 16248 120 16528
rect 880 16248 39200 16528
rect 13 15168 39200 16248
rect 13 14888 39120 15168
rect 13 14488 39200 14888
rect 13 14208 120 14488
rect 880 14208 39200 14488
rect 13 13808 39200 14208
rect 13 13528 39120 13808
rect 13 13128 39200 13528
rect 13 12848 120 13128
rect 880 12848 39200 13128
rect 13 11768 39200 12848
rect 13 11488 39120 11768
rect 13 11088 39200 11488
rect 13 10808 120 11088
rect 880 10808 39200 11088
rect 13 10408 39200 10808
rect 13 10128 39120 10408
rect 13 9728 39200 10128
rect 13 9448 120 9728
rect 880 9448 39200 9728
rect 13 9048 39200 9448
rect 13 8768 39120 9048
rect 13 8368 39200 8768
rect 13 8088 120 8368
rect 880 8088 39200 8368
rect 13 7008 39200 8088
rect 13 6728 39120 7008
rect 13 6328 39200 6728
rect 13 6048 120 6328
rect 880 6048 39200 6328
rect 13 5648 39200 6048
rect 13 5368 39120 5648
rect 13 4968 39200 5368
rect 13 4688 120 4968
rect 880 4688 39200 4968
rect 13 3608 39200 4688
rect 13 3328 39120 3608
rect 13 2928 39200 3328
rect 13 2648 120 2928
rect 880 2648 39200 2928
rect 13 2248 39200 2648
rect 13 1968 39120 2248
rect 13 1568 39200 1968
rect 13 1288 120 1568
rect 880 1288 39200 1568
rect 13 208 39200 1288
rect 13 35 39120 208
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 1899 3979 4128 36685
rect 4608 3979 15949 36685
<< labels >>
rlabel metal2 s 7102 39200 7158 39800 6 ccff_head
port 1 nsew signal input
rlabel metal2 s 3882 39200 3938 39800 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 200 27888 800 28008 6 chanx_left_in[0]
port 3 nsew signal input
rlabel metal3 s 39200 11568 39800 11688 6 chanx_left_in[10]
port 4 nsew signal input
rlabel metal3 s 39200 25168 39800 25288 6 chanx_left_in[11]
port 5 nsew signal input
rlabel metal2 s 22558 39200 22614 39800 6 chanx_left_in[12]
port 6 nsew signal input
rlabel metal2 s 10322 200 10378 800 6 chanx_left_in[13]
port 7 nsew signal input
rlabel metal2 s 15474 200 15530 800 6 chanx_left_in[14]
port 8 nsew signal input
rlabel metal2 s 32218 200 32274 800 6 chanx_left_in[15]
port 9 nsew signal input
rlabel metal3 s 200 1368 800 1488 6 chanx_left_in[16]
port 10 nsew signal input
rlabel metal3 s 39200 31288 39800 31408 6 chanx_left_in[17]
port 11 nsew signal input
rlabel metal2 s 4526 200 4582 800 6 chanx_left_in[18]
port 12 nsew signal input
rlabel metal2 s 34150 200 34206 800 6 chanx_left_in[1]
port 13 nsew signal input
rlabel metal3 s 200 32648 800 32768 6 chanx_left_in[2]
port 14 nsew signal input
rlabel metal2 s 33506 39200 33562 39800 6 chanx_left_in[3]
port 15 nsew signal input
rlabel metal3 s 39200 19728 39800 19848 6 chanx_left_in[4]
port 16 nsew signal input
rlabel metal2 s 11610 39200 11666 39800 6 chanx_left_in[5]
port 17 nsew signal input
rlabel metal3 s 200 37408 800 37528 6 chanx_left_in[6]
port 18 nsew signal input
rlabel metal3 s 200 25848 800 25968 6 chanx_left_in[7]
port 19 nsew signal input
rlabel metal2 s 38658 200 38714 800 6 chanx_left_in[8]
port 20 nsew signal input
rlabel metal3 s 200 17688 800 17808 6 chanx_left_in[9]
port 21 nsew signal input
rlabel metal3 s 39200 34688 39800 34808 6 chanx_left_out[0]
port 22 nsew signal output
rlabel metal3 s 39200 5448 39800 5568 6 chanx_left_out[10]
port 23 nsew signal output
rlabel metal2 s 25778 39200 25834 39800 6 chanx_left_out[11]
port 24 nsew signal output
rlabel metal3 s 200 21088 800 21208 6 chanx_left_out[12]
port 25 nsew signal output
rlabel metal2 s 14830 39200 14886 39800 6 chanx_left_out[13]
port 26 nsew signal output
rlabel metal2 s 16118 39200 16174 39800 6 chanx_left_out[14]
port 27 nsew signal output
rlabel metal2 s 28998 39200 29054 39800 6 chanx_left_out[15]
port 28 nsew signal output
rlabel metal3 s 200 29248 800 29368 6 chanx_left_out[16]
port 29 nsew signal output
rlabel metal3 s 39200 38088 39800 38208 6 chanx_left_out[17]
port 30 nsew signal output
rlabel metal3 s 39200 33328 39800 33448 6 chanx_left_out[18]
port 31 nsew signal output
rlabel metal3 s 39200 36728 39800 36848 6 chanx_left_out[1]
port 32 nsew signal output
rlabel metal3 s 39200 8848 39800 8968 6 chanx_left_out[2]
port 33 nsew signal output
rlabel metal2 s 23846 39200 23902 39800 6 chanx_left_out[3]
port 34 nsew signal output
rlabel metal2 s 18050 39200 18106 39800 6 chanx_left_out[4]
port 35 nsew signal output
rlabel metal3 s 200 4768 800 4888 6 chanx_left_out[5]
port 36 nsew signal output
rlabel metal3 s 200 39448 800 39568 6 chanx_left_out[6]
port 37 nsew signal output
rlabel metal2 s 9034 200 9090 800 6 chanx_left_out[7]
port 38 nsew signal output
rlabel metal3 s 39200 28568 39800 28688 6 chanx_left_out[8]
port 39 nsew signal output
rlabel metal2 s 37370 200 37426 800 6 chanx_left_out[9]
port 40 nsew signal output
rlabel metal3 s 39200 14968 39800 15088 6 chany_top_in[0]
port 41 nsew signal input
rlabel metal2 s 20626 39200 20682 39800 6 chany_top_in[10]
port 42 nsew signal input
rlabel metal2 s 12898 39200 12954 39800 6 chany_top_in[11]
port 43 nsew signal input
rlabel metal3 s 39200 8 39800 128 6 chany_top_in[12]
port 44 nsew signal input
rlabel metal3 s 39200 29928 39800 30048 6 chany_top_in[13]
port 45 nsew signal input
rlabel metal2 s 38014 39200 38070 39800 6 chany_top_in[14]
port 46 nsew signal input
rlabel metal3 s 200 6128 800 6248 6 chany_top_in[15]
port 47 nsew signal input
rlabel metal2 s 13542 200 13598 800 6 chany_top_in[16]
port 48 nsew signal input
rlabel metal3 s 39200 6808 39800 6928 6 chany_top_in[17]
port 49 nsew signal input
rlabel metal3 s 200 22448 800 22568 6 chany_top_in[18]
port 50 nsew signal input
rlabel metal3 s 200 2728 800 2848 6 chany_top_in[1]
port 51 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 chany_top_in[2]
port 52 nsew signal input
rlabel metal2 s 10322 39200 10378 39800 6 chany_top_in[3]
port 53 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 chany_top_in[4]
port 54 nsew signal input
rlabel metal2 s 34794 39200 34850 39800 6 chany_top_in[5]
port 55 nsew signal input
rlabel metal2 s 24490 200 24546 800 6 chany_top_in[6]
port 56 nsew signal input
rlabel metal2 s 2594 200 2650 800 6 chany_top_in[7]
port 57 nsew signal input
rlabel metal3 s 200 19728 800 19848 6 chany_top_in[8]
port 58 nsew signal input
rlabel metal2 s 35438 200 35494 800 6 chany_top_in[9]
port 59 nsew signal input
rlabel metal3 s 39200 17008 39800 17128 6 chany_top_out[0]
port 60 nsew signal output
rlabel metal3 s 39200 10208 39800 10328 6 chany_top_out[10]
port 61 nsew signal output
rlabel metal2 s 27710 200 27766 800 6 chany_top_out[11]
port 62 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 chany_top_out[12]
port 63 nsew signal output
rlabel metal3 s 39200 2048 39800 2168 6 chany_top_out[13]
port 64 nsew signal output
rlabel metal2 s 5170 39200 5226 39800 6 chany_top_out[14]
port 65 nsew signal output
rlabel metal3 s 39200 13608 39800 13728 6 chany_top_out[15]
port 66 nsew signal output
rlabel metal3 s 200 16328 800 16448 6 chany_top_out[16]
port 67 nsew signal output
rlabel metal2 s 30930 200 30986 800 6 chany_top_out[17]
port 68 nsew signal output
rlabel metal3 s 39200 26528 39800 26648 6 chany_top_out[18]
port 69 nsew signal output
rlabel metal2 s 18694 200 18750 800 6 chany_top_out[1]
port 70 nsew signal output
rlabel metal3 s 200 24488 800 24608 6 chany_top_out[2]
port 71 nsew signal output
rlabel metal2 s 19982 200 20038 800 6 chany_top_out[3]
port 72 nsew signal output
rlabel metal2 s 18 200 74 800 6 chany_top_out[4]
port 73 nsew signal output
rlabel metal2 s 23202 200 23258 800 6 chany_top_out[5]
port 74 nsew signal output
rlabel metal3 s 200 8168 800 8288 6 chany_top_out[6]
port 75 nsew signal output
rlabel metal2 s 19338 39200 19394 39800 6 chany_top_out[7]
port 76 nsew signal output
rlabel metal3 s 200 12928 800 13048 6 chany_top_out[8]
port 77 nsew signal output
rlabel metal2 s 662 39200 718 39800 6 chany_top_out[9]
port 78 nsew signal output
rlabel metal2 s 5814 200 5870 800 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 79 nsew signal input
rlabel metal2 s 1306 200 1362 800 6 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 80 nsew signal input
rlabel metal2 s 36726 39200 36782 39800 6 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 81 nsew signal input
rlabel metal2 s 27066 39200 27122 39800 6 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 82 nsew signal input
rlabel metal2 s 16762 200 16818 800 6 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_
port 83 nsew signal input
rlabel metal2 s 39302 39200 39358 39800 6 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_
port 84 nsew signal input
rlabel metal3 s 39200 3408 39800 3528 6 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_
port 85 nsew signal input
rlabel metal3 s 200 9528 800 9648 6 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_
port 86 nsew signal input
rlabel metal3 s 39200 21768 39800 21888 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 87 nsew signal input
rlabel metal2 s 7746 200 7802 800 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 88 nsew signal input
rlabel metal2 s 12254 200 12310 800 6 pReset
port 89 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 prog_clk
port 90 nsew signal input
rlabel metal3 s 39200 23128 39800 23248 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 91 nsew signal input
rlabel metal2 s 21270 200 21326 800 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 92 nsew signal input
rlabel metal2 s 31574 39200 31630 39800 6 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 93 nsew signal input
rlabel metal2 s 30286 39200 30342 39800 6 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 94 nsew signal input
rlabel metal2 s 1950 39200 2006 39800 6 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 95 nsew signal input
rlabel metal2 s 8390 39200 8446 39800 6 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 96 nsew signal input
rlabel metal2 s 26422 200 26478 800 6 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 97 nsew signal input
rlabel metal3 s 200 10888 800 11008 6 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 98 nsew signal input
rlabel metal3 s 200 36048 800 36168 6 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 99 nsew signal input
rlabel metal3 s 39200 18368 39800 18488 6 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 100 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 101 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 101 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 102 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2154554
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/sb_4__0_/runs/22_12_30_10_29/results/signoff/sb_4__0_.magic.gds
string GDS_START 138996
<< end >>

