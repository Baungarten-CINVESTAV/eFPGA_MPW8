magic
tech sky130A
magscale 1 2
timestamp 1672416474
<< viali >>
rect 2881 37417 2915 37451
rect 9505 37417 9539 37451
rect 16221 37417 16255 37451
rect 21373 37417 21407 37451
rect 2329 37349 2363 37383
rect 22293 37349 22327 37383
rect 5549 37281 5583 37315
rect 6745 37281 6779 37315
rect 7205 37281 7239 37315
rect 11161 37281 11195 37315
rect 11713 37281 11747 37315
rect 13737 37281 13771 37315
rect 17509 37281 17543 37315
rect 18245 37281 18279 37315
rect 22753 37281 22787 37315
rect 23489 37281 23523 37315
rect 24869 37281 24903 37315
rect 35081 37281 35115 37315
rect 35541 37281 35575 37315
rect 2145 37213 2179 37247
rect 3065 37213 3099 37247
rect 3985 37213 4019 37247
rect 4813 37213 4847 37247
rect 5365 37213 5399 37247
rect 7481 37213 7515 37247
rect 8585 37213 8619 37247
rect 9229 37213 9263 37247
rect 10885 37213 10919 37247
rect 12541 37213 12575 37247
rect 13001 37213 13035 37247
rect 14381 37213 14415 37247
rect 16865 37213 16899 37247
rect 17693 37213 17727 37247
rect 19441 37213 19475 37247
rect 22109 37213 22143 37247
rect 22937 37213 22971 37247
rect 24685 37213 24719 37247
rect 27169 37213 27203 37247
rect 28733 37213 28767 37247
rect 29745 37213 29779 37247
rect 32321 37213 32355 37247
rect 33885 37213 33919 37247
rect 35817 37213 35851 37247
rect 4169 37077 4203 37111
rect 12357 37077 12391 37111
rect 14473 37077 14507 37111
rect 17049 37077 17083 37111
rect 19625 37077 19659 37111
rect 27353 37077 27387 37111
rect 28549 37077 28583 37111
rect 29929 37077 29963 37111
rect 32505 37077 32539 37111
rect 33701 37077 33735 37111
rect 1685 36873 1719 36907
rect 2329 36873 2363 36907
rect 4077 36873 4111 36907
rect 18889 36873 18923 36907
rect 24501 36873 24535 36907
rect 35081 36873 35115 36907
rect 36277 36873 36311 36907
rect 1869 36737 1903 36771
rect 4261 36737 4295 36771
rect 17601 36737 17635 36771
rect 18705 36737 18739 36771
rect 22569 36737 22603 36771
rect 23213 36737 23247 36771
rect 23857 36737 23891 36771
rect 34897 36737 34931 36771
rect 36093 36737 36127 36771
rect 17785 36601 17819 36635
rect 22753 36601 22787 36635
rect 23397 36601 23431 36635
rect 28825 36533 28859 36567
rect 33977 36533 34011 36567
rect 2237 36329 2271 36363
rect 36277 36329 36311 36363
rect 1593 36125 1627 36159
rect 36093 36125 36127 36159
rect 1777 35989 1811 36023
rect 36093 35649 36127 35683
rect 36277 35445 36311 35479
rect 36185 35241 36219 35275
rect 1869 35037 1903 35071
rect 36001 35037 36035 35071
rect 1685 34901 1719 34935
rect 35449 34901 35483 34935
rect 36093 33473 36127 33507
rect 36277 33337 36311 33371
rect 35541 33269 35575 33303
rect 1685 32793 1719 32827
rect 1777 32725 1811 32759
rect 1685 32521 1719 32555
rect 3985 31977 4019 32011
rect 36093 31841 36127 31875
rect 1869 31773 1903 31807
rect 4169 31773 4203 31807
rect 4629 31773 4663 31807
rect 36369 31773 36403 31807
rect 1685 31637 1719 31671
rect 1961 31433 1995 31467
rect 23581 31433 23615 31467
rect 27629 31433 27663 31467
rect 36369 31365 36403 31399
rect 2053 31297 2087 31331
rect 2513 31297 2547 31331
rect 19809 31297 19843 31331
rect 22937 31297 22971 31331
rect 27445 31297 27479 31331
rect 28089 31297 28123 31331
rect 19901 31093 19935 31127
rect 23029 31093 23063 31127
rect 1777 30889 1811 30923
rect 1961 30685 1995 30719
rect 36093 30209 36127 30243
rect 35633 30005 35667 30039
rect 36277 30005 36311 30039
rect 6009 29801 6043 29835
rect 1869 29597 1903 29631
rect 6101 29597 6135 29631
rect 6561 29597 6595 29631
rect 11989 29597 12023 29631
rect 1685 29461 1719 29495
rect 12081 29461 12115 29495
rect 35633 28033 35667 28067
rect 36277 28033 36311 28067
rect 36185 27829 36219 27863
rect 1869 27421 1903 27455
rect 1685 27285 1719 27319
rect 26801 26537 26835 26571
rect 36277 26469 36311 26503
rect 26617 26333 26651 26367
rect 36093 26333 36127 26367
rect 27353 26265 27387 26299
rect 1593 25245 1627 25279
rect 1869 25245 1903 25279
rect 1593 24905 1627 24939
rect 1593 24157 1627 24191
rect 1869 24157 1903 24191
rect 36093 24157 36127 24191
rect 36369 24157 36403 24191
rect 1593 23817 1627 23851
rect 7297 23817 7331 23851
rect 36369 23817 36403 23851
rect 6745 23681 6779 23715
rect 12265 23681 12299 23715
rect 12081 23545 12115 23579
rect 6561 23477 6595 23511
rect 12725 23477 12759 23511
rect 4721 23273 4755 23307
rect 4905 23069 4939 23103
rect 5457 22933 5491 22967
rect 36093 22593 36127 22627
rect 36277 22457 36311 22491
rect 1593 21981 1627 22015
rect 1777 21845 1811 21879
rect 1593 21641 1627 21675
rect 18981 21505 19015 21539
rect 18889 21301 18923 21335
rect 19625 21301 19659 21335
rect 35633 21097 35667 21131
rect 8401 20893 8435 20927
rect 9137 20893 9171 20927
rect 9781 20893 9815 20927
rect 35449 20893 35483 20927
rect 36093 20893 36127 20927
rect 8493 20825 8527 20859
rect 9229 20757 9263 20791
rect 36277 20757 36311 20791
rect 35725 20213 35759 20247
rect 29929 20009 29963 20043
rect 1593 19805 1627 19839
rect 1869 19805 1903 19839
rect 29745 19805 29779 19839
rect 30389 19805 30423 19839
rect 1593 19465 1627 19499
rect 34897 19465 34931 19499
rect 34713 19329 34747 19363
rect 35357 19329 35391 19363
rect 31033 18921 31067 18955
rect 30941 18717 30975 18751
rect 36093 18717 36127 18751
rect 1685 18649 1719 18683
rect 1869 18649 1903 18683
rect 23581 18581 23615 18615
rect 36277 18581 36311 18615
rect 1593 18377 1627 18411
rect 24593 18377 24627 18411
rect 26157 18241 26191 18275
rect 27353 18241 27387 18275
rect 22845 18173 22879 18207
rect 25973 18105 26007 18139
rect 22109 18037 22143 18071
rect 23305 18037 23339 18071
rect 24041 18037 24075 18071
rect 25053 18037 25087 18071
rect 27261 18037 27295 18071
rect 21373 17833 21407 17867
rect 21925 17833 21959 17867
rect 33241 17833 33275 17867
rect 22845 17697 22879 17731
rect 23121 17697 23155 17731
rect 23857 17629 23891 17663
rect 24685 17629 24719 17663
rect 25513 17629 25547 17663
rect 25973 17629 26007 17663
rect 33149 17629 33183 17663
rect 23029 17561 23063 17595
rect 20913 17493 20947 17527
rect 23765 17493 23799 17527
rect 24685 17493 24719 17527
rect 25421 17493 25455 17527
rect 26525 17493 26559 17527
rect 25237 17289 25271 17323
rect 24501 17221 24535 17255
rect 24593 17221 24627 17255
rect 20545 17153 20579 17187
rect 21281 17153 21315 17187
rect 22109 17153 22143 17187
rect 22845 17153 22879 17187
rect 25329 17153 25363 17187
rect 26433 17153 26467 17187
rect 36093 17153 36127 17187
rect 22293 17085 22327 17119
rect 25789 17085 25823 17119
rect 24041 17017 24075 17051
rect 36277 17017 36311 17051
rect 20637 16949 20671 16983
rect 21373 16949 21407 16983
rect 22937 16949 22971 16983
rect 26525 16949 26559 16983
rect 27905 16745 27939 16779
rect 19625 16609 19659 16643
rect 20729 16609 20763 16643
rect 22569 16609 22603 16643
rect 22753 16609 22787 16643
rect 24685 16609 24719 16643
rect 26249 16609 26283 16643
rect 26709 16609 26743 16643
rect 1869 16541 1903 16575
rect 20269 16541 20303 16575
rect 21005 16541 21039 16575
rect 23673 16541 23707 16575
rect 24777 16541 24811 16575
rect 25421 16541 25455 16575
rect 27445 16541 27479 16575
rect 21833 16473 21867 16507
rect 26617 16473 26651 16507
rect 1685 16405 1719 16439
rect 20177 16405 20211 16439
rect 21925 16405 21959 16439
rect 23213 16405 23247 16439
rect 23857 16405 23891 16439
rect 25329 16405 25363 16439
rect 27353 16405 27387 16439
rect 11713 16201 11747 16235
rect 19073 16201 19107 16235
rect 21465 16201 21499 16235
rect 22569 16133 22603 16167
rect 24961 16133 24995 16167
rect 25053 16133 25087 16167
rect 11897 16065 11931 16099
rect 12449 16065 12483 16099
rect 19625 16065 19659 16099
rect 20269 16065 20303 16099
rect 23581 16065 23615 16099
rect 26065 16065 26099 16099
rect 27353 16065 27387 16099
rect 27813 16065 27847 16099
rect 20453 15997 20487 16031
rect 22477 15997 22511 16031
rect 24409 15997 24443 16031
rect 26249 15997 26283 16031
rect 28457 15997 28491 16031
rect 23029 15929 23063 15963
rect 19717 15861 19751 15895
rect 20913 15861 20947 15895
rect 23673 15861 23707 15895
rect 25605 15861 25639 15895
rect 27261 15861 27295 15895
rect 27905 15861 27939 15895
rect 36369 15861 36403 15895
rect 18889 15657 18923 15691
rect 29009 15657 29043 15691
rect 33609 15657 33643 15691
rect 20821 15521 20855 15555
rect 22569 15521 22603 15555
rect 23213 15521 23247 15555
rect 25145 15521 25179 15555
rect 27721 15521 27755 15555
rect 36093 15521 36127 15555
rect 18337 15453 18371 15487
rect 27169 15453 27203 15487
rect 27621 15453 27655 15487
rect 31677 15453 31711 15487
rect 33425 15453 33459 15487
rect 36369 15453 36403 15487
rect 19993 15385 20027 15419
rect 20177 15385 20211 15419
rect 20913 15385 20947 15419
rect 21465 15385 21499 15419
rect 21925 15385 21959 15419
rect 22477 15385 22511 15419
rect 23305 15385 23339 15419
rect 23857 15385 23891 15419
rect 25329 15385 25363 15419
rect 25421 15385 25455 15419
rect 26525 15385 26559 15419
rect 26617 15385 26651 15419
rect 31585 15385 31619 15419
rect 19533 15317 19567 15351
rect 28273 15317 28307 15351
rect 32229 15317 32263 15351
rect 19073 15113 19107 15147
rect 27169 15113 27203 15147
rect 29193 15113 29227 15147
rect 36093 15113 36127 15147
rect 20269 15045 20303 15079
rect 21373 15045 21407 15079
rect 22293 15045 22327 15079
rect 25237 15045 25271 15079
rect 27905 15045 27939 15079
rect 17233 14977 17267 15011
rect 17877 14977 17911 15011
rect 18981 14977 19015 15011
rect 19625 14977 19659 15011
rect 19809 14977 19843 15011
rect 20729 14977 20763 15011
rect 20913 14977 20947 15011
rect 23489 14977 23523 15011
rect 25881 14977 25915 15011
rect 26065 14977 26099 15011
rect 27997 14977 28031 15011
rect 28641 14977 28675 15011
rect 29285 14977 29319 15011
rect 35909 14977 35943 15011
rect 18521 14909 18555 14943
rect 22201 14909 22235 14943
rect 23673 14909 23707 14943
rect 25329 14909 25363 14943
rect 28549 14909 28583 14943
rect 29745 14909 29779 14943
rect 22753 14841 22787 14875
rect 23857 14841 23891 14875
rect 24777 14841 24811 14875
rect 17693 14773 17727 14807
rect 26249 14773 26283 14807
rect 18153 14569 18187 14603
rect 22293 14569 22327 14603
rect 22845 14569 22879 14603
rect 24685 14569 24719 14603
rect 20085 14433 20119 14467
rect 20821 14433 20855 14467
rect 21649 14433 21683 14467
rect 23581 14433 23615 14467
rect 25973 14433 26007 14467
rect 29101 14433 29135 14467
rect 1869 14365 1903 14399
rect 18705 14365 18739 14399
rect 19901 14365 19935 14399
rect 22201 14365 22235 14399
rect 23397 14365 23431 14399
rect 24777 14365 24811 14399
rect 26157 14365 26191 14399
rect 28549 14365 28583 14399
rect 29009 14365 29043 14399
rect 29929 14365 29963 14399
rect 21557 14297 21591 14331
rect 26617 14297 26651 14331
rect 27169 14297 27203 14331
rect 27261 14297 27295 14331
rect 27905 14297 27939 14331
rect 27997 14297 28031 14331
rect 29837 14297 29871 14331
rect 1685 14229 1719 14263
rect 18797 14229 18831 14263
rect 19441 14229 19475 14263
rect 24041 14229 24075 14263
rect 25513 14229 25547 14263
rect 30481 14229 30515 14263
rect 17049 14025 17083 14059
rect 17693 14025 17727 14059
rect 19441 14025 19475 14059
rect 22109 14025 22143 14059
rect 22753 14025 22787 14059
rect 24501 14025 24535 14059
rect 28825 14025 28859 14059
rect 30205 14025 30239 14059
rect 30849 14025 30883 14059
rect 20085 13957 20119 13991
rect 20177 13957 20211 13991
rect 21281 13957 21315 13991
rect 23765 13957 23799 13991
rect 25697 13957 25731 13991
rect 25789 13957 25823 13991
rect 27629 13957 27663 13991
rect 27721 13957 27755 13991
rect 18153 13889 18187 13923
rect 21373 13889 21407 13923
rect 22017 13889 22051 13923
rect 24593 13889 24627 13923
rect 26525 13889 26559 13923
rect 28917 13889 28951 13923
rect 29653 13889 29687 13923
rect 30113 13889 30147 13923
rect 30941 13889 30975 13923
rect 18797 13821 18831 13855
rect 18981 13821 19015 13855
rect 20729 13821 20763 13855
rect 23397 13821 23431 13855
rect 23857 13821 23891 13855
rect 25513 13821 25547 13855
rect 29561 13821 29595 13855
rect 26433 13753 26467 13787
rect 28181 13753 28215 13787
rect 18245 13685 18279 13719
rect 17601 13481 17635 13515
rect 18797 13481 18831 13515
rect 22293 13481 22327 13515
rect 21649 13413 21683 13447
rect 29101 13413 29135 13447
rect 29929 13413 29963 13447
rect 17049 13345 17083 13379
rect 19533 13345 19567 13379
rect 21097 13345 21131 13379
rect 26065 13345 26099 13379
rect 26617 13345 26651 13379
rect 30389 13345 30423 13379
rect 18061 13277 18095 13311
rect 18889 13277 18923 13311
rect 22201 13277 22235 13311
rect 24777 13277 24811 13311
rect 29009 13277 29043 13311
rect 29745 13277 29779 13311
rect 31769 13277 31803 13311
rect 36093 13277 36127 13311
rect 19625 13209 19659 13243
rect 20177 13209 20211 13243
rect 21189 13209 21223 13243
rect 22937 13209 22971 13243
rect 23489 13209 23523 13243
rect 23581 13209 23615 13243
rect 25421 13209 25455 13243
rect 25973 13209 26007 13243
rect 27169 13209 27203 13243
rect 27261 13209 27295 13243
rect 27813 13209 27847 13243
rect 28365 13209 28399 13243
rect 28457 13209 28491 13243
rect 31677 13209 31711 13243
rect 18153 13141 18187 13175
rect 24593 13141 24627 13175
rect 36277 13141 36311 13175
rect 2421 12937 2455 12971
rect 18521 12937 18555 12971
rect 21189 12937 21223 12971
rect 28549 12937 28583 12971
rect 22569 12869 22603 12903
rect 22661 12869 22695 12903
rect 23857 12869 23891 12903
rect 25421 12869 25455 12903
rect 27445 12869 27479 12903
rect 1869 12801 1903 12835
rect 2513 12801 2547 12835
rect 17417 12801 17451 12835
rect 18061 12801 18095 12835
rect 18981 12801 19015 12835
rect 19165 12801 19199 12835
rect 20637 12801 20671 12835
rect 21281 12801 21315 12835
rect 26065 12801 26099 12835
rect 26157 12801 26191 12835
rect 27997 12801 28031 12835
rect 28641 12801 28675 12835
rect 29101 12801 29135 12835
rect 17877 12733 17911 12767
rect 22385 12733 22419 12767
rect 23765 12733 23799 12767
rect 24869 12733 24903 12767
rect 25513 12733 25547 12767
rect 27353 12733 27387 12767
rect 3065 12665 3099 12699
rect 24317 12665 24351 12699
rect 29745 12665 29779 12699
rect 1685 12597 1719 12631
rect 17325 12597 17359 12631
rect 19625 12597 19659 12631
rect 20545 12597 20579 12631
rect 29193 12597 29227 12631
rect 17693 12393 17727 12427
rect 20637 12393 20671 12427
rect 21189 12393 21223 12427
rect 27905 12393 27939 12427
rect 28549 12393 28583 12427
rect 29101 12393 29135 12427
rect 18889 12325 18923 12359
rect 19809 12325 19843 12359
rect 21833 12325 21867 12359
rect 29745 12325 29779 12359
rect 12725 12257 12759 12291
rect 19441 12257 19475 12291
rect 22385 12257 22419 12291
rect 23581 12257 23615 12291
rect 24685 12257 24719 12291
rect 25697 12257 25731 12291
rect 26709 12257 26743 12291
rect 8125 12189 8159 12223
rect 12633 12189 12667 12223
rect 17785 12189 17819 12223
rect 18245 12189 18279 12223
rect 18429 12189 18463 12223
rect 19625 12189 19659 12223
rect 20545 12189 20579 12223
rect 24777 12189 24811 12223
rect 27353 12189 27387 12223
rect 27813 12189 27847 12223
rect 28641 12189 28675 12223
rect 30389 12189 30423 12223
rect 22293 12121 22327 12155
rect 22937 12121 22971 12155
rect 23489 12121 23523 12155
rect 25789 12121 25823 12155
rect 7941 12053 7975 12087
rect 13277 12053 13311 12087
rect 27261 12053 27295 12087
rect 17601 11849 17635 11883
rect 18153 11849 18187 11883
rect 21189 11849 21223 11883
rect 23305 11849 23339 11883
rect 27261 11849 27295 11883
rect 28549 11849 28583 11883
rect 29837 11849 29871 11883
rect 8309 11781 8343 11815
rect 20085 11781 20119 11815
rect 22569 11781 22603 11815
rect 25053 11781 25087 11815
rect 25145 11781 25179 11815
rect 26249 11781 26283 11815
rect 14289 11713 14323 11747
rect 17693 11713 17727 11747
rect 21097 11713 21131 11747
rect 23397 11713 23431 11747
rect 25697 11713 25731 11747
rect 27353 11713 27387 11747
rect 27813 11713 27847 11747
rect 28457 11713 28491 11747
rect 29101 11713 29135 11747
rect 29745 11713 29779 11747
rect 19257 11645 19291 11679
rect 19441 11645 19475 11679
rect 19993 11645 20027 11679
rect 20637 11645 20671 11679
rect 22385 11645 22419 11679
rect 22661 11645 22695 11679
rect 24133 11645 24167 11679
rect 26341 11645 26375 11679
rect 27905 11645 27939 11679
rect 14105 11577 14139 11611
rect 14841 11577 14875 11611
rect 29193 11577 29227 11611
rect 19073 11509 19107 11543
rect 17509 11305 17543 11339
rect 18153 11305 18187 11339
rect 18797 11305 18831 11339
rect 24685 11305 24719 11339
rect 30481 11305 30515 11339
rect 19533 11169 19567 11203
rect 21097 11169 21131 11203
rect 21741 11169 21775 11203
rect 22937 11169 22971 11203
rect 25789 11169 25823 11203
rect 27077 11169 27111 11203
rect 27721 11169 27755 11203
rect 29837 11169 29871 11203
rect 1869 11101 1903 11135
rect 16957 11101 16991 11135
rect 17601 11101 17635 11135
rect 18061 11101 18095 11135
rect 18889 11101 18923 11135
rect 23397 11101 23431 11135
rect 24777 11101 24811 11135
rect 28549 11101 28583 11135
rect 29929 11101 29963 11135
rect 30389 11101 30423 11135
rect 36093 11101 36127 11135
rect 16865 11033 16899 11067
rect 19625 11033 19659 11067
rect 20545 11033 20579 11067
rect 21189 11033 21223 11067
rect 22293 11033 22327 11067
rect 22385 11033 22419 11067
rect 25513 11033 25547 11067
rect 25605 11033 25639 11067
rect 27169 11033 27203 11067
rect 35633 11033 35667 11067
rect 36277 11033 36311 11067
rect 1685 10965 1719 10999
rect 23581 10965 23615 10999
rect 28641 10965 28675 10999
rect 17417 10761 17451 10795
rect 28825 10761 28859 10795
rect 30113 10761 30147 10795
rect 18705 10693 18739 10727
rect 20269 10693 20303 10727
rect 22017 10693 22051 10727
rect 22937 10693 22971 10727
rect 24501 10693 24535 10727
rect 25789 10693 25823 10727
rect 25881 10693 25915 10727
rect 27261 10693 27295 10727
rect 27353 10693 27387 10727
rect 29469 10693 29503 10727
rect 17877 10625 17911 10659
rect 28917 10625 28951 10659
rect 29561 10625 29595 10659
rect 30021 10625 30055 10659
rect 18613 10557 18647 10591
rect 19625 10557 19659 10591
rect 20177 10557 20211 10591
rect 21189 10557 21223 10591
rect 23029 10557 23063 10591
rect 23581 10557 23615 10591
rect 24593 10557 24627 10591
rect 27721 10557 27755 10591
rect 26341 10489 26375 10523
rect 17969 10421 18003 10455
rect 25145 10421 25179 10455
rect 36369 10421 36403 10455
rect 7573 10217 7607 10251
rect 18153 10217 18187 10251
rect 18797 10217 18831 10251
rect 25329 10217 25363 10251
rect 27721 10217 27755 10251
rect 28365 10217 28399 10251
rect 22201 10149 22235 10183
rect 26433 10149 26467 10183
rect 26985 10149 27019 10183
rect 22845 10081 22879 10115
rect 23121 10081 23155 10115
rect 23949 10081 23983 10115
rect 36093 10081 36127 10115
rect 7665 10013 7699 10047
rect 18245 10013 18279 10047
rect 18889 10013 18923 10047
rect 25329 10013 25363 10047
rect 27169 10013 27203 10047
rect 27629 10013 27663 10047
rect 28457 10013 28491 10047
rect 29101 10013 29135 10047
rect 36369 10013 36403 10047
rect 8217 9945 8251 9979
rect 19717 9945 19751 9979
rect 19809 9945 19843 9979
rect 20729 9945 20763 9979
rect 21649 9945 21683 9979
rect 21741 9945 21775 9979
rect 22946 9945 22980 9979
rect 25881 9945 25915 9979
rect 25982 9945 26016 9979
rect 29009 9945 29043 9979
rect 17601 9877 17635 9911
rect 34989 9877 35023 9911
rect 19441 9673 19475 9707
rect 17601 9605 17635 9639
rect 20177 9605 20211 9639
rect 20269 9605 20303 9639
rect 20821 9605 20855 9639
rect 26525 9605 26559 9639
rect 27905 9605 27939 9639
rect 36369 9605 36403 9639
rect 17141 9537 17175 9571
rect 18153 9537 18187 9571
rect 18981 9537 19015 9571
rect 21281 9537 21315 9571
rect 21373 9537 21407 9571
rect 26625 9537 26659 9571
rect 27169 9537 27203 9571
rect 27997 9537 28031 9571
rect 18797 9469 18831 9503
rect 22017 9469 22051 9503
rect 22293 9469 22327 9503
rect 24225 9469 24259 9503
rect 24501 9469 24535 9503
rect 27261 9401 27295 9435
rect 28549 9401 28583 9435
rect 18245 9333 18279 9367
rect 23765 9333 23799 9367
rect 25973 9333 26007 9367
rect 29009 9333 29043 9367
rect 33057 9333 33091 9367
rect 33793 9333 33827 9367
rect 34253 9333 34287 9367
rect 35173 9333 35207 9367
rect 35817 9333 35851 9367
rect 2421 9129 2455 9163
rect 18889 9129 18923 9163
rect 26341 9129 26375 9163
rect 32321 9129 32355 9163
rect 32873 9129 32907 9163
rect 18429 8993 18463 9027
rect 19441 8993 19475 9027
rect 20453 8993 20487 9027
rect 22845 8993 22879 9027
rect 24593 8993 24627 9027
rect 24869 8993 24903 9027
rect 26801 8993 26835 9027
rect 1869 8925 1903 8959
rect 17785 8925 17819 8959
rect 18245 8925 18279 8959
rect 33701 8925 33735 8959
rect 34253 8925 34287 8959
rect 17693 8857 17727 8891
rect 20361 8857 20395 8891
rect 22569 8857 22603 8891
rect 23305 8857 23339 8891
rect 23857 8857 23891 8891
rect 23949 8857 23983 8891
rect 27077 8857 27111 8891
rect 35909 8857 35943 8891
rect 1685 8789 1719 8823
rect 21097 8789 21131 8823
rect 28549 8789 28583 8823
rect 29101 8789 29135 8823
rect 34897 8789 34931 8823
rect 17877 8517 17911 8551
rect 18613 8517 18647 8551
rect 19901 8517 19935 8551
rect 31769 8517 31803 8551
rect 32505 8517 32539 8551
rect 17785 8449 17819 8483
rect 19625 8449 19659 8483
rect 23857 8449 23891 8483
rect 24317 8449 24351 8483
rect 27353 8449 27387 8483
rect 33241 8449 33275 8483
rect 18521 8381 18555 8415
rect 24593 8381 24627 8415
rect 27261 8381 27295 8415
rect 27905 8381 27939 8415
rect 29653 8381 29687 8415
rect 29929 8381 29963 8415
rect 19073 8313 19107 8347
rect 22109 8313 22143 8347
rect 30389 8313 30423 8347
rect 33149 8313 33183 8347
rect 33793 8313 33827 8347
rect 34989 8313 35023 8347
rect 36277 8313 36311 8347
rect 21373 8245 21407 8279
rect 23593 8245 23627 8279
rect 26065 8245 26099 8279
rect 34253 8245 34287 8279
rect 35449 8245 35483 8279
rect 23305 8041 23339 8075
rect 23949 8041 23983 8075
rect 24685 8041 24719 8075
rect 26598 8041 26632 8075
rect 31769 8041 31803 8075
rect 22661 7973 22695 8007
rect 28089 7973 28123 8007
rect 20085 7905 20119 7939
rect 20913 7905 20947 7939
rect 25329 7905 25363 7939
rect 25881 7905 25915 7939
rect 26341 7905 26375 7939
rect 33609 7905 33643 7939
rect 34897 7905 34931 7939
rect 36093 7905 36127 7939
rect 18061 7837 18095 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 19901 7837 19935 7871
rect 23397 7837 23431 7871
rect 24041 7837 24075 7871
rect 24777 7837 24811 7871
rect 33057 7837 33091 7871
rect 33149 7837 33183 7871
rect 36369 7837 36403 7871
rect 17601 7769 17635 7803
rect 21189 7769 21223 7803
rect 31217 7769 31251 7803
rect 18153 7701 18187 7735
rect 19441 7701 19475 7735
rect 28733 7701 28767 7735
rect 29745 7701 29779 7735
rect 32321 7701 32355 7735
rect 34161 7701 34195 7735
rect 22109 7497 22143 7531
rect 22753 7497 22787 7531
rect 25789 7497 25823 7531
rect 26433 7497 26467 7531
rect 29745 7497 29779 7531
rect 36369 7497 36403 7531
rect 17325 7429 17359 7463
rect 18245 7429 18279 7463
rect 19073 7429 19107 7463
rect 27169 7429 27203 7463
rect 33793 7429 33827 7463
rect 35449 7429 35483 7463
rect 1869 7361 1903 7395
rect 20453 7361 20487 7395
rect 22201 7361 22235 7395
rect 22661 7361 22695 7395
rect 23489 7361 23523 7395
rect 30665 7361 30699 7395
rect 31217 7361 31251 7395
rect 32597 7361 32631 7395
rect 33241 7361 33275 7395
rect 33885 7361 33919 7395
rect 34345 7361 34379 7395
rect 34897 7361 34931 7395
rect 18337 7293 18371 7327
rect 18981 7293 19015 7327
rect 19993 7293 20027 7327
rect 20637 7293 20671 7327
rect 23397 7293 23431 7327
rect 24041 7293 24075 7327
rect 24317 7293 24351 7327
rect 28917 7293 28951 7327
rect 29193 7293 29227 7327
rect 20821 7225 20855 7259
rect 32505 7225 32539 7259
rect 1685 7157 1719 7191
rect 31769 7157 31803 7191
rect 33149 7157 33183 7191
rect 35541 6953 35575 6987
rect 20085 6885 20119 6919
rect 17417 6817 17451 6851
rect 20821 6817 20855 6851
rect 22845 6817 22879 6851
rect 23305 6817 23339 6851
rect 23949 6817 23983 6851
rect 24685 6817 24719 6851
rect 25237 6817 25271 6851
rect 25697 6817 25731 6851
rect 32873 6817 32907 6851
rect 34161 6817 34195 6851
rect 9137 6749 9171 6783
rect 17509 6749 17543 6783
rect 17969 6749 18003 6783
rect 18061 6749 18095 6783
rect 18797 6749 18831 6783
rect 31493 6749 31527 6783
rect 32321 6749 32355 6783
rect 32965 6749 32999 6783
rect 33609 6749 33643 6783
rect 34253 6749 34287 6783
rect 35081 6749 35115 6783
rect 36093 6749 36127 6783
rect 19533 6681 19567 6715
rect 19625 6681 19659 6715
rect 21097 6681 21131 6715
rect 25973 6681 26007 6715
rect 9229 6613 9263 6647
rect 18705 6613 18739 6647
rect 27445 6613 27479 6647
rect 28089 6613 28123 6647
rect 28641 6613 28675 6647
rect 29193 6613 29227 6647
rect 29745 6613 29779 6647
rect 30757 6613 30791 6647
rect 32229 6613 32263 6647
rect 33517 6613 33551 6647
rect 34989 6613 35023 6647
rect 1777 6409 1811 6443
rect 18613 6409 18647 6443
rect 31677 6409 31711 6443
rect 32597 6409 32631 6443
rect 34529 6409 34563 6443
rect 36277 6409 36311 6443
rect 19993 6341 20027 6375
rect 24869 6341 24903 6375
rect 35725 6341 35759 6375
rect 1961 6273 1995 6307
rect 17417 6273 17451 6307
rect 17969 6273 18003 6307
rect 19257 6273 19291 6307
rect 19717 6273 19751 6307
rect 23857 6273 23891 6307
rect 24593 6273 24627 6307
rect 31769 6273 31803 6307
rect 32689 6273 32723 6307
rect 33333 6273 33367 6307
rect 33977 6273 34011 6307
rect 34621 6273 34655 6307
rect 35265 6273 35299 6307
rect 19073 6205 19107 6239
rect 22109 6205 22143 6239
rect 23581 6205 23615 6239
rect 26617 6205 26651 6239
rect 27813 6205 27847 6239
rect 29285 6205 29319 6239
rect 29561 6205 29595 6239
rect 33241 6205 33275 6239
rect 18061 6137 18095 6171
rect 33885 6137 33919 6171
rect 21465 6069 21499 6103
rect 27169 6069 27203 6103
rect 30021 6069 30055 6103
rect 30573 6069 30607 6103
rect 35173 6069 35207 6103
rect 2329 5865 2363 5899
rect 17325 5865 17359 5899
rect 18613 5865 18647 5899
rect 29101 5865 29135 5899
rect 30002 5865 30036 5899
rect 31493 5865 31527 5899
rect 32045 5865 32079 5899
rect 33333 5865 33367 5899
rect 23397 5797 23431 5831
rect 32689 5797 32723 5831
rect 33977 5797 34011 5831
rect 20821 5729 20855 5763
rect 22845 5729 22879 5763
rect 27353 5729 27387 5763
rect 36093 5729 36127 5763
rect 1869 5661 1903 5695
rect 17233 5661 17267 5695
rect 17877 5661 17911 5695
rect 18521 5661 18555 5695
rect 20177 5661 20211 5695
rect 29745 5661 29779 5695
rect 32137 5661 32171 5695
rect 32781 5661 32815 5695
rect 33425 5661 33459 5695
rect 34069 5661 34103 5695
rect 35081 5661 35115 5695
rect 36369 5661 36403 5695
rect 19533 5593 19567 5627
rect 19625 5593 19659 5627
rect 21097 5593 21131 5627
rect 23949 5593 23983 5627
rect 24685 5593 24719 5627
rect 26709 5593 26743 5627
rect 27629 5593 27663 5627
rect 1685 5525 1719 5559
rect 16681 5525 16715 5559
rect 17969 5525 18003 5559
rect 25513 5525 25547 5559
rect 26065 5525 26099 5559
rect 34989 5525 35023 5559
rect 19073 5321 19107 5355
rect 19717 5321 19751 5355
rect 28917 5321 28951 5355
rect 34253 5321 34287 5355
rect 34897 5321 34931 5355
rect 35449 5321 35483 5355
rect 17417 5253 17451 5287
rect 18337 5253 18371 5287
rect 30389 5253 30423 5287
rect 14565 5185 14599 5219
rect 15209 5185 15243 5219
rect 18981 5185 19015 5219
rect 19625 5185 19659 5219
rect 27169 5185 27203 5219
rect 30481 5185 30515 5219
rect 31033 5185 31067 5219
rect 31125 5185 31159 5219
rect 31769 5185 31803 5219
rect 32413 5185 32447 5219
rect 32505 5185 32539 5219
rect 33149 5185 33183 5219
rect 33793 5185 33827 5219
rect 35909 5185 35943 5219
rect 17325 5117 17359 5151
rect 33701 5117 33735 5151
rect 14657 5049 14691 5083
rect 22017 5049 22051 5083
rect 24961 5049 24995 5083
rect 33057 5049 33091 5083
rect 23029 4981 23063 5015
rect 23673 4981 23707 5015
rect 24133 4981 24167 5015
rect 25513 4981 25547 5015
rect 26065 4981 26099 5015
rect 26525 4981 26559 5015
rect 27432 4981 27466 5015
rect 29653 4981 29687 5015
rect 31677 4981 31711 5015
rect 16773 4777 16807 4811
rect 22661 4777 22695 4811
rect 35449 4777 35483 4811
rect 18153 4709 18187 4743
rect 29745 4709 29779 4743
rect 15117 4641 15151 4675
rect 17325 4641 17359 4675
rect 20913 4641 20947 4675
rect 21189 4641 21223 4675
rect 23121 4641 23155 4675
rect 23765 4641 23799 4675
rect 24685 4641 24719 4675
rect 25237 4641 25271 4675
rect 25789 4641 25823 4675
rect 26341 4641 26375 4675
rect 26893 4641 26927 4675
rect 27353 4641 27387 4675
rect 31217 4641 31251 4675
rect 32597 4641 32631 4675
rect 13093 4573 13127 4607
rect 13553 4573 13587 4607
rect 14289 4573 14323 4607
rect 14841 4573 14875 4607
rect 16865 4573 16899 4607
rect 31493 4573 31527 4607
rect 32689 4573 32723 4607
rect 33333 4573 33367 4607
rect 33977 4573 34011 4607
rect 34897 4573 34931 4607
rect 36093 4573 36127 4607
rect 13645 4505 13679 4539
rect 27629 4505 27663 4539
rect 33241 4505 33275 4539
rect 29101 4437 29135 4471
rect 32045 4437 32079 4471
rect 33885 4437 33919 4471
rect 36277 4437 36311 4471
rect 13461 4233 13495 4267
rect 21373 4233 21407 4267
rect 29929 4165 29963 4199
rect 13921 4097 13955 4131
rect 14841 4097 14875 4131
rect 15761 4097 15795 4131
rect 17785 4097 17819 4131
rect 17877 4097 17911 4131
rect 18981 4097 19015 4131
rect 19073 4097 19107 4131
rect 22109 4097 22143 4131
rect 26065 4097 26099 4131
rect 26525 4097 26559 4131
rect 32413 4097 32447 4131
rect 32505 4097 32539 4131
rect 33057 4097 33091 4131
rect 33149 4097 33183 4131
rect 33793 4097 33827 4131
rect 35909 4097 35943 4131
rect 14197 4029 14231 4063
rect 15117 4029 15151 4063
rect 22385 4029 22419 4063
rect 24317 4029 24351 4063
rect 25789 4029 25823 4063
rect 27445 4029 27479 4063
rect 28917 4029 28951 4063
rect 29193 4029 29227 4063
rect 29653 4029 29687 4063
rect 34345 3961 34379 3995
rect 23857 3893 23891 3927
rect 31401 3893 31435 3927
rect 33701 3893 33735 3927
rect 34805 3893 34839 3927
rect 35449 3893 35483 3927
rect 14289 3689 14323 3723
rect 20453 3689 20487 3723
rect 29101 3689 29135 3723
rect 32689 3689 32723 3723
rect 34897 3689 34931 3723
rect 10333 3621 10367 3655
rect 22661 3621 22695 3655
rect 29745 3621 29779 3655
rect 33333 3621 33367 3655
rect 36093 3621 36127 3655
rect 15117 3553 15151 3587
rect 18061 3553 18095 3587
rect 23765 3553 23799 3587
rect 24041 3553 24075 3587
rect 24593 3553 24627 3587
rect 26801 3553 26835 3587
rect 31493 3553 31527 3587
rect 1869 3485 1903 3519
rect 10517 3485 10551 3519
rect 14841 3485 14875 3519
rect 20913 3485 20947 3519
rect 32137 3485 32171 3519
rect 32781 3485 32815 3519
rect 33425 3485 33459 3519
rect 34069 3485 34103 3519
rect 36277 3485 36311 3519
rect 21189 3417 21223 3451
rect 24869 3417 24903 3451
rect 27077 3417 27111 3451
rect 31217 3417 31251 3451
rect 33977 3417 34011 3451
rect 1685 3349 1719 3383
rect 26341 3349 26375 3383
rect 28549 3349 28583 3383
rect 32045 3349 32079 3383
rect 35541 3349 35575 3383
rect 12541 3145 12575 3179
rect 13277 3145 13311 3179
rect 16957 3145 16991 3179
rect 19717 3145 19751 3179
rect 33149 3145 33183 3179
rect 22017 3077 22051 3111
rect 25881 3077 25915 3111
rect 26433 3077 26467 3111
rect 26617 3077 26651 3111
rect 34989 3077 35023 3111
rect 1869 3009 1903 3043
rect 11897 3009 11931 3043
rect 12725 3009 12759 3043
rect 14289 3009 14323 3043
rect 14841 3009 14875 3043
rect 16129 3009 16163 3043
rect 21465 3009 21499 3043
rect 22937 3009 22971 3043
rect 23857 3009 23891 3043
rect 28917 3009 28951 3043
rect 29377 3009 29411 3043
rect 31677 3009 31711 3043
rect 31769 3009 31803 3043
rect 32321 3009 32355 3043
rect 33241 3009 33275 3043
rect 33885 3009 33919 3043
rect 36093 3009 36127 3043
rect 21189 2941 21223 2975
rect 24133 2941 24167 2975
rect 28641 2941 28675 2975
rect 29653 2941 29687 2975
rect 33793 2941 33827 2975
rect 36369 2941 36403 2975
rect 15945 2873 15979 2907
rect 27169 2873 27203 2907
rect 32505 2873 32539 2907
rect 34805 2873 34839 2907
rect 1685 2805 1719 2839
rect 11713 2805 11747 2839
rect 14105 2805 14139 2839
rect 22753 2805 22787 2839
rect 31125 2805 31159 2839
rect 2513 2601 2547 2635
rect 4721 2601 4755 2635
rect 19441 2601 19475 2635
rect 22017 2601 22051 2635
rect 29101 2601 29135 2635
rect 31493 2601 31527 2635
rect 33701 2601 33735 2635
rect 36185 2601 36219 2635
rect 9413 2533 9447 2567
rect 23765 2465 23799 2499
rect 24593 2465 24627 2499
rect 24869 2465 24903 2499
rect 26341 2465 26375 2499
rect 27353 2465 27387 2499
rect 27629 2465 27663 2499
rect 29745 2465 29779 2499
rect 30021 2465 30055 2499
rect 35173 2465 35207 2499
rect 1869 2397 1903 2431
rect 2329 2397 2363 2431
rect 4261 2397 4295 2431
rect 5549 2397 5583 2431
rect 6837 2397 6871 2431
rect 11989 2397 12023 2431
rect 14565 2397 14599 2431
rect 15853 2397 15887 2431
rect 17785 2397 17819 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 32321 2397 32355 2431
rect 32597 2397 32631 2431
rect 33793 2397 33827 2431
rect 34897 2397 34931 2431
rect 2973 2329 3007 2363
rect 9229 2329 9263 2363
rect 9965 2329 9999 2363
rect 10517 2329 10551 2363
rect 23489 2329 23523 2363
rect 1685 2261 1719 2295
rect 4077 2261 4111 2295
rect 5365 2261 5399 2295
rect 6653 2261 6687 2295
rect 8493 2261 8527 2295
rect 10609 2261 10643 2295
rect 11805 2261 11839 2295
rect 14381 2261 14415 2295
rect 15669 2261 15703 2295
rect 17601 2261 17635 2295
rect 18337 2261 18371 2295
rect 20821 2261 20855 2295
<< metal1 >>
rect 1104 37562 36892 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36892 37562
rect 1104 37488 36892 37510
rect 14 37408 20 37460
rect 72 37448 78 37460
rect 2869 37451 2927 37457
rect 2869 37448 2881 37451
rect 72 37420 2881 37448
rect 72 37408 78 37420
rect 2869 37417 2881 37420
rect 2915 37417 2927 37451
rect 2869 37411 2927 37417
rect 9493 37451 9551 37457
rect 9493 37417 9505 37451
rect 9539 37448 9551 37451
rect 13538 37448 13544 37460
rect 9539 37420 13544 37448
rect 9539 37417 9551 37420
rect 9493 37411 9551 37417
rect 13538 37408 13544 37420
rect 13596 37408 13602 37460
rect 16114 37408 16120 37460
rect 16172 37448 16178 37460
rect 16209 37451 16267 37457
rect 16209 37448 16221 37451
rect 16172 37420 16221 37448
rect 16172 37408 16178 37420
rect 16209 37417 16221 37420
rect 16255 37417 16267 37451
rect 16209 37411 16267 37417
rect 21266 37408 21272 37460
rect 21324 37448 21330 37460
rect 21361 37451 21419 37457
rect 21361 37448 21373 37451
rect 21324 37420 21373 37448
rect 21324 37408 21330 37420
rect 21361 37417 21373 37420
rect 21407 37417 21419 37451
rect 21361 37411 21419 37417
rect 2317 37383 2375 37389
rect 2317 37349 2329 37383
rect 2363 37380 2375 37383
rect 2363 37352 21312 37380
rect 2363 37349 2375 37352
rect 2317 37343 2375 37349
rect 5534 37312 5540 37324
rect 5495 37284 5540 37312
rect 5534 37272 5540 37284
rect 5592 37272 5598 37324
rect 6733 37315 6791 37321
rect 6733 37281 6745 37315
rect 6779 37312 6791 37315
rect 7098 37312 7104 37324
rect 6779 37284 7104 37312
rect 6779 37281 6791 37284
rect 6733 37275 6791 37281
rect 7098 37272 7104 37284
rect 7156 37312 7162 37324
rect 7193 37315 7251 37321
rect 7193 37312 7205 37315
rect 7156 37284 7205 37312
rect 7156 37272 7162 37284
rect 7193 37281 7205 37284
rect 7239 37281 7251 37315
rect 7193 37275 7251 37281
rect 10318 37272 10324 37324
rect 10376 37312 10382 37324
rect 11149 37315 11207 37321
rect 11149 37312 11161 37315
rect 10376 37284 11161 37312
rect 10376 37272 10382 37284
rect 11149 37281 11161 37284
rect 11195 37312 11207 37315
rect 11701 37315 11759 37321
rect 11701 37312 11713 37315
rect 11195 37284 11713 37312
rect 11195 37281 11207 37284
rect 11149 37275 11207 37281
rect 11701 37281 11713 37284
rect 11747 37281 11759 37315
rect 11701 37275 11759 37281
rect 13725 37315 13783 37321
rect 13725 37281 13737 37315
rect 13771 37312 13783 37315
rect 13771 37284 14228 37312
rect 13771 37281 13783 37284
rect 13725 37275 13783 37281
rect 14200 37256 14228 37284
rect 16114 37272 16120 37324
rect 16172 37312 16178 37324
rect 16172 37284 16574 37312
rect 16172 37272 16178 37284
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2133 37247 2191 37253
rect 2133 37244 2145 37247
rect 2004 37216 2145 37244
rect 2004 37204 2010 37216
rect 2133 37213 2145 37216
rect 2179 37213 2191 37247
rect 3050 37244 3056 37256
rect 3011 37216 3056 37244
rect 2133 37207 2191 37213
rect 3050 37204 3056 37216
rect 3108 37204 3114 37256
rect 3970 37244 3976 37256
rect 3931 37216 3976 37244
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 4801 37247 4859 37253
rect 4801 37213 4813 37247
rect 4847 37244 4859 37247
rect 5166 37244 5172 37256
rect 4847 37216 5172 37244
rect 4847 37213 4859 37216
rect 4801 37207 4859 37213
rect 5166 37204 5172 37216
rect 5224 37244 5230 37256
rect 5353 37247 5411 37253
rect 5353 37244 5365 37247
rect 5224 37216 5365 37244
rect 5224 37204 5230 37216
rect 5353 37213 5365 37216
rect 5399 37213 5411 37247
rect 7466 37244 7472 37256
rect 7427 37216 7472 37244
rect 5353 37207 5411 37213
rect 7466 37204 7472 37216
rect 7524 37204 7530 37256
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37244 8631 37247
rect 9030 37244 9036 37256
rect 8619 37216 9036 37244
rect 8619 37213 8631 37216
rect 8573 37207 8631 37213
rect 9030 37204 9036 37216
rect 9088 37244 9094 37256
rect 9217 37247 9275 37253
rect 9217 37244 9229 37247
rect 9088 37216 9229 37244
rect 9088 37204 9094 37216
rect 9217 37213 9229 37216
rect 9263 37213 9275 37247
rect 10870 37244 10876 37256
rect 10831 37216 10876 37244
rect 9217 37207 9275 37213
rect 10870 37204 10876 37216
rect 10928 37204 10934 37256
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 12529 37247 12587 37253
rect 12529 37244 12541 37247
rect 12492 37216 12541 37244
rect 12492 37204 12498 37216
rect 12529 37213 12541 37216
rect 12575 37244 12587 37247
rect 12989 37247 13047 37253
rect 12989 37244 13001 37247
rect 12575 37216 13001 37244
rect 12575 37213 12587 37216
rect 12529 37207 12587 37213
rect 12989 37213 13001 37216
rect 13035 37213 13047 37247
rect 12989 37207 13047 37213
rect 14182 37204 14188 37256
rect 14240 37244 14246 37256
rect 14369 37247 14427 37253
rect 14369 37244 14381 37247
rect 14240 37216 14381 37244
rect 14240 37204 14246 37216
rect 14369 37213 14381 37216
rect 14415 37213 14427 37247
rect 16546 37244 16574 37284
rect 17034 37272 17040 37324
rect 17092 37312 17098 37324
rect 17497 37315 17555 37321
rect 17497 37312 17509 37315
rect 17092 37284 17509 37312
rect 17092 37272 17098 37284
rect 17497 37281 17509 37284
rect 17543 37281 17555 37315
rect 18233 37315 18291 37321
rect 18233 37312 18245 37315
rect 17497 37275 17555 37281
rect 17696 37284 18245 37312
rect 16853 37247 16911 37253
rect 16853 37244 16865 37247
rect 16546 37216 16865 37244
rect 14369 37207 14427 37213
rect 16853 37213 16865 37216
rect 16899 37213 16911 37247
rect 16853 37207 16911 37213
rect 17402 37204 17408 37256
rect 17460 37244 17466 37256
rect 17696 37253 17724 37284
rect 18233 37281 18245 37284
rect 18279 37281 18291 37315
rect 18233 37275 18291 37281
rect 17681 37247 17739 37253
rect 17681 37244 17693 37247
rect 17460 37216 17693 37244
rect 17460 37204 17466 37216
rect 17681 37213 17693 37216
rect 17727 37213 17739 37247
rect 17681 37207 17739 37213
rect 18874 37204 18880 37256
rect 18932 37244 18938 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 18932 37216 19441 37244
rect 18932 37204 18938 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 8938 37136 8944 37188
rect 8996 37176 9002 37188
rect 21284 37176 21312 37352
rect 21376 37312 21404 37411
rect 22281 37383 22339 37389
rect 22281 37349 22293 37383
rect 22327 37380 22339 37383
rect 25498 37380 25504 37392
rect 22327 37352 25504 37380
rect 22327 37349 22339 37352
rect 22281 37343 22339 37349
rect 25498 37340 25504 37352
rect 25556 37340 25562 37392
rect 21376 37284 22140 37312
rect 22112 37253 22140 37284
rect 22646 37272 22652 37324
rect 22704 37312 22710 37324
rect 22741 37315 22799 37321
rect 22741 37312 22753 37315
rect 22704 37284 22753 37312
rect 22704 37272 22710 37284
rect 22741 37281 22753 37284
rect 22787 37281 22799 37315
rect 23477 37315 23535 37321
rect 23477 37312 23489 37315
rect 22741 37275 22799 37281
rect 22940 37284 23489 37312
rect 22097 37247 22155 37253
rect 22097 37213 22109 37247
rect 22143 37213 22155 37247
rect 22097 37207 22155 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22940 37253 22968 37284
rect 23477 37281 23489 37284
rect 23523 37281 23535 37315
rect 24854 37312 24860 37324
rect 24815 37284 24860 37312
rect 23477 37275 23535 37281
rect 24854 37272 24860 37284
rect 24912 37272 24918 37324
rect 35069 37315 35127 37321
rect 35069 37281 35081 37315
rect 35115 37312 35127 37315
rect 35526 37312 35532 37324
rect 35115 37284 35532 37312
rect 35115 37281 35127 37284
rect 35069 37275 35127 37281
rect 35526 37272 35532 37284
rect 35584 37272 35590 37324
rect 22925 37247 22983 37253
rect 22925 37244 22937 37247
rect 22612 37216 22937 37244
rect 22612 37204 22618 37216
rect 22925 37213 22937 37216
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24673 37247 24731 37253
rect 24673 37244 24685 37247
rect 24544 37216 24685 37244
rect 24544 37204 24550 37216
rect 24673 37213 24685 37216
rect 24719 37213 24731 37247
rect 24673 37207 24731 37213
rect 26786 37204 26792 37256
rect 26844 37244 26850 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 26844 37216 27169 37244
rect 26844 37204 26850 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 28721 37247 28779 37253
rect 28721 37213 28733 37247
rect 28767 37244 28779 37247
rect 28810 37244 28816 37256
rect 28767 37216 28816 37244
rect 28767 37213 28779 37216
rect 28721 37207 28779 37213
rect 28810 37204 28816 37216
rect 28868 37204 28874 37256
rect 29730 37244 29736 37256
rect 29691 37216 29736 37244
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 32309 37247 32367 37253
rect 32309 37213 32321 37247
rect 32355 37213 32367 37247
rect 32309 37207 32367 37213
rect 23198 37176 23204 37188
rect 8996 37148 12388 37176
rect 21284 37148 23204 37176
rect 8996 37136 9002 37148
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 12360 37117 12388 37148
rect 23198 37136 23204 37148
rect 23256 37136 23262 37188
rect 28626 37136 28632 37188
rect 28684 37176 28690 37188
rect 32324 37176 32352 37207
rect 33594 37204 33600 37256
rect 33652 37244 33658 37256
rect 33873 37247 33931 37253
rect 33873 37244 33885 37247
rect 33652 37216 33885 37244
rect 33652 37204 33658 37216
rect 33873 37213 33885 37216
rect 33919 37213 33931 37247
rect 35802 37244 35808 37256
rect 35763 37216 35808 37244
rect 33873 37207 33931 37213
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 28684 37148 32352 37176
rect 28684 37136 28690 37148
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3936 37080 4169 37108
rect 3936 37068 3942 37080
rect 4157 37077 4169 37080
rect 4203 37077 4215 37111
rect 4157 37071 4215 37077
rect 12345 37111 12403 37117
rect 12345 37077 12357 37111
rect 12391 37077 12403 37111
rect 14458 37108 14464 37120
rect 14419 37080 14464 37108
rect 12345 37071 12403 37077
rect 14458 37068 14464 37080
rect 14516 37068 14522 37120
rect 17037 37111 17095 37117
rect 17037 37077 17049 37111
rect 17083 37108 17095 37111
rect 19242 37108 19248 37120
rect 17083 37080 19248 37108
rect 17083 37077 17095 37080
rect 17037 37071 17095 37077
rect 19242 37068 19248 37080
rect 19300 37068 19306 37120
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19613 37111 19671 37117
rect 19613 37108 19625 37111
rect 19392 37080 19625 37108
rect 19392 37068 19398 37080
rect 19613 37077 19625 37080
rect 19659 37077 19671 37111
rect 19613 37071 19671 37077
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 26476 37080 27353 37108
rect 26476 37068 26482 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28350 37068 28356 37120
rect 28408 37108 28414 37120
rect 28537 37111 28595 37117
rect 28537 37108 28549 37111
rect 28408 37080 28549 37108
rect 28408 37068 28414 37080
rect 28537 37077 28549 37080
rect 28583 37077 28595 37111
rect 28537 37071 28595 37077
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29696 37080 29929 37108
rect 29696 37068 29702 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 31754 37068 31760 37120
rect 31812 37108 31818 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 31812 37080 32505 37108
rect 31812 37068 31818 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33689 37111 33747 37117
rect 33689 37108 33701 37111
rect 33560 37080 33701 37108
rect 33560 37068 33566 37080
rect 33689 37077 33701 37080
rect 33735 37077 33747 37111
rect 33689 37071 33747 37077
rect 1104 37018 36892 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 36892 37018
rect 1104 36944 36892 36966
rect 1670 36904 1676 36916
rect 1631 36876 1676 36904
rect 1670 36864 1676 36876
rect 1728 36864 1734 36916
rect 1946 36864 1952 36916
rect 2004 36904 2010 36916
rect 2317 36907 2375 36913
rect 2317 36904 2329 36907
rect 2004 36876 2329 36904
rect 2004 36864 2010 36876
rect 2317 36873 2329 36876
rect 2363 36873 2375 36907
rect 2317 36867 2375 36873
rect 3050 36864 3056 36916
rect 3108 36904 3114 36916
rect 4065 36907 4123 36913
rect 4065 36904 4077 36907
rect 3108 36876 4077 36904
rect 3108 36864 3114 36876
rect 4065 36873 4077 36876
rect 4111 36873 4123 36907
rect 18874 36904 18880 36916
rect 18835 36876 18880 36904
rect 4065 36867 4123 36873
rect 18874 36864 18880 36876
rect 18932 36864 18938 36916
rect 24486 36904 24492 36916
rect 24447 36876 24492 36904
rect 24486 36864 24492 36876
rect 24544 36864 24550 36916
rect 34790 36864 34796 36916
rect 34848 36904 34854 36916
rect 35069 36907 35127 36913
rect 35069 36904 35081 36907
rect 34848 36876 35081 36904
rect 34848 36864 34854 36876
rect 35069 36873 35081 36876
rect 35115 36873 35127 36907
rect 36262 36904 36268 36916
rect 36223 36876 36268 36904
rect 35069 36867 35127 36873
rect 36262 36864 36268 36876
rect 36320 36864 36326 36916
rect 10870 36796 10876 36848
rect 10928 36836 10934 36848
rect 10928 36808 18736 36836
rect 10928 36796 10934 36808
rect 1762 36728 1768 36780
rect 1820 36768 1826 36780
rect 1857 36771 1915 36777
rect 1857 36768 1869 36771
rect 1820 36740 1869 36768
rect 1820 36728 1826 36740
rect 1857 36737 1869 36740
rect 1903 36737 1915 36771
rect 1857 36731 1915 36737
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36768 4307 36771
rect 7466 36768 7472 36780
rect 4295 36740 7472 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 7466 36728 7472 36740
rect 7524 36768 7530 36780
rect 11054 36768 11060 36780
rect 7524 36740 11060 36768
rect 7524 36728 7530 36740
rect 11054 36728 11060 36740
rect 11112 36728 11118 36780
rect 17586 36768 17592 36780
rect 17547 36740 17592 36768
rect 17586 36728 17592 36740
rect 17644 36728 17650 36780
rect 18708 36777 18736 36808
rect 19242 36796 19248 36848
rect 19300 36836 19306 36848
rect 19300 36808 22600 36836
rect 19300 36796 19306 36808
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36768 18751 36771
rect 19426 36768 19432 36780
rect 18739 36740 19432 36768
rect 18739 36737 18751 36740
rect 18693 36731 18751 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 22572 36777 22600 36808
rect 22664 36808 26234 36836
rect 22557 36771 22615 36777
rect 22557 36737 22569 36771
rect 22603 36737 22615 36771
rect 22557 36731 22615 36737
rect 17773 36635 17831 36641
rect 17773 36601 17785 36635
rect 17819 36632 17831 36635
rect 22664 36632 22692 36808
rect 23198 36768 23204 36780
rect 23159 36740 23204 36768
rect 23198 36728 23204 36740
rect 23256 36768 23262 36780
rect 23382 36768 23388 36780
rect 23256 36740 23388 36768
rect 23256 36728 23262 36740
rect 23382 36728 23388 36740
rect 23440 36768 23446 36780
rect 23845 36771 23903 36777
rect 23845 36768 23857 36771
rect 23440 36740 23857 36768
rect 23440 36728 23446 36740
rect 23845 36737 23857 36740
rect 23891 36737 23903 36771
rect 26206 36768 26234 36808
rect 34885 36771 34943 36777
rect 34885 36768 34897 36771
rect 26206 36740 34897 36768
rect 23845 36731 23903 36737
rect 34885 36737 34897 36740
rect 34931 36737 34943 36771
rect 34885 36731 34943 36737
rect 35986 36728 35992 36780
rect 36044 36768 36050 36780
rect 36081 36771 36139 36777
rect 36081 36768 36093 36771
rect 36044 36740 36093 36768
rect 36044 36728 36050 36740
rect 36081 36737 36093 36740
rect 36127 36737 36139 36771
rect 36081 36731 36139 36737
rect 22756 36672 25084 36700
rect 22756 36641 22784 36672
rect 17819 36604 22692 36632
rect 22741 36635 22799 36641
rect 17819 36601 17831 36604
rect 17773 36595 17831 36601
rect 22741 36601 22753 36635
rect 22787 36601 22799 36635
rect 22741 36595 22799 36601
rect 23385 36635 23443 36641
rect 23385 36601 23397 36635
rect 23431 36632 23443 36635
rect 25056 36632 25084 36672
rect 29730 36632 29736 36644
rect 23431 36604 24992 36632
rect 25056 36604 29736 36632
rect 23431 36601 23443 36604
rect 23385 36595 23443 36601
rect 24964 36564 24992 36604
rect 29730 36592 29736 36604
rect 29788 36592 29794 36644
rect 28626 36564 28632 36576
rect 24964 36536 28632 36564
rect 28626 36524 28632 36536
rect 28684 36524 28690 36576
rect 28810 36564 28816 36576
rect 28771 36536 28816 36564
rect 28810 36524 28816 36536
rect 28868 36524 28874 36576
rect 33594 36524 33600 36576
rect 33652 36564 33658 36576
rect 33965 36567 34023 36573
rect 33965 36564 33977 36567
rect 33652 36536 33977 36564
rect 33652 36524 33658 36536
rect 33965 36533 33977 36536
rect 34011 36533 34023 36567
rect 33965 36527 34023 36533
rect 1104 36474 36892 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36892 36474
rect 1104 36400 36892 36422
rect 2225 36363 2283 36369
rect 2225 36329 2237 36363
rect 2271 36360 2283 36363
rect 2774 36360 2780 36372
rect 2271 36332 2780 36360
rect 2271 36329 2283 36332
rect 2225 36323 2283 36329
rect 1581 36159 1639 36165
rect 1581 36125 1593 36159
rect 1627 36156 1639 36159
rect 2240 36156 2268 36323
rect 2774 36320 2780 36332
rect 2832 36320 2838 36372
rect 36265 36363 36323 36369
rect 36265 36329 36277 36363
rect 36311 36360 36323 36363
rect 36722 36360 36728 36372
rect 36311 36332 36728 36360
rect 36311 36329 36323 36332
rect 36265 36323 36323 36329
rect 36722 36320 36728 36332
rect 36780 36320 36786 36372
rect 1627 36128 2268 36156
rect 1627 36125 1639 36128
rect 1581 36119 1639 36125
rect 32306 36116 32312 36168
rect 32364 36156 32370 36168
rect 36081 36159 36139 36165
rect 36081 36156 36093 36159
rect 32364 36128 36093 36156
rect 32364 36116 32370 36128
rect 36081 36125 36093 36128
rect 36127 36125 36139 36159
rect 36081 36119 36139 36125
rect 17586 36088 17592 36100
rect 1780 36060 17592 36088
rect 1780 36029 1808 36060
rect 17586 36048 17592 36060
rect 17644 36048 17650 36100
rect 1765 36023 1823 36029
rect 1765 35989 1777 36023
rect 1811 35989 1823 36023
rect 1765 35983 1823 35989
rect 1104 35930 36892 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 36892 35930
rect 1104 35856 36892 35878
rect 36078 35680 36084 35692
rect 36039 35652 36084 35680
rect 36078 35640 36084 35652
rect 36136 35640 36142 35692
rect 36262 35476 36268 35488
rect 36223 35448 36268 35476
rect 36262 35436 36268 35448
rect 36320 35436 36326 35488
rect 1104 35386 36892 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36892 35386
rect 1104 35312 36892 35334
rect 36078 35232 36084 35284
rect 36136 35272 36142 35284
rect 36173 35275 36231 35281
rect 36173 35272 36185 35275
rect 36136 35244 36185 35272
rect 36136 35232 36142 35244
rect 36173 35241 36185 35244
rect 36219 35241 36231 35275
rect 36173 35235 36231 35241
rect 1857 35071 1915 35077
rect 1857 35037 1869 35071
rect 1903 35068 1915 35071
rect 2682 35068 2688 35080
rect 1903 35040 2688 35068
rect 1903 35037 1915 35040
rect 1857 35031 1915 35037
rect 2682 35028 2688 35040
rect 2740 35028 2746 35080
rect 35989 35071 36047 35077
rect 35989 35068 36001 35071
rect 35866 35040 36001 35068
rect 1670 34932 1676 34944
rect 1631 34904 1676 34932
rect 1670 34892 1676 34904
rect 1728 34892 1734 34944
rect 35434 34932 35440 34944
rect 35395 34904 35440 34932
rect 35434 34892 35440 34904
rect 35492 34932 35498 34944
rect 35866 34932 35894 35040
rect 35989 35037 36001 35040
rect 36035 35037 36047 35071
rect 35989 35031 36047 35037
rect 35492 34904 35894 34932
rect 35492 34892 35498 34904
rect 1104 34842 36892 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 36892 34842
rect 1104 34768 36892 34790
rect 1104 34298 36892 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36892 34298
rect 1104 34224 36892 34246
rect 1104 33754 36892 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 36892 33754
rect 1104 33680 36892 33702
rect 35526 33464 35532 33516
rect 35584 33504 35590 33516
rect 36081 33507 36139 33513
rect 36081 33504 36093 33507
rect 35584 33476 36093 33504
rect 35584 33464 35590 33476
rect 36081 33473 36093 33476
rect 36127 33473 36139 33507
rect 36081 33467 36139 33473
rect 36262 33368 36268 33380
rect 36223 33340 36268 33368
rect 36262 33328 36268 33340
rect 36320 33328 36326 33380
rect 35526 33300 35532 33312
rect 35487 33272 35532 33300
rect 35526 33260 35532 33272
rect 35584 33260 35590 33312
rect 1104 33210 36892 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36892 33210
rect 1104 33136 36892 33158
rect 1670 32824 1676 32836
rect 1631 32796 1676 32824
rect 1670 32784 1676 32796
rect 1728 32784 1734 32836
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32756 1823 32759
rect 17862 32756 17868 32768
rect 1811 32728 17868 32756
rect 1811 32725 1823 32728
rect 1765 32719 1823 32725
rect 17862 32716 17868 32728
rect 17920 32716 17926 32768
rect 1104 32666 36892 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 36892 32666
rect 1104 32592 36892 32614
rect 1670 32552 1676 32564
rect 1631 32524 1676 32552
rect 1670 32512 1676 32524
rect 1728 32512 1734 32564
rect 1104 32122 36892 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36892 32122
rect 1104 32048 36892 32070
rect 3970 32008 3976 32020
rect 3931 31980 3976 32008
rect 3970 31968 3976 31980
rect 4028 31968 4034 32020
rect 36081 31875 36139 31881
rect 36081 31841 36093 31875
rect 36127 31872 36139 31875
rect 36446 31872 36452 31884
rect 36127 31844 36452 31872
rect 36127 31841 36139 31844
rect 36081 31835 36139 31841
rect 36446 31832 36452 31844
rect 36504 31832 36510 31884
rect 1854 31804 1860 31816
rect 1815 31776 1860 31804
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 4157 31807 4215 31813
rect 4157 31773 4169 31807
rect 4203 31804 4215 31807
rect 4614 31804 4620 31816
rect 4203 31776 4620 31804
rect 4203 31773 4215 31776
rect 4157 31767 4215 31773
rect 4614 31764 4620 31776
rect 4672 31764 4678 31816
rect 36354 31804 36360 31816
rect 36315 31776 36360 31804
rect 36354 31764 36360 31776
rect 36412 31764 36418 31816
rect 1670 31668 1676 31680
rect 1631 31640 1676 31668
rect 1670 31628 1676 31640
rect 1728 31628 1734 31680
rect 1104 31578 36892 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 36892 31578
rect 1104 31504 36892 31526
rect 1854 31424 1860 31476
rect 1912 31464 1918 31476
rect 1949 31467 2007 31473
rect 1949 31464 1961 31467
rect 1912 31436 1961 31464
rect 1912 31424 1918 31436
rect 1949 31433 1961 31436
rect 1995 31433 2007 31467
rect 1949 31427 2007 31433
rect 23382 31424 23388 31476
rect 23440 31464 23446 31476
rect 23569 31467 23627 31473
rect 23569 31464 23581 31467
rect 23440 31436 23581 31464
rect 23440 31424 23446 31436
rect 23569 31433 23581 31436
rect 23615 31433 23627 31467
rect 23569 31427 23627 31433
rect 27617 31467 27675 31473
rect 27617 31433 27629 31467
rect 27663 31464 27675 31467
rect 32306 31464 32312 31476
rect 27663 31436 32312 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 32306 31424 32312 31436
rect 32364 31424 32370 31476
rect 2038 31328 2044 31340
rect 1999 31300 2044 31328
rect 2038 31288 2044 31300
rect 2096 31328 2102 31340
rect 2501 31331 2559 31337
rect 2501 31328 2513 31331
rect 2096 31300 2513 31328
rect 2096 31288 2102 31300
rect 2501 31297 2513 31300
rect 2547 31297 2559 31331
rect 2501 31291 2559 31297
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19797 31331 19855 31337
rect 19797 31328 19809 31331
rect 19484 31300 19809 31328
rect 19484 31288 19490 31300
rect 19797 31297 19809 31300
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 22925 31331 22983 31337
rect 22925 31297 22937 31331
rect 22971 31328 22983 31331
rect 23400 31328 23428 31424
rect 36354 31396 36360 31408
rect 36315 31368 36360 31396
rect 36354 31356 36360 31368
rect 36412 31356 36418 31408
rect 27430 31328 27436 31340
rect 22971 31300 23428 31328
rect 27391 31300 27436 31328
rect 22971 31297 22983 31300
rect 22925 31291 22983 31297
rect 27430 31288 27436 31300
rect 27488 31328 27494 31340
rect 28077 31331 28135 31337
rect 28077 31328 28089 31331
rect 27488 31300 28089 31328
rect 27488 31288 27494 31300
rect 28077 31297 28089 31300
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 19889 31127 19947 31133
rect 19889 31093 19901 31127
rect 19935 31124 19947 31127
rect 19978 31124 19984 31136
rect 19935 31096 19984 31124
rect 19935 31093 19947 31096
rect 19889 31087 19947 31093
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 23014 31124 23020 31136
rect 22975 31096 23020 31124
rect 23014 31084 23020 31096
rect 23072 31084 23078 31136
rect 1104 31034 36892 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36892 31034
rect 1104 30960 36892 30982
rect 1762 30920 1768 30932
rect 1723 30892 1768 30920
rect 1762 30880 1768 30892
rect 1820 30880 1826 30932
rect 1854 30676 1860 30728
rect 1912 30716 1918 30728
rect 1949 30719 2007 30725
rect 1949 30716 1961 30719
rect 1912 30688 1961 30716
rect 1912 30676 1918 30688
rect 1949 30685 1961 30688
rect 1995 30685 2007 30719
rect 1949 30679 2007 30685
rect 1104 30490 36892 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 36892 30490
rect 1104 30416 36892 30438
rect 35618 30200 35624 30252
rect 35676 30240 35682 30252
rect 36081 30243 36139 30249
rect 36081 30240 36093 30243
rect 35676 30212 36093 30240
rect 35676 30200 35682 30212
rect 36081 30209 36093 30212
rect 36127 30209 36139 30243
rect 36081 30203 36139 30209
rect 35618 30036 35624 30048
rect 35579 30008 35624 30036
rect 35618 29996 35624 30008
rect 35676 29996 35682 30048
rect 36262 30036 36268 30048
rect 36223 30008 36268 30036
rect 36262 29996 36268 30008
rect 36320 29996 36326 30048
rect 1104 29946 36892 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36892 29946
rect 1104 29872 36892 29894
rect 2682 29792 2688 29844
rect 2740 29832 2746 29844
rect 5997 29835 6055 29841
rect 5997 29832 6009 29835
rect 2740 29804 6009 29832
rect 2740 29792 2746 29804
rect 5997 29801 6009 29804
rect 6043 29801 6055 29835
rect 5997 29795 6055 29801
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29628 1915 29631
rect 1946 29628 1952 29640
rect 1903 29600 1952 29628
rect 1903 29597 1915 29600
rect 1857 29591 1915 29597
rect 1946 29588 1952 29600
rect 2004 29588 2010 29640
rect 6086 29628 6092 29640
rect 6047 29600 6092 29628
rect 6086 29588 6092 29600
rect 6144 29628 6150 29640
rect 6549 29631 6607 29637
rect 6549 29628 6561 29631
rect 6144 29600 6561 29628
rect 6144 29588 6150 29600
rect 6549 29597 6561 29600
rect 6595 29597 6607 29631
rect 6549 29591 6607 29597
rect 11054 29588 11060 29640
rect 11112 29628 11118 29640
rect 11977 29631 12035 29637
rect 11977 29628 11989 29631
rect 11112 29600 11989 29628
rect 11112 29588 11118 29600
rect 11977 29597 11989 29600
rect 12023 29597 12035 29631
rect 11977 29591 12035 29597
rect 1670 29492 1676 29504
rect 1631 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29452 1734 29504
rect 12069 29495 12127 29501
rect 12069 29461 12081 29495
rect 12115 29492 12127 29495
rect 17218 29492 17224 29504
rect 12115 29464 17224 29492
rect 12115 29461 12127 29464
rect 12069 29455 12127 29461
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 1104 29402 36892 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 36892 29402
rect 1104 29328 36892 29350
rect 1104 28858 36892 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36892 28858
rect 1104 28784 36892 28806
rect 1104 28314 36892 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 36892 28314
rect 1104 28240 36892 28262
rect 35621 28067 35679 28073
rect 35621 28033 35633 28067
rect 35667 28064 35679 28067
rect 36262 28064 36268 28076
rect 35667 28036 36268 28064
rect 35667 28033 35679 28036
rect 35621 28027 35679 28033
rect 36262 28024 36268 28036
rect 36320 28024 36326 28076
rect 36170 27860 36176 27872
rect 36131 27832 36176 27860
rect 36170 27820 36176 27832
rect 36228 27820 36234 27872
rect 1104 27770 36892 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36892 27770
rect 1104 27696 36892 27718
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27452 1915 27455
rect 3694 27452 3700 27464
rect 1903 27424 3700 27452
rect 1903 27421 1915 27424
rect 1857 27415 1915 27421
rect 3694 27412 3700 27424
rect 3752 27412 3758 27464
rect 1670 27316 1676 27328
rect 1631 27288 1676 27316
rect 1670 27276 1676 27288
rect 1728 27276 1734 27328
rect 1104 27226 36892 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 36892 27226
rect 1104 27152 36892 27174
rect 1104 26682 36892 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36892 26682
rect 1104 26608 36892 26630
rect 26786 26568 26792 26580
rect 26747 26540 26792 26568
rect 26786 26528 26792 26540
rect 26844 26528 26850 26580
rect 35802 26460 35808 26512
rect 35860 26500 35866 26512
rect 36265 26503 36323 26509
rect 36265 26500 36277 26503
rect 35860 26472 36277 26500
rect 35860 26460 35866 26472
rect 36265 26469 36277 26472
rect 36311 26469 36323 26503
rect 36265 26463 36323 26469
rect 26605 26367 26663 26373
rect 26605 26333 26617 26367
rect 26651 26364 26663 26367
rect 26651 26336 27384 26364
rect 26651 26333 26663 26336
rect 26605 26327 26663 26333
rect 27356 26305 27384 26336
rect 35342 26324 35348 26376
rect 35400 26364 35406 26376
rect 36081 26367 36139 26373
rect 36081 26364 36093 26367
rect 35400 26336 36093 26364
rect 35400 26324 35406 26336
rect 36081 26333 36093 26336
rect 36127 26333 36139 26367
rect 36081 26327 36139 26333
rect 27341 26299 27399 26305
rect 27341 26265 27353 26299
rect 27387 26296 27399 26299
rect 27614 26296 27620 26308
rect 27387 26268 27620 26296
rect 27387 26265 27399 26268
rect 27341 26259 27399 26265
rect 27614 26256 27620 26268
rect 27672 26256 27678 26308
rect 1104 26138 36892 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 36892 26138
rect 1104 26064 36892 26086
rect 1104 25594 36892 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36892 25594
rect 1104 25520 36892 25542
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 1854 25276 1860 25288
rect 1815 25248 1860 25276
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 1104 25050 36892 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 36892 25050
rect 1104 24976 36892 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 1104 24506 36892 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36892 24506
rect 1104 24432 36892 24454
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 4614 24188 4620 24200
rect 1903 24160 4620 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 36081 24191 36139 24197
rect 36081 24188 36093 24191
rect 30432 24160 36093 24188
rect 30432 24148 30438 24160
rect 36081 24157 36093 24160
rect 36127 24157 36139 24191
rect 36354 24188 36360 24200
rect 36315 24160 36360 24188
rect 36081 24151 36139 24157
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 1104 23962 36892 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 36892 23962
rect 1104 23888 36892 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 7285 23851 7343 23857
rect 7285 23848 7297 23851
rect 6886 23820 7297 23848
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23712 6791 23715
rect 6886 23712 6914 23820
rect 7285 23817 7297 23820
rect 7331 23848 7343 23851
rect 8938 23848 8944 23860
rect 7331 23820 8944 23848
rect 7331 23817 7343 23820
rect 7285 23811 7343 23817
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 36354 23848 36360 23860
rect 36315 23820 36360 23848
rect 36354 23808 36360 23820
rect 36412 23808 36418 23860
rect 6779 23684 6914 23712
rect 12253 23715 12311 23721
rect 6779 23681 6791 23684
rect 6733 23675 6791 23681
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 12710 23712 12716 23724
rect 12299 23684 12716 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 1946 23536 1952 23588
rect 2004 23576 2010 23588
rect 12069 23579 12127 23585
rect 12069 23576 12081 23579
rect 2004 23548 12081 23576
rect 2004 23536 2010 23548
rect 12069 23545 12081 23548
rect 12115 23545 12127 23579
rect 12069 23539 12127 23545
rect 6546 23508 6552 23520
rect 6507 23480 6552 23508
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 12710 23508 12716 23520
rect 12671 23480 12716 23508
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 1104 23418 36892 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36892 23418
rect 1104 23344 36892 23366
rect 3694 23264 3700 23316
rect 3752 23304 3758 23316
rect 4709 23307 4767 23313
rect 4709 23304 4721 23307
rect 3752 23276 4721 23304
rect 3752 23264 3758 23276
rect 4709 23273 4721 23276
rect 4755 23273 4767 23307
rect 4709 23267 4767 23273
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23100 4951 23103
rect 4939 23072 5488 23100
rect 4939 23069 4951 23072
rect 4893 23063 4951 23069
rect 5460 22973 5488 23072
rect 5445 22967 5503 22973
rect 5445 22933 5457 22967
rect 5491 22964 5503 22967
rect 13262 22964 13268 22976
rect 5491 22936 13268 22964
rect 5491 22933 5503 22936
rect 5445 22927 5503 22933
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 1104 22874 36892 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 36892 22874
rect 1104 22800 36892 22822
rect 36078 22624 36084 22636
rect 36039 22596 36084 22624
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 36262 22488 36268 22500
rect 36223 22460 36268 22488
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 1104 22330 36892 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36892 22330
rect 1104 22256 36892 22278
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 1765 21879 1823 21885
rect 1765 21845 1777 21879
rect 1811 21876 1823 21879
rect 24578 21876 24584 21888
rect 1811 21848 24584 21876
rect 1811 21845 1823 21848
rect 1765 21839 1823 21845
rect 24578 21836 24584 21848
rect 24636 21876 24642 21888
rect 27430 21876 27436 21888
rect 24636 21848 27436 21876
rect 24636 21836 24642 21848
rect 27430 21836 27436 21848
rect 27488 21836 27494 21888
rect 1104 21786 36892 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 36892 21786
rect 1104 21712 36892 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21536 19027 21539
rect 19015 21508 19656 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 2314 21292 2320 21344
rect 2372 21332 2378 21344
rect 19628 21341 19656 21508
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 2372 21304 18889 21332
rect 2372 21292 2378 21304
rect 18877 21301 18889 21304
rect 18923 21301 18935 21335
rect 18877 21295 18935 21301
rect 19613 21335 19671 21341
rect 19613 21301 19625 21335
rect 19659 21332 19671 21335
rect 35710 21332 35716 21344
rect 19659 21304 35716 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 35710 21292 35716 21304
rect 35768 21292 35774 21344
rect 1104 21242 36892 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36892 21242
rect 1104 21168 36892 21190
rect 35621 21131 35679 21137
rect 35621 21097 35633 21131
rect 35667 21128 35679 21131
rect 35986 21128 35992 21140
rect 35667 21100 35992 21128
rect 35667 21097 35679 21100
rect 35621 21091 35679 21097
rect 35986 21088 35992 21100
rect 36044 21088 36050 21140
rect 4614 20952 4620 21004
rect 4672 20992 4678 21004
rect 4672 20964 9168 20992
rect 4672 20952 4678 20964
rect 1854 20884 1860 20936
rect 1912 20924 1918 20936
rect 9140 20933 9168 20964
rect 8389 20927 8447 20933
rect 8389 20924 8401 20927
rect 1912 20896 8401 20924
rect 1912 20884 1918 20896
rect 8389 20893 8401 20896
rect 8435 20893 8447 20927
rect 8389 20887 8447 20893
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20924 9183 20927
rect 9769 20927 9827 20933
rect 9769 20924 9781 20927
rect 9171 20896 9781 20924
rect 9171 20893 9183 20896
rect 9125 20887 9183 20893
rect 9769 20893 9781 20896
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 35437 20927 35495 20933
rect 35437 20893 35449 20927
rect 35483 20924 35495 20927
rect 35710 20924 35716 20936
rect 35483 20896 35716 20924
rect 35483 20893 35495 20896
rect 35437 20887 35495 20893
rect 35710 20884 35716 20896
rect 35768 20884 35774 20936
rect 36081 20927 36139 20933
rect 36081 20924 36093 20927
rect 35866 20896 36093 20924
rect 8481 20859 8539 20865
rect 8481 20825 8493 20859
rect 8527 20856 8539 20859
rect 17954 20856 17960 20868
rect 8527 20828 17960 20856
rect 8527 20825 8539 20828
rect 8481 20819 8539 20825
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 33134 20816 33140 20868
rect 33192 20856 33198 20868
rect 35866 20856 35894 20896
rect 36081 20893 36093 20896
rect 36127 20893 36139 20927
rect 36081 20887 36139 20893
rect 33192 20828 35894 20856
rect 33192 20816 33198 20828
rect 9214 20788 9220 20800
rect 9175 20760 9220 20788
rect 9214 20748 9220 20760
rect 9272 20748 9278 20800
rect 36262 20788 36268 20800
rect 36223 20760 36268 20788
rect 36262 20748 36268 20760
rect 36320 20748 36326 20800
rect 1104 20698 36892 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 36892 20698
rect 1104 20624 36892 20646
rect 35710 20244 35716 20256
rect 35671 20216 35716 20244
rect 35710 20204 35716 20216
rect 35768 20204 35774 20256
rect 1104 20154 36892 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36892 20154
rect 1104 20080 36892 20102
rect 29917 20043 29975 20049
rect 29917 20009 29929 20043
rect 29963 20040 29975 20043
rect 33134 20040 33140 20052
rect 29963 20012 33140 20040
rect 29963 20009 29975 20012
rect 29917 20003 29975 20009
rect 33134 20000 33140 20012
rect 33192 20000 33198 20052
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19836 1915 19839
rect 21358 19836 21364 19848
rect 1903 19808 21364 19836
rect 1903 19805 1915 19808
rect 1857 19799 1915 19805
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 29730 19836 29736 19848
rect 29691 19808 29736 19836
rect 29730 19796 29736 19808
rect 29788 19836 29794 19848
rect 30377 19839 30435 19845
rect 30377 19836 30389 19839
rect 29788 19808 30389 19836
rect 29788 19796 29794 19808
rect 30377 19805 30389 19808
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 1104 19610 36892 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 36892 19610
rect 1104 19536 36892 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 34885 19499 34943 19505
rect 34885 19465 34897 19499
rect 34931 19496 34943 19499
rect 36078 19496 36084 19508
rect 34931 19468 36084 19496
rect 34931 19465 34943 19468
rect 34885 19459 34943 19465
rect 36078 19456 36084 19468
rect 36136 19456 36142 19508
rect 34606 19320 34612 19372
rect 34664 19360 34670 19372
rect 34701 19363 34759 19369
rect 34701 19360 34713 19363
rect 34664 19332 34713 19360
rect 34664 19320 34670 19332
rect 34701 19329 34713 19332
rect 34747 19360 34759 19363
rect 35345 19363 35403 19369
rect 35345 19360 35357 19363
rect 34747 19332 35357 19360
rect 34747 19329 34759 19332
rect 34701 19323 34759 19329
rect 35345 19329 35357 19332
rect 35391 19329 35403 19363
rect 35345 19323 35403 19329
rect 1104 19066 36892 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36892 19066
rect 1104 18992 36892 19014
rect 31021 18955 31079 18961
rect 31021 18921 31033 18955
rect 31067 18952 31079 18955
rect 35342 18952 35348 18964
rect 31067 18924 35348 18952
rect 31067 18921 31079 18924
rect 31021 18915 31079 18921
rect 35342 18912 35348 18924
rect 35400 18912 35406 18964
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 30929 18751 30987 18757
rect 30929 18748 30941 18751
rect 28592 18720 30941 18748
rect 28592 18708 28598 18720
rect 30929 18717 30941 18720
rect 30975 18717 30987 18751
rect 30929 18711 30987 18717
rect 34514 18708 34520 18760
rect 34572 18748 34578 18760
rect 36081 18751 36139 18757
rect 36081 18748 36093 18751
rect 34572 18720 36093 18748
rect 34572 18708 34578 18720
rect 36081 18717 36093 18720
rect 36127 18717 36139 18751
rect 36081 18711 36139 18717
rect 1578 18640 1584 18692
rect 1636 18680 1642 18692
rect 1673 18683 1731 18689
rect 1673 18680 1685 18683
rect 1636 18652 1685 18680
rect 1636 18640 1642 18652
rect 1673 18649 1685 18652
rect 1719 18649 1731 18683
rect 1673 18643 1731 18649
rect 1857 18683 1915 18689
rect 1857 18649 1869 18683
rect 1903 18680 1915 18683
rect 2682 18680 2688 18692
rect 1903 18652 2688 18680
rect 1903 18649 1915 18652
rect 1857 18643 1915 18649
rect 2682 18640 2688 18652
rect 2740 18640 2746 18692
rect 23566 18612 23572 18624
rect 23527 18584 23572 18612
rect 23566 18572 23572 18584
rect 23624 18572 23630 18624
rect 36262 18612 36268 18624
rect 36223 18584 36268 18612
rect 36262 18572 36268 18584
rect 36320 18572 36326 18624
rect 1104 18522 36892 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 36892 18522
rect 1104 18448 36892 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 24578 18408 24584 18420
rect 24539 18380 24584 18408
rect 24578 18368 24584 18380
rect 24636 18368 24642 18420
rect 26145 18275 26203 18281
rect 26145 18241 26157 18275
rect 26191 18272 26203 18275
rect 27341 18275 27399 18281
rect 27341 18272 27353 18275
rect 26191 18244 27353 18272
rect 26191 18241 26203 18244
rect 26145 18235 26203 18241
rect 27341 18241 27353 18244
rect 27387 18272 27399 18275
rect 30374 18272 30380 18284
rect 27387 18244 30380 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 22833 18207 22891 18213
rect 22833 18173 22845 18207
rect 22879 18204 22891 18207
rect 23106 18204 23112 18216
rect 22879 18176 23112 18204
rect 22879 18173 22891 18176
rect 22833 18167 22891 18173
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 25682 18096 25688 18148
rect 25740 18136 25746 18148
rect 25961 18139 26019 18145
rect 25961 18136 25973 18139
rect 25740 18108 25973 18136
rect 25740 18096 25746 18108
rect 25961 18105 25973 18108
rect 26007 18105 26019 18139
rect 25961 18099 26019 18105
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 22002 18068 22008 18080
rect 5592 18040 22008 18068
rect 5592 18028 5598 18040
rect 22002 18028 22008 18040
rect 22060 18068 22066 18080
rect 22097 18071 22155 18077
rect 22097 18068 22109 18071
rect 22060 18040 22109 18068
rect 22060 18028 22066 18040
rect 22097 18037 22109 18040
rect 22143 18037 22155 18071
rect 22097 18031 22155 18037
rect 22830 18028 22836 18080
rect 22888 18068 22894 18080
rect 23293 18071 23351 18077
rect 23293 18068 23305 18071
rect 22888 18040 23305 18068
rect 22888 18028 22894 18040
rect 23293 18037 23305 18040
rect 23339 18037 23351 18071
rect 23293 18031 23351 18037
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 24029 18071 24087 18077
rect 24029 18068 24041 18071
rect 23900 18040 24041 18068
rect 23900 18028 23906 18040
rect 24029 18037 24041 18040
rect 24075 18068 24087 18071
rect 24762 18068 24768 18080
rect 24075 18040 24768 18068
rect 24075 18037 24087 18040
rect 24029 18031 24087 18037
rect 24762 18028 24768 18040
rect 24820 18068 24826 18080
rect 25041 18071 25099 18077
rect 25041 18068 25053 18071
rect 24820 18040 25053 18068
rect 24820 18028 24826 18040
rect 25041 18037 25053 18040
rect 25087 18037 25099 18071
rect 25041 18031 25099 18037
rect 26694 18028 26700 18080
rect 26752 18068 26758 18080
rect 27249 18071 27307 18077
rect 27249 18068 27261 18071
rect 26752 18040 27261 18068
rect 26752 18028 26758 18040
rect 27249 18037 27261 18040
rect 27295 18037 27307 18071
rect 27249 18031 27307 18037
rect 1104 17978 36892 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36892 17978
rect 1104 17904 36892 17926
rect 21358 17864 21364 17876
rect 21319 17836 21364 17864
rect 21358 17824 21364 17836
rect 21416 17864 21422 17876
rect 21913 17867 21971 17873
rect 21913 17864 21925 17867
rect 21416 17836 21925 17864
rect 21416 17824 21422 17836
rect 21913 17833 21925 17836
rect 21959 17833 21971 17867
rect 21913 17827 21971 17833
rect 33229 17867 33287 17873
rect 33229 17833 33241 17867
rect 33275 17864 33287 17867
rect 34514 17864 34520 17876
rect 33275 17836 34520 17864
rect 33275 17833 33287 17836
rect 33229 17827 33287 17833
rect 34514 17824 34520 17836
rect 34572 17824 34578 17876
rect 23198 17796 23204 17808
rect 22848 17768 23204 17796
rect 22848 17737 22876 17768
rect 23198 17756 23204 17768
rect 23256 17756 23262 17808
rect 22833 17731 22891 17737
rect 22833 17697 22845 17731
rect 22879 17697 22891 17731
rect 23106 17728 23112 17740
rect 23067 17700 23112 17728
rect 22833 17691 22891 17697
rect 23106 17688 23112 17700
rect 23164 17688 23170 17740
rect 23842 17660 23848 17672
rect 23803 17632 23848 17660
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 24578 17620 24584 17672
rect 24636 17660 24642 17672
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24636 17632 24685 17660
rect 24636 17620 24642 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 25498 17660 25504 17672
rect 25459 17632 25504 17660
rect 24673 17623 24731 17629
rect 25498 17620 25504 17632
rect 25556 17660 25562 17672
rect 25961 17663 26019 17669
rect 25961 17660 25973 17663
rect 25556 17632 25973 17660
rect 25556 17620 25562 17632
rect 25961 17629 25973 17632
rect 26007 17660 26019 17663
rect 29730 17660 29736 17672
rect 26007 17632 29736 17660
rect 26007 17629 26019 17632
rect 25961 17623 26019 17629
rect 29730 17620 29736 17632
rect 29788 17620 29794 17672
rect 33137 17663 33195 17669
rect 33137 17660 33149 17663
rect 31726 17632 33149 17660
rect 23017 17595 23075 17601
rect 23017 17561 23029 17595
rect 23063 17561 23075 17595
rect 23017 17555 23075 17561
rect 20898 17524 20904 17536
rect 20859 17496 20904 17524
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 23032 17524 23060 17555
rect 27798 17552 27804 17604
rect 27856 17592 27862 17604
rect 31726 17592 31754 17632
rect 33137 17629 33149 17632
rect 33183 17629 33195 17663
rect 33137 17623 33195 17629
rect 27856 17564 31754 17592
rect 27856 17552 27862 17564
rect 23753 17527 23811 17533
rect 23753 17524 23765 17527
rect 23032 17496 23765 17524
rect 23753 17493 23765 17496
rect 23799 17493 23811 17527
rect 23753 17487 23811 17493
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24636 17496 24685 17524
rect 24636 17484 24642 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24673 17487 24731 17493
rect 25409 17527 25467 17533
rect 25409 17493 25421 17527
rect 25455 17524 25467 17527
rect 25866 17524 25872 17536
rect 25455 17496 25872 17524
rect 25455 17493 25467 17496
rect 25409 17487 25467 17493
rect 25866 17484 25872 17496
rect 25924 17484 25930 17536
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 26513 17527 26571 17533
rect 26513 17524 26525 17527
rect 26200 17496 26525 17524
rect 26200 17484 26206 17496
rect 26513 17493 26525 17496
rect 26559 17493 26571 17527
rect 26513 17487 26571 17493
rect 1104 17434 36892 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 36892 17434
rect 1104 17360 36892 17382
rect 25225 17323 25283 17329
rect 25225 17320 25237 17323
rect 24504 17292 25237 17320
rect 24504 17261 24532 17292
rect 25225 17289 25237 17292
rect 25271 17289 25283 17323
rect 25225 17283 25283 17289
rect 24489 17255 24547 17261
rect 24489 17221 24501 17255
rect 24535 17221 24547 17255
rect 24489 17215 24547 17221
rect 24578 17212 24584 17264
rect 24636 17252 24642 17264
rect 27430 17252 27436 17264
rect 24636 17224 24681 17252
rect 25332 17224 27436 17252
rect 24636 17212 24642 17224
rect 20533 17187 20591 17193
rect 20533 17153 20545 17187
rect 20579 17153 20591 17187
rect 20533 17147 20591 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 21358 17184 21364 17196
rect 21315 17156 21364 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 20548 17116 20576 17147
rect 21358 17144 21364 17156
rect 21416 17184 21422 17196
rect 22097 17187 22155 17193
rect 22097 17184 22109 17187
rect 21416 17156 22109 17184
rect 21416 17144 21422 17156
rect 22097 17153 22109 17156
rect 22143 17153 22155 17187
rect 22830 17184 22836 17196
rect 22791 17156 22836 17184
rect 22097 17147 22155 17153
rect 22830 17144 22836 17156
rect 22888 17144 22894 17196
rect 25332 17193 25360 17224
rect 27430 17212 27436 17224
rect 27488 17212 27494 17264
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 26142 17184 26148 17196
rect 25464 17156 26148 17184
rect 25464 17144 25470 17156
rect 26142 17144 26148 17156
rect 26200 17184 26206 17196
rect 26421 17187 26479 17193
rect 26421 17184 26433 17187
rect 26200 17156 26433 17184
rect 26200 17144 26206 17156
rect 26421 17153 26433 17156
rect 26467 17153 26479 17187
rect 36078 17184 36084 17196
rect 36039 17156 36084 17184
rect 26421 17147 26479 17153
rect 36078 17144 36084 17156
rect 36136 17144 36142 17196
rect 20898 17116 20904 17128
rect 20548 17088 20904 17116
rect 20898 17076 20904 17088
rect 20956 17116 20962 17128
rect 21634 17116 21640 17128
rect 20956 17088 21640 17116
rect 20956 17076 20962 17088
rect 21634 17076 21640 17088
rect 21692 17076 21698 17128
rect 22281 17119 22339 17125
rect 22281 17085 22293 17119
rect 22327 17116 22339 17119
rect 25774 17116 25780 17128
rect 22327 17088 25636 17116
rect 25735 17088 25780 17116
rect 22327 17085 22339 17088
rect 22281 17079 22339 17085
rect 23198 17008 23204 17060
rect 23256 17048 23262 17060
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 23256 17020 24041 17048
rect 23256 17008 23262 17020
rect 24029 17017 24041 17020
rect 24075 17017 24087 17051
rect 25608 17048 25636 17088
rect 25774 17076 25780 17088
rect 25832 17076 25838 17128
rect 35618 17116 35624 17128
rect 26344 17088 35624 17116
rect 26234 17048 26240 17060
rect 25608 17020 26240 17048
rect 24029 17011 24087 17017
rect 26234 17008 26240 17020
rect 26292 17008 26298 17060
rect 20625 16983 20683 16989
rect 20625 16949 20637 16983
rect 20671 16980 20683 16983
rect 20990 16980 20996 16992
rect 20671 16952 20996 16980
rect 20671 16949 20683 16952
rect 20625 16943 20683 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21358 16980 21364 16992
rect 21319 16952 21364 16980
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 22925 16983 22983 16989
rect 22925 16949 22937 16983
rect 22971 16980 22983 16983
rect 26344 16980 26372 17088
rect 35618 17076 35624 17088
rect 35676 17076 35682 17128
rect 26418 17008 26424 17060
rect 26476 17048 26482 17060
rect 35526 17048 35532 17060
rect 26476 17020 35532 17048
rect 26476 17008 26482 17020
rect 35526 17008 35532 17020
rect 35584 17008 35590 17060
rect 36262 17048 36268 17060
rect 36223 17020 36268 17048
rect 36262 17008 36268 17020
rect 36320 17008 36326 17060
rect 22971 16952 26372 16980
rect 26513 16983 26571 16989
rect 22971 16949 22983 16952
rect 22925 16943 22983 16949
rect 26513 16949 26525 16983
rect 26559 16980 26571 16983
rect 26602 16980 26608 16992
rect 26559 16952 26608 16980
rect 26559 16949 26571 16952
rect 26513 16943 26571 16949
rect 26602 16940 26608 16952
rect 26660 16940 26666 16992
rect 1104 16890 36892 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36892 16890
rect 1104 16816 36892 16838
rect 25406 16776 25412 16788
rect 22066 16748 25412 16776
rect 22066 16708 22094 16748
rect 25406 16736 25412 16748
rect 25464 16736 25470 16788
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 27893 16779 27951 16785
rect 27893 16776 27905 16779
rect 27672 16748 27905 16776
rect 27672 16736 27678 16748
rect 27893 16745 27905 16748
rect 27939 16745 27951 16779
rect 27893 16739 27951 16745
rect 27522 16708 27528 16720
rect 20272 16680 22094 16708
rect 25424 16680 27528 16708
rect 19613 16643 19671 16649
rect 19613 16609 19625 16643
rect 19659 16640 19671 16643
rect 20272 16640 20300 16680
rect 20714 16640 20720 16652
rect 19659 16612 20300 16640
rect 20675 16612 20720 16640
rect 19659 16609 19671 16612
rect 19613 16603 19671 16609
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 11698 16572 11704 16584
rect 1903 16544 11704 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 20272 16581 20300 16612
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 22557 16643 22615 16649
rect 22557 16640 22569 16643
rect 21416 16612 22569 16640
rect 21416 16600 21422 16612
rect 22557 16609 22569 16612
rect 22603 16609 22615 16643
rect 22557 16603 22615 16609
rect 22741 16643 22799 16649
rect 22741 16609 22753 16643
rect 22787 16640 22799 16643
rect 24673 16643 24731 16649
rect 24673 16640 24685 16643
rect 22787 16612 24685 16640
rect 22787 16609 22799 16612
rect 22741 16603 22799 16609
rect 24673 16609 24685 16612
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16572 21051 16575
rect 21039 16544 21956 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 21818 16504 21824 16516
rect 21779 16476 21824 16504
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 21928 16504 21956 16544
rect 22002 16532 22008 16584
rect 22060 16572 22066 16584
rect 23566 16572 23572 16584
rect 22060 16544 23572 16572
rect 22060 16532 22066 16544
rect 23566 16532 23572 16544
rect 23624 16572 23630 16584
rect 23661 16575 23719 16581
rect 23661 16572 23673 16575
rect 23624 16544 23673 16572
rect 23624 16532 23630 16544
rect 23661 16541 23673 16544
rect 23707 16541 23719 16575
rect 24762 16572 24768 16584
rect 24675 16544 24768 16572
rect 23661 16535 23719 16541
rect 24762 16532 24768 16544
rect 24820 16532 24826 16584
rect 25424 16581 25452 16680
rect 27522 16668 27528 16680
rect 27580 16668 27586 16720
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 26237 16643 26295 16649
rect 26237 16640 26249 16643
rect 26108 16612 26249 16640
rect 26108 16600 26114 16612
rect 26237 16609 26249 16612
rect 26283 16609 26295 16643
rect 26694 16640 26700 16652
rect 26655 16612 26700 16640
rect 26237 16603 26295 16609
rect 26694 16600 26700 16612
rect 26752 16600 26758 16652
rect 28994 16640 29000 16652
rect 28966 16600 29000 16640
rect 29052 16600 29058 16652
rect 25409 16575 25467 16581
rect 25409 16541 25421 16575
rect 25455 16541 25467 16575
rect 27430 16572 27436 16584
rect 27391 16544 27436 16572
rect 25409 16535 25467 16541
rect 27430 16532 27436 16544
rect 27488 16572 27494 16584
rect 28966 16572 28994 16600
rect 27488 16544 28994 16572
rect 27488 16532 27494 16544
rect 22094 16504 22100 16516
rect 21928 16476 22100 16504
rect 22094 16464 22100 16476
rect 22152 16504 22158 16516
rect 22646 16504 22652 16516
rect 22152 16476 22652 16504
rect 22152 16464 22158 16476
rect 22646 16464 22652 16476
rect 22704 16464 22710 16516
rect 24780 16504 24808 16532
rect 26326 16504 26332 16516
rect 24780 16476 26332 16504
rect 26326 16464 26332 16476
rect 26384 16464 26390 16516
rect 26602 16504 26608 16516
rect 26563 16476 26608 16504
rect 26602 16464 26608 16476
rect 26660 16464 26666 16516
rect 27154 16464 27160 16516
rect 27212 16504 27218 16516
rect 27798 16504 27804 16516
rect 27212 16476 27804 16504
rect 27212 16464 27218 16476
rect 27798 16464 27804 16476
rect 27856 16504 27862 16516
rect 28166 16504 28172 16516
rect 27856 16476 28172 16504
rect 27856 16464 27862 16476
rect 28166 16464 28172 16476
rect 28224 16464 28230 16516
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 20162 16436 20168 16448
rect 20123 16408 20168 16436
rect 20162 16396 20168 16408
rect 20220 16396 20226 16448
rect 21910 16436 21916 16448
rect 21871 16408 21916 16436
rect 21910 16396 21916 16408
rect 21968 16396 21974 16448
rect 23201 16439 23259 16445
rect 23201 16405 23213 16439
rect 23247 16436 23259 16439
rect 23474 16436 23480 16448
rect 23247 16408 23480 16436
rect 23247 16405 23259 16408
rect 23201 16399 23259 16405
rect 23474 16396 23480 16408
rect 23532 16396 23538 16448
rect 23842 16436 23848 16448
rect 23803 16408 23848 16436
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25317 16439 25375 16445
rect 25317 16436 25329 16439
rect 24912 16408 25329 16436
rect 24912 16396 24918 16408
rect 25317 16405 25329 16408
rect 25363 16405 25375 16439
rect 25317 16399 25375 16405
rect 26142 16396 26148 16448
rect 26200 16436 26206 16448
rect 27341 16439 27399 16445
rect 27341 16436 27353 16439
rect 26200 16408 27353 16436
rect 26200 16396 26206 16408
rect 27341 16405 27353 16408
rect 27387 16405 27399 16439
rect 27341 16399 27399 16405
rect 1104 16346 36892 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 36892 16346
rect 1104 16272 36892 16294
rect 11698 16232 11704 16244
rect 11659 16204 11704 16232
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 17276 16204 19073 16232
rect 17276 16192 17282 16204
rect 19061 16201 19073 16204
rect 19107 16232 19119 16235
rect 19334 16232 19340 16244
rect 19107 16204 19340 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 21453 16235 21511 16241
rect 21453 16201 21465 16235
rect 21499 16232 21511 16235
rect 22094 16232 22100 16244
rect 21499 16204 22100 16232
rect 21499 16201 21511 16204
rect 21453 16195 21511 16201
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 27338 16232 27344 16244
rect 22204 16204 23612 16232
rect 9214 16124 9220 16176
rect 9272 16164 9278 16176
rect 9272 16136 20300 16164
rect 9272 16124 9278 16136
rect 20272 16105 20300 16136
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 11931 16068 12449 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16065 20315 16099
rect 22204 16096 22232 16204
rect 22554 16164 22560 16176
rect 22515 16136 22560 16164
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 23584 16105 23612 16204
rect 24964 16204 27344 16232
rect 24964 16173 24992 16204
rect 27338 16192 27344 16204
rect 27396 16192 27402 16244
rect 24949 16167 25007 16173
rect 24949 16133 24961 16167
rect 24995 16133 25007 16167
rect 24949 16127 25007 16133
rect 25041 16167 25099 16173
rect 25041 16133 25053 16167
rect 25087 16164 25099 16167
rect 25774 16164 25780 16176
rect 25087 16136 25780 16164
rect 25087 16133 25099 16136
rect 25041 16127 25099 16133
rect 25774 16124 25780 16136
rect 25832 16124 25838 16176
rect 26786 16124 26792 16176
rect 26844 16164 26850 16176
rect 26844 16136 27660 16164
rect 26844 16124 26850 16136
rect 27632 16108 27660 16136
rect 20257 16059 20315 16065
rect 20364 16068 22232 16096
rect 23569 16099 23627 16105
rect 12452 15960 12480 16059
rect 19628 16028 19656 16059
rect 20070 16028 20076 16040
rect 19628 16000 20076 16028
rect 20070 15988 20076 16000
rect 20128 16028 20134 16040
rect 20364 16028 20392 16068
rect 23569 16065 23581 16099
rect 23615 16065 23627 16099
rect 23569 16059 23627 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26142 16096 26148 16108
rect 26099 16068 26148 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 26326 16056 26332 16108
rect 26384 16096 26390 16108
rect 26602 16096 26608 16108
rect 26384 16068 26608 16096
rect 26384 16056 26390 16068
rect 26602 16056 26608 16068
rect 26660 16096 26666 16108
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 26660 16068 27353 16096
rect 26660 16056 26666 16068
rect 27341 16065 27353 16068
rect 27387 16096 27399 16099
rect 27387 16068 27568 16096
rect 27387 16065 27399 16068
rect 27341 16059 27399 16065
rect 20128 16000 20392 16028
rect 20441 16031 20499 16037
rect 20128 15988 20134 16000
rect 20441 15997 20453 16031
rect 20487 16028 20499 16031
rect 20530 16028 20536 16040
rect 20487 16000 20536 16028
rect 20487 15997 20499 16000
rect 20441 15991 20499 15997
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 16028 22523 16031
rect 23842 16028 23848 16040
rect 22511 16000 23848 16028
rect 22511 15997 22523 16000
rect 22465 15991 22523 15997
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 24394 16028 24400 16040
rect 24355 16000 24400 16028
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 26237 16031 26295 16037
rect 26237 15997 26249 16031
rect 26283 16028 26295 16031
rect 27540 16028 27568 16068
rect 27614 16056 27620 16108
rect 27672 16096 27678 16108
rect 27801 16099 27859 16105
rect 27801 16096 27813 16099
rect 27672 16068 27813 16096
rect 27672 16056 27678 16068
rect 27801 16065 27813 16068
rect 27847 16065 27859 16099
rect 27801 16059 27859 16065
rect 28445 16031 28503 16037
rect 28445 16028 28457 16031
rect 26283 16000 27476 16028
rect 27540 16000 28457 16028
rect 26283 15997 26295 16000
rect 26237 15991 26295 15997
rect 22002 15960 22008 15972
rect 12452 15932 22008 15960
rect 22002 15920 22008 15932
rect 22060 15920 22066 15972
rect 23017 15963 23075 15969
rect 23017 15929 23029 15963
rect 23063 15960 23075 15963
rect 23290 15960 23296 15972
rect 23063 15932 23296 15960
rect 23063 15929 23075 15932
rect 23017 15923 23075 15929
rect 23290 15920 23296 15932
rect 23348 15920 23354 15972
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 23532 15932 24440 15960
rect 23532 15920 23538 15932
rect 19705 15895 19763 15901
rect 19705 15861 19717 15895
rect 19751 15892 19763 15895
rect 20806 15892 20812 15904
rect 19751 15864 20812 15892
rect 19751 15861 19763 15864
rect 19705 15855 19763 15861
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 20901 15895 20959 15901
rect 20901 15861 20913 15895
rect 20947 15892 20959 15895
rect 21082 15892 21088 15904
rect 20947 15864 21088 15892
rect 20947 15861 20959 15864
rect 20901 15855 20959 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 23658 15892 23664 15904
rect 23619 15864 23664 15892
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 24412 15892 24440 15932
rect 27448 15904 27476 16000
rect 28445 15997 28457 16000
rect 28491 15997 28503 16031
rect 28445 15991 28503 15997
rect 25593 15895 25651 15901
rect 25593 15892 25605 15895
rect 24412 15864 25605 15892
rect 25593 15861 25605 15864
rect 25639 15892 25651 15895
rect 26510 15892 26516 15904
rect 25639 15864 26516 15892
rect 25639 15861 25651 15864
rect 25593 15855 25651 15861
rect 26510 15852 26516 15864
rect 26568 15852 26574 15904
rect 27246 15892 27252 15904
rect 27207 15864 27252 15892
rect 27246 15852 27252 15864
rect 27304 15852 27310 15904
rect 27430 15852 27436 15904
rect 27488 15892 27494 15904
rect 27893 15895 27951 15901
rect 27893 15892 27905 15895
rect 27488 15864 27905 15892
rect 27488 15852 27494 15864
rect 27893 15861 27905 15864
rect 27939 15861 27951 15895
rect 36354 15892 36360 15904
rect 36315 15864 36360 15892
rect 27893 15855 27951 15861
rect 36354 15852 36360 15864
rect 36412 15852 36418 15904
rect 1104 15802 36892 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36892 15802
rect 1104 15728 36892 15750
rect 18877 15691 18935 15697
rect 18877 15657 18889 15691
rect 18923 15688 18935 15691
rect 19334 15688 19340 15700
rect 18923 15660 19340 15688
rect 18923 15657 18935 15660
rect 18877 15651 18935 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 27982 15688 27988 15700
rect 21692 15660 27988 15688
rect 21692 15648 21698 15660
rect 27982 15648 27988 15660
rect 28040 15688 28046 15700
rect 28997 15691 29055 15697
rect 28997 15688 29009 15691
rect 28040 15660 29009 15688
rect 28040 15648 28046 15660
rect 28997 15657 29009 15660
rect 29043 15657 29055 15691
rect 33594 15688 33600 15700
rect 33555 15660 33600 15688
rect 28997 15651 29055 15657
rect 33594 15648 33600 15660
rect 33652 15648 33658 15700
rect 28074 15580 28080 15632
rect 28132 15620 28138 15632
rect 28132 15592 31754 15620
rect 28132 15580 28138 15592
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 20809 15555 20867 15561
rect 20809 15552 20821 15555
rect 19392 15524 20821 15552
rect 19392 15512 19398 15524
rect 20809 15521 20821 15524
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22557 15555 22615 15561
rect 22557 15552 22569 15555
rect 22152 15524 22569 15552
rect 22152 15512 22158 15524
rect 22557 15521 22569 15524
rect 22603 15552 22615 15555
rect 23201 15555 23259 15561
rect 23201 15552 23213 15555
rect 22603 15524 23213 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 23201 15521 23213 15524
rect 23247 15521 23259 15555
rect 23201 15515 23259 15521
rect 23290 15512 23296 15564
rect 23348 15552 23354 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 23348 15524 25145 15552
rect 23348 15512 23354 15524
rect 25133 15521 25145 15524
rect 25179 15552 25191 15555
rect 25222 15552 25228 15564
rect 25179 15524 25228 15552
rect 25179 15521 25191 15524
rect 25133 15515 25191 15521
rect 25222 15512 25228 15524
rect 25280 15512 25286 15564
rect 27706 15512 27712 15564
rect 27764 15552 27770 15564
rect 31726 15552 31754 15592
rect 36081 15555 36139 15561
rect 36081 15552 36093 15555
rect 27764 15524 27809 15552
rect 31726 15524 36093 15552
rect 27764 15512 27770 15524
rect 36081 15521 36093 15524
rect 36127 15521 36139 15555
rect 36081 15515 36139 15521
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15484 18383 15487
rect 19058 15484 19064 15496
rect 18371 15456 19064 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 27154 15444 27160 15496
rect 27212 15484 27218 15496
rect 27212 15456 27257 15484
rect 27212 15444 27218 15456
rect 27606 15444 27612 15496
rect 27664 15484 27670 15496
rect 31665 15487 31723 15493
rect 27664 15456 27709 15484
rect 27664 15444 27670 15456
rect 31665 15453 31677 15487
rect 31711 15484 31723 15487
rect 33410 15484 33416 15496
rect 31711 15456 32260 15484
rect 33371 15456 33416 15484
rect 31711 15453 31723 15456
rect 31665 15447 31723 15453
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 6886 15388 19993 15416
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 6886 15348 6914 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 20165 15419 20223 15425
rect 20165 15385 20177 15419
rect 20211 15385 20223 15419
rect 20165 15379 20223 15385
rect 4764 15320 6914 15348
rect 19521 15351 19579 15357
rect 4764 15308 4770 15320
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 20180 15348 20208 15379
rect 20898 15376 20904 15428
rect 20956 15416 20962 15428
rect 21453 15419 21511 15425
rect 20956 15388 21001 15416
rect 20956 15376 20962 15388
rect 21453 15385 21465 15419
rect 21499 15416 21511 15419
rect 21726 15416 21732 15428
rect 21499 15388 21732 15416
rect 21499 15385 21511 15388
rect 21453 15379 21511 15385
rect 21726 15376 21732 15388
rect 21784 15416 21790 15428
rect 21913 15419 21971 15425
rect 21913 15416 21925 15419
rect 21784 15388 21925 15416
rect 21784 15376 21790 15388
rect 21913 15385 21925 15388
rect 21959 15385 21971 15419
rect 22462 15416 22468 15428
rect 22423 15388 22468 15416
rect 21913 15379 21971 15385
rect 22462 15376 22468 15388
rect 22520 15376 22526 15428
rect 23293 15419 23351 15425
rect 23293 15385 23305 15419
rect 23339 15416 23351 15419
rect 23566 15416 23572 15428
rect 23339 15388 23572 15416
rect 23339 15385 23351 15388
rect 23293 15379 23351 15385
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 23845 15419 23903 15425
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 24302 15416 24308 15428
rect 23891 15388 24308 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 24302 15376 24308 15388
rect 24360 15376 24366 15428
rect 25317 15419 25375 15425
rect 25317 15385 25329 15419
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 25409 15419 25467 15425
rect 25409 15385 25421 15419
rect 25455 15416 25467 15419
rect 26326 15416 26332 15428
rect 25455 15388 26332 15416
rect 25455 15385 25467 15388
rect 25409 15379 25467 15385
rect 22186 15348 22192 15360
rect 19567 15320 22192 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 25332 15348 25360 15379
rect 26326 15376 26332 15388
rect 26384 15376 26390 15428
rect 26510 15416 26516 15428
rect 26471 15388 26516 15416
rect 26510 15376 26516 15388
rect 26568 15376 26574 15428
rect 26605 15419 26663 15425
rect 26605 15385 26617 15419
rect 26651 15416 26663 15419
rect 26970 15416 26976 15428
rect 26651 15388 26976 15416
rect 26651 15385 26663 15388
rect 26605 15379 26663 15385
rect 26970 15376 26976 15388
rect 27028 15376 27034 15428
rect 27890 15376 27896 15428
rect 27948 15416 27954 15428
rect 31573 15419 31631 15425
rect 31573 15416 31585 15419
rect 27948 15388 31585 15416
rect 27948 15376 27954 15388
rect 31573 15385 31585 15388
rect 31619 15385 31631 15419
rect 31573 15379 31631 15385
rect 27522 15348 27528 15360
rect 25332 15320 27528 15348
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 28258 15348 28264 15360
rect 28219 15320 28264 15348
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 32232 15357 32260 15456
rect 33410 15444 33416 15456
rect 33468 15444 33474 15496
rect 36354 15484 36360 15496
rect 36315 15456 36360 15484
rect 36354 15444 36360 15456
rect 36412 15444 36418 15496
rect 32217 15351 32275 15357
rect 32217 15317 32229 15351
rect 32263 15348 32275 15351
rect 35526 15348 35532 15360
rect 32263 15320 35532 15348
rect 32263 15317 32275 15320
rect 32217 15311 32275 15317
rect 35526 15308 35532 15320
rect 35584 15308 35590 15360
rect 1104 15258 36892 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 36892 15258
rect 1104 15184 36892 15206
rect 19061 15147 19119 15153
rect 19061 15113 19073 15147
rect 19107 15144 19119 15147
rect 20530 15144 20536 15156
rect 19107 15116 20536 15144
rect 19107 15113 19119 15116
rect 19061 15107 19119 15113
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 24946 15144 24952 15156
rect 22888 15116 24952 15144
rect 22888 15104 22894 15116
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 26326 15104 26332 15156
rect 26384 15144 26390 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 26384 15116 27169 15144
rect 26384 15104 26390 15116
rect 27157 15113 27169 15116
rect 27203 15113 27215 15147
rect 27157 15107 27215 15113
rect 27522 15104 27528 15156
rect 27580 15144 27586 15156
rect 29181 15147 29239 15153
rect 29181 15144 29193 15147
rect 27580 15116 29193 15144
rect 27580 15104 27586 15116
rect 29181 15113 29193 15116
rect 29227 15113 29239 15147
rect 36078 15144 36084 15156
rect 36039 15116 36084 15144
rect 29181 15107 29239 15113
rect 36078 15104 36084 15116
rect 36136 15104 36142 15156
rect 20257 15079 20315 15085
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 21082 15076 21088 15088
rect 20303 15048 21088 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 21082 15036 21088 15048
rect 21140 15076 21146 15088
rect 21361 15079 21419 15085
rect 21361 15076 21373 15079
rect 21140 15048 21373 15076
rect 21140 15036 21146 15048
rect 21361 15045 21373 15048
rect 21407 15045 21419 15079
rect 21361 15039 21419 15045
rect 22281 15079 22339 15085
rect 22281 15045 22293 15079
rect 22327 15076 22339 15079
rect 23658 15076 23664 15088
rect 22327 15048 23664 15076
rect 22327 15045 22339 15048
rect 22281 15039 22339 15045
rect 23658 15036 23664 15048
rect 23716 15036 23722 15088
rect 25225 15079 25283 15085
rect 25225 15045 25237 15079
rect 25271 15076 25283 15079
rect 27893 15079 27951 15085
rect 27893 15076 27905 15079
rect 25271 15048 27905 15076
rect 25271 15045 25283 15048
rect 25225 15039 25283 15045
rect 27893 15045 27905 15048
rect 27939 15045 27951 15079
rect 27893 15039 27951 15045
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17862 15008 17868 15020
rect 17267 14980 17868 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 18969 15011 19027 15017
rect 18969 14977 18981 15011
rect 19015 15008 19027 15011
rect 19058 15008 19064 15020
rect 19015 14980 19064 15008
rect 19015 14977 19027 14980
rect 18969 14971 19027 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19392 14980 19625 15008
rect 19392 14968 19398 14980
rect 19613 14977 19625 14980
rect 19659 14977 19671 15011
rect 19613 14971 19671 14977
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 20162 15008 20168 15020
rect 19843 14980 20168 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20714 15008 20720 15020
rect 20675 14980 20720 15008
rect 20714 14968 20720 14980
rect 20772 14968 20778 15020
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 20990 15008 20996 15020
rect 20947 14980 20996 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 23014 14968 23020 15020
rect 23072 15008 23078 15020
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 23072 14980 23489 15008
rect 23072 14968 23078 14980
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 25866 15008 25872 15020
rect 25827 14980 25872 15008
rect 23477 14971 23535 14977
rect 25866 14968 25872 14980
rect 25924 14968 25930 15020
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 15008 26111 15011
rect 27246 15008 27252 15020
rect 26099 14980 27252 15008
rect 26099 14977 26111 14980
rect 26053 14971 26111 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 27982 15008 27988 15020
rect 27943 14980 27988 15008
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 28629 15011 28687 15017
rect 28629 14977 28641 15011
rect 28675 14977 28687 15011
rect 28629 14971 28687 14977
rect 18506 14940 18512 14952
rect 18467 14912 18512 14940
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 19978 14900 19984 14952
rect 20036 14940 20042 14952
rect 22189 14943 22247 14949
rect 22189 14940 22201 14943
rect 20036 14912 22201 14940
rect 20036 14900 20042 14912
rect 22189 14909 22201 14912
rect 22235 14940 22247 14943
rect 22830 14940 22836 14952
rect 22235 14912 22836 14940
rect 22235 14909 22247 14912
rect 22189 14903 22247 14909
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 23661 14943 23719 14949
rect 23661 14909 23673 14943
rect 23707 14940 23719 14943
rect 24854 14940 24860 14952
rect 23707 14912 24860 14940
rect 23707 14909 23719 14912
rect 23661 14903 23719 14909
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 25314 14940 25320 14952
rect 25275 14912 25320 14940
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 27338 14900 27344 14952
rect 27396 14940 27402 14952
rect 28537 14943 28595 14949
rect 28537 14940 28549 14943
rect 27396 14912 28549 14940
rect 27396 14900 27402 14912
rect 28537 14909 28549 14912
rect 28583 14909 28595 14943
rect 28644 14940 28672 14971
rect 28718 14968 28724 15020
rect 28776 15008 28782 15020
rect 29273 15011 29331 15017
rect 29273 15008 29285 15011
rect 28776 14980 29285 15008
rect 28776 14968 28782 14980
rect 29273 14977 29285 14980
rect 29319 14977 29331 15011
rect 29273 14971 29331 14977
rect 35897 15011 35955 15017
rect 35897 14977 35909 15011
rect 35943 15008 35955 15011
rect 35986 15008 35992 15020
rect 35943 14980 35992 15008
rect 35943 14977 35955 14980
rect 35897 14971 35955 14977
rect 35986 14968 35992 14980
rect 36044 14968 36050 15020
rect 29086 14940 29092 14952
rect 28644 14912 29092 14940
rect 28537 14903 28595 14909
rect 29086 14900 29092 14912
rect 29144 14940 29150 14952
rect 29733 14943 29791 14949
rect 29733 14940 29745 14943
rect 29144 14912 29745 14940
rect 29144 14900 29150 14912
rect 29733 14909 29745 14912
rect 29779 14909 29791 14943
rect 29733 14903 29791 14909
rect 22741 14875 22799 14881
rect 22741 14841 22753 14875
rect 22787 14841 22799 14875
rect 22741 14835 22799 14841
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 17460 14776 17693 14804
rect 17460 14764 17466 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 22756 14804 22784 14835
rect 23474 14832 23480 14884
rect 23532 14872 23538 14884
rect 23845 14875 23903 14881
rect 23845 14872 23857 14875
rect 23532 14844 23857 14872
rect 23532 14832 23538 14844
rect 23845 14841 23857 14844
rect 23891 14841 23903 14875
rect 23845 14835 23903 14841
rect 24765 14875 24823 14881
rect 24765 14841 24777 14875
rect 24811 14872 24823 14875
rect 25130 14872 25136 14884
rect 24811 14844 25136 14872
rect 24811 14841 24823 14844
rect 24765 14835 24823 14841
rect 25130 14832 25136 14844
rect 25188 14872 25194 14884
rect 26050 14872 26056 14884
rect 25188 14844 26056 14872
rect 25188 14832 25194 14844
rect 26050 14832 26056 14844
rect 26108 14832 26114 14884
rect 26142 14832 26148 14884
rect 26200 14872 26206 14884
rect 26878 14872 26884 14884
rect 26200 14844 26884 14872
rect 26200 14832 26206 14844
rect 26878 14832 26884 14844
rect 26936 14872 26942 14884
rect 30834 14872 30840 14884
rect 26936 14844 30840 14872
rect 26936 14832 26942 14844
rect 30834 14832 30840 14844
rect 30892 14832 30898 14884
rect 24394 14804 24400 14816
rect 22756 14776 24400 14804
rect 17681 14767 17739 14773
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 26234 14804 26240 14816
rect 26195 14776 26240 14804
rect 26234 14764 26240 14776
rect 26292 14764 26298 14816
rect 1104 14714 36892 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36892 14714
rect 1104 14640 36892 14662
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 17920 14572 18153 14600
rect 17920 14560 17926 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 18141 14563 18199 14569
rect 22281 14603 22339 14609
rect 22281 14569 22293 14603
rect 22327 14600 22339 14603
rect 22554 14600 22560 14612
rect 22327 14572 22560 14600
rect 22327 14569 22339 14572
rect 22281 14563 22339 14569
rect 1854 14396 1860 14408
rect 1815 14368 1860 14396
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 18156 14396 18184 14563
rect 22554 14560 22560 14572
rect 22612 14560 22618 14612
rect 22830 14600 22836 14612
rect 22791 14572 22836 14600
rect 22830 14560 22836 14572
rect 22888 14560 22894 14612
rect 23566 14560 23572 14612
rect 23624 14600 23630 14612
rect 24673 14603 24731 14609
rect 24673 14600 24685 14603
rect 23624 14572 24685 14600
rect 23624 14560 23630 14572
rect 24673 14569 24685 14572
rect 24719 14569 24731 14603
rect 24673 14563 24731 14569
rect 26602 14560 26608 14612
rect 26660 14600 26666 14612
rect 27890 14600 27896 14612
rect 26660 14572 27896 14600
rect 26660 14560 26666 14572
rect 27890 14560 27896 14572
rect 27948 14560 27954 14612
rect 27706 14532 27712 14544
rect 23584 14504 27712 14532
rect 18506 14424 18512 14476
rect 18564 14464 18570 14476
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 18564 14436 20085 14464
rect 18564 14424 18570 14436
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20806 14464 20812 14476
rect 20767 14436 20812 14464
rect 20073 14427 20131 14433
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 21082 14424 21088 14476
rect 21140 14464 21146 14476
rect 23584 14473 23612 14504
rect 27706 14492 27712 14504
rect 27764 14492 27770 14544
rect 27982 14492 27988 14544
rect 28040 14532 28046 14544
rect 30006 14532 30012 14544
rect 28040 14504 30012 14532
rect 28040 14492 28046 14504
rect 30006 14492 30012 14504
rect 30064 14492 30070 14544
rect 21637 14467 21695 14473
rect 21637 14464 21649 14467
rect 21140 14436 21649 14464
rect 21140 14424 21146 14436
rect 21637 14433 21649 14436
rect 21683 14433 21695 14467
rect 21637 14427 21695 14433
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14433 23627 14467
rect 23569 14427 23627 14433
rect 25961 14467 26019 14473
rect 25961 14433 25973 14467
rect 26007 14464 26019 14467
rect 29089 14467 29147 14473
rect 29089 14464 29101 14467
rect 26007 14436 29101 14464
rect 26007 14433 26019 14436
rect 25961 14427 26019 14433
rect 29089 14433 29101 14436
rect 29135 14433 29147 14467
rect 29089 14427 29147 14433
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 18156 14368 18705 14396
rect 18693 14365 18705 14368
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20714 14396 20720 14408
rect 19935 14368 20720 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 21818 14356 21824 14408
rect 21876 14396 21882 14408
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 21876 14368 22201 14396
rect 21876 14356 21882 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 23382 14396 23388 14408
rect 23343 14368 23388 14396
rect 22189 14359 22247 14365
rect 2038 14288 2044 14340
rect 2096 14328 2102 14340
rect 20806 14328 20812 14340
rect 2096 14300 20812 14328
rect 2096 14288 2102 14300
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 21545 14331 21603 14337
rect 21545 14297 21557 14331
rect 21591 14297 21603 14331
rect 22204 14328 22232 14359
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 24762 14396 24768 14408
rect 23492 14368 24768 14396
rect 23492 14328 23520 14368
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 26142 14396 26148 14408
rect 26103 14368 26148 14396
rect 26142 14356 26148 14368
rect 26200 14356 26206 14408
rect 28534 14356 28540 14408
rect 28592 14396 28598 14408
rect 28592 14368 28637 14396
rect 28592 14356 28598 14368
rect 28994 14356 29000 14408
rect 29052 14396 29058 14408
rect 29546 14396 29552 14408
rect 29052 14368 29552 14396
rect 29052 14356 29058 14368
rect 29546 14356 29552 14368
rect 29604 14356 29610 14408
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14396 29975 14399
rect 29963 14368 30512 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 22204 14300 23520 14328
rect 21545 14291 21603 14297
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 18785 14263 18843 14269
rect 18785 14229 18797 14263
rect 18831 14260 18843 14263
rect 19334 14260 19340 14272
rect 18831 14232 19340 14260
rect 18831 14229 18843 14232
rect 18785 14223 18843 14229
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 21560 14260 21588 14291
rect 24394 14288 24400 14340
rect 24452 14328 24458 14340
rect 26602 14328 26608 14340
rect 24452 14300 26608 14328
rect 24452 14288 24458 14300
rect 26602 14288 26608 14300
rect 26660 14288 26666 14340
rect 27157 14331 27215 14337
rect 27157 14297 27169 14331
rect 27203 14297 27215 14331
rect 27157 14291 27215 14297
rect 27249 14331 27307 14337
rect 27249 14297 27261 14331
rect 27295 14328 27307 14331
rect 27706 14328 27712 14340
rect 27295 14300 27712 14328
rect 27295 14297 27307 14300
rect 27249 14291 27307 14297
rect 22278 14260 22284 14272
rect 19484 14232 19529 14260
rect 21560 14232 22284 14260
rect 19484 14220 19490 14232
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 24029 14263 24087 14269
rect 24029 14229 24041 14263
rect 24075 14260 24087 14263
rect 25501 14263 25559 14269
rect 25501 14260 25513 14263
rect 24075 14232 25513 14260
rect 24075 14229 24087 14232
rect 24029 14223 24087 14229
rect 25501 14229 25513 14232
rect 25547 14260 25559 14263
rect 26234 14260 26240 14272
rect 25547 14232 26240 14260
rect 25547 14229 25559 14232
rect 25501 14223 25559 14229
rect 26234 14220 26240 14232
rect 26292 14220 26298 14272
rect 27172 14260 27200 14291
rect 27706 14288 27712 14300
rect 27764 14288 27770 14340
rect 27890 14328 27896 14340
rect 27851 14300 27896 14328
rect 27890 14288 27896 14300
rect 27948 14288 27954 14340
rect 27982 14288 27988 14340
rect 28040 14328 28046 14340
rect 28040 14300 28085 14328
rect 28040 14288 28046 14300
rect 28626 14288 28632 14340
rect 28684 14328 28690 14340
rect 29825 14331 29883 14337
rect 29825 14328 29837 14331
rect 28684 14300 29837 14328
rect 28684 14288 28690 14300
rect 29825 14297 29837 14300
rect 29871 14297 29883 14331
rect 29825 14291 29883 14297
rect 29730 14260 29736 14272
rect 27172 14232 29736 14260
rect 29730 14220 29736 14232
rect 29788 14220 29794 14272
rect 30484 14269 30512 14368
rect 30469 14263 30527 14269
rect 30469 14229 30481 14263
rect 30515 14260 30527 14263
rect 34606 14260 34612 14272
rect 30515 14232 34612 14260
rect 30515 14229 30527 14232
rect 30469 14223 30527 14229
rect 34606 14220 34612 14232
rect 34664 14220 34670 14272
rect 1104 14170 36892 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 36892 14170
rect 1104 14096 36892 14118
rect 17034 14056 17040 14068
rect 16995 14028 17040 14056
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 17954 14056 17960 14068
rect 17727 14028 17960 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 22738 14056 22744 14068
rect 22152 14028 22197 14056
rect 22699 14028 22744 14056
rect 22152 14016 22158 14028
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 23382 14016 23388 14068
rect 23440 14056 23446 14068
rect 24489 14059 24547 14065
rect 24489 14056 24501 14059
rect 23440 14028 24501 14056
rect 23440 14016 23446 14028
rect 24489 14025 24501 14028
rect 24535 14025 24547 14059
rect 27798 14056 27804 14068
rect 24489 14019 24547 14025
rect 25700 14028 27804 14056
rect 17052 13920 17080 14016
rect 19334 13948 19340 14000
rect 19392 13988 19398 14000
rect 20073 13991 20131 13997
rect 20073 13988 20085 13991
rect 19392 13960 20085 13988
rect 19392 13948 19398 13960
rect 20073 13957 20085 13960
rect 20119 13957 20131 13991
rect 20073 13951 20131 13957
rect 20165 13991 20223 13997
rect 20165 13957 20177 13991
rect 20211 13988 20223 13991
rect 21269 13991 21327 13997
rect 21269 13988 21281 13991
rect 20211 13960 21281 13988
rect 20211 13957 20223 13960
rect 20165 13951 20223 13957
rect 21269 13957 21281 13960
rect 21315 13957 21327 13991
rect 21269 13951 21327 13957
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17052 13892 18153 13920
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 21818 13920 21824 13932
rect 21407 13892 21824 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22002 13880 22008 13932
rect 22060 13920 22066 13932
rect 22756 13920 22784 14016
rect 23750 13988 23756 14000
rect 23711 13960 23756 13988
rect 23750 13948 23756 13960
rect 23808 13948 23814 14000
rect 25700 13997 25728 14028
rect 27798 14016 27804 14028
rect 27856 14016 27862 14068
rect 28810 14056 28816 14068
rect 28771 14028 28816 14056
rect 28810 14016 28816 14028
rect 28868 14016 28874 14068
rect 28994 14016 29000 14068
rect 29052 14016 29058 14068
rect 29730 14016 29736 14068
rect 29788 14056 29794 14068
rect 30193 14059 30251 14065
rect 30193 14056 30205 14059
rect 29788 14028 30205 14056
rect 29788 14016 29794 14028
rect 30193 14025 30205 14028
rect 30239 14025 30251 14059
rect 30834 14056 30840 14068
rect 30795 14028 30840 14056
rect 30193 14019 30251 14025
rect 30834 14016 30840 14028
rect 30892 14016 30898 14068
rect 25685 13991 25743 13997
rect 25685 13957 25697 13991
rect 25731 13957 25743 13991
rect 25685 13951 25743 13957
rect 25774 13948 25780 14000
rect 25832 13988 25838 14000
rect 25832 13960 25877 13988
rect 25832 13948 25838 13960
rect 26234 13948 26240 14000
rect 26292 13988 26298 14000
rect 27617 13991 27675 13997
rect 27617 13988 27629 13991
rect 26292 13960 27629 13988
rect 26292 13948 26298 13960
rect 27617 13957 27629 13960
rect 27663 13957 27675 13991
rect 27617 13951 27675 13957
rect 27709 13991 27767 13997
rect 27709 13957 27721 13991
rect 27755 13988 27767 13991
rect 29012 13988 29040 14016
rect 27755 13960 29040 13988
rect 27755 13957 27767 13960
rect 27709 13951 27767 13957
rect 22060 13892 22784 13920
rect 24581 13923 24639 13929
rect 22060 13880 22066 13892
rect 24581 13889 24593 13923
rect 24627 13920 24639 13923
rect 24854 13920 24860 13932
rect 24627 13892 24860 13920
rect 24627 13889 24639 13892
rect 24581 13883 24639 13889
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 25958 13880 25964 13932
rect 26016 13920 26022 13932
rect 26513 13923 26571 13929
rect 26513 13920 26525 13923
rect 26016 13892 26525 13920
rect 26016 13880 26022 13892
rect 26513 13889 26525 13892
rect 26559 13920 26571 13923
rect 28905 13923 28963 13929
rect 26559 13892 27476 13920
rect 26559 13889 26571 13892
rect 26513 13883 26571 13889
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18782 13852 18788 13864
rect 18012 13824 18788 13852
rect 18012 13812 18018 13824
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 18966 13852 18972 13864
rect 18927 13824 18972 13852
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 22922 13852 22928 13864
rect 20763 13824 22928 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 22922 13812 22928 13824
rect 22980 13812 22986 13864
rect 23385 13855 23443 13861
rect 23385 13821 23397 13855
rect 23431 13821 23443 13855
rect 23385 13815 23443 13821
rect 21174 13744 21180 13796
rect 21232 13784 21238 13796
rect 23400 13784 23428 13815
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 23845 13855 23903 13861
rect 23845 13852 23857 13855
rect 23532 13824 23857 13852
rect 23532 13812 23538 13824
rect 23845 13821 23857 13824
rect 23891 13852 23903 13855
rect 23891 13824 25452 13852
rect 23891 13821 23903 13824
rect 23845 13815 23903 13821
rect 23658 13784 23664 13796
rect 21232 13756 23336 13784
rect 23400 13756 23664 13784
rect 21232 13744 21238 13756
rect 18230 13716 18236 13728
rect 18191 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 22370 13716 22376 13728
rect 18380 13688 22376 13716
rect 18380 13676 18386 13688
rect 22370 13676 22376 13688
rect 22428 13676 22434 13728
rect 23308 13716 23336 13756
rect 23658 13744 23664 13756
rect 23716 13744 23722 13796
rect 25424 13784 25452 13824
rect 25498 13812 25504 13864
rect 25556 13852 25562 13864
rect 26602 13852 26608 13864
rect 25556 13824 26608 13852
rect 25556 13812 25562 13824
rect 26602 13812 26608 13824
rect 26660 13812 26666 13864
rect 26421 13787 26479 13793
rect 26421 13784 26433 13787
rect 25424 13756 26433 13784
rect 26421 13753 26433 13756
rect 26467 13753 26479 13787
rect 27448 13784 27476 13892
rect 28905 13889 28917 13923
rect 28951 13920 28963 13923
rect 29362 13920 29368 13932
rect 28951 13892 29368 13920
rect 28951 13889 28963 13892
rect 28905 13883 28963 13889
rect 29362 13880 29368 13892
rect 29420 13880 29426 13932
rect 29641 13923 29699 13929
rect 29641 13889 29653 13923
rect 29687 13889 29699 13923
rect 29641 13883 29699 13889
rect 30101 13923 30159 13929
rect 30101 13889 30113 13923
rect 30147 13889 30159 13923
rect 30101 13883 30159 13889
rect 30929 13923 30987 13929
rect 30929 13889 30941 13923
rect 30975 13920 30987 13923
rect 33410 13920 33416 13932
rect 30975 13892 33416 13920
rect 30975 13889 30987 13892
rect 30929 13883 30987 13889
rect 27706 13812 27712 13864
rect 27764 13852 27770 13864
rect 29549 13855 29607 13861
rect 29549 13852 29561 13855
rect 27764 13824 29561 13852
rect 27764 13812 27770 13824
rect 29549 13821 29561 13824
rect 29595 13821 29607 13855
rect 29549 13815 29607 13821
rect 27522 13784 27528 13796
rect 27448 13756 27528 13784
rect 26421 13747 26479 13753
rect 27522 13744 27528 13756
rect 27580 13744 27586 13796
rect 28166 13784 28172 13796
rect 28127 13756 28172 13784
rect 28166 13744 28172 13756
rect 28224 13744 28230 13796
rect 28810 13744 28816 13796
rect 28868 13784 28874 13796
rect 29656 13784 29684 13883
rect 30116 13852 30144 13883
rect 33410 13880 33416 13892
rect 33468 13880 33474 13932
rect 28868 13756 29684 13784
rect 29748 13824 30144 13852
rect 28868 13744 28874 13756
rect 28442 13716 28448 13728
rect 23308 13688 28448 13716
rect 28442 13676 28448 13688
rect 28500 13676 28506 13728
rect 28902 13676 28908 13728
rect 28960 13716 28966 13728
rect 29748 13716 29776 13824
rect 28960 13688 29776 13716
rect 28960 13676 28966 13688
rect 1104 13626 36892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36892 13626
rect 1104 13552 36892 13574
rect 17589 13515 17647 13521
rect 17589 13481 17601 13515
rect 17635 13512 17647 13515
rect 17954 13512 17960 13524
rect 17635 13484 17960 13512
rect 17635 13481 17647 13484
rect 17589 13475 17647 13481
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 18785 13515 18843 13521
rect 18785 13481 18797 13515
rect 18831 13512 18843 13515
rect 18966 13512 18972 13524
rect 18831 13484 18972 13512
rect 18831 13481 18843 13484
rect 18785 13475 18843 13481
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 22186 13512 22192 13524
rect 19260 13484 22192 13512
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 19260 13376 19288 13484
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22281 13515 22339 13521
rect 22281 13481 22293 13515
rect 22327 13512 22339 13515
rect 22462 13512 22468 13524
rect 22327 13484 22468 13512
rect 22327 13481 22339 13484
rect 22281 13475 22339 13481
rect 22462 13472 22468 13484
rect 22520 13472 22526 13524
rect 25038 13472 25044 13524
rect 25096 13512 25102 13524
rect 25958 13512 25964 13524
rect 25096 13484 25964 13512
rect 25096 13472 25102 13484
rect 25958 13472 25964 13484
rect 26016 13472 26022 13524
rect 26050 13472 26056 13524
rect 26108 13512 26114 13524
rect 28626 13512 28632 13524
rect 26108 13484 28632 13512
rect 26108 13472 26114 13484
rect 28626 13472 28632 13484
rect 28684 13472 28690 13524
rect 21637 13447 21695 13453
rect 21637 13413 21649 13447
rect 21683 13444 21695 13447
rect 23658 13444 23664 13456
rect 21683 13416 23664 13444
rect 21683 13413 21695 13416
rect 21637 13407 21695 13413
rect 23658 13404 23664 13416
rect 23716 13404 23722 13456
rect 29089 13447 29147 13453
rect 29089 13444 29101 13447
rect 24228 13416 29101 13444
rect 17083 13348 19288 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19521 13379 19579 13385
rect 19521 13376 19533 13379
rect 19392 13348 19533 13376
rect 19392 13336 19398 13348
rect 19521 13345 19533 13348
rect 19567 13345 19579 13379
rect 19521 13339 19579 13345
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13376 21143 13379
rect 23382 13376 23388 13388
rect 21131 13348 23388 13376
rect 21131 13345 21143 13348
rect 21085 13339 21143 13345
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13308 18107 13311
rect 18322 13308 18328 13320
rect 18095 13280 18328 13308
rect 18095 13277 18107 13280
rect 18049 13271 18107 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 22186 13308 22192 13320
rect 18923 13280 19288 13308
rect 22147 13280 22192 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 19150 13172 19156 13184
rect 18187 13144 19156 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 19260 13172 19288 13280
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 19392 13212 19625 13240
rect 19392 13200 19398 13212
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 20162 13240 20168 13252
rect 20123 13212 20168 13240
rect 19613 13203 19671 13209
rect 20162 13200 20168 13212
rect 20220 13200 20226 13252
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 21177 13243 21235 13249
rect 21177 13240 21189 13243
rect 20680 13212 21189 13240
rect 20680 13200 20686 13212
rect 21177 13209 21189 13212
rect 21223 13209 21235 13243
rect 22922 13240 22928 13252
rect 22883 13212 22928 13240
rect 21177 13203 21235 13209
rect 22922 13200 22928 13212
rect 22980 13200 22986 13252
rect 23477 13243 23535 13249
rect 23477 13209 23489 13243
rect 23523 13209 23535 13243
rect 23477 13203 23535 13209
rect 20438 13172 20444 13184
rect 19260 13144 20444 13172
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 23492 13172 23520 13203
rect 23566 13200 23572 13252
rect 23624 13240 23630 13252
rect 23624 13212 23669 13240
rect 23624 13200 23630 13212
rect 24228 13172 24256 13416
rect 29089 13413 29101 13416
rect 29135 13413 29147 13447
rect 29089 13407 29147 13413
rect 29917 13447 29975 13453
rect 29917 13413 29929 13447
rect 29963 13444 29975 13447
rect 29963 13416 35894 13444
rect 29963 13413 29975 13416
rect 29917 13407 29975 13413
rect 25774 13336 25780 13388
rect 25832 13376 25838 13388
rect 26050 13376 26056 13388
rect 25832 13348 26056 13376
rect 25832 13336 25838 13348
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 26602 13376 26608 13388
rect 26563 13348 26608 13376
rect 26602 13336 26608 13348
rect 26660 13336 26666 13388
rect 28442 13336 28448 13388
rect 28500 13376 28506 13388
rect 30377 13379 30435 13385
rect 30377 13376 30389 13379
rect 28500 13348 30389 13376
rect 28500 13336 28506 13348
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 25038 13308 25044 13320
rect 24811 13280 25044 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 28997 13311 29055 13317
rect 28997 13277 29009 13311
rect 29043 13308 29055 13311
rect 29178 13308 29184 13320
rect 29043 13280 29184 13308
rect 29043 13277 29055 13280
rect 28997 13271 29055 13277
rect 29178 13268 29184 13280
rect 29236 13268 29242 13320
rect 29748 13317 29776 13348
rect 30377 13345 30389 13348
rect 30423 13345 30435 13379
rect 35866 13376 35894 13416
rect 35866 13348 36124 13376
rect 30377 13339 30435 13345
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13277 29791 13311
rect 29733 13271 29791 13277
rect 31757 13311 31815 13317
rect 31757 13277 31769 13311
rect 31803 13308 31815 13311
rect 35986 13308 35992 13320
rect 31803 13280 35992 13308
rect 31803 13277 31815 13280
rect 31757 13271 31815 13277
rect 35986 13268 35992 13280
rect 36044 13268 36050 13320
rect 36096 13317 36124 13348
rect 36081 13311 36139 13317
rect 36081 13277 36093 13311
rect 36127 13277 36139 13311
rect 36081 13271 36139 13277
rect 24302 13200 24308 13252
rect 24360 13240 24366 13252
rect 25314 13240 25320 13252
rect 24360 13212 25320 13240
rect 24360 13200 24366 13212
rect 25314 13200 25320 13212
rect 25372 13240 25378 13252
rect 25409 13243 25467 13249
rect 25409 13240 25421 13243
rect 25372 13212 25421 13240
rect 25372 13200 25378 13212
rect 25409 13209 25421 13212
rect 25455 13209 25467 13243
rect 25958 13240 25964 13252
rect 25919 13212 25964 13240
rect 25409 13203 25467 13209
rect 25958 13200 25964 13212
rect 26016 13200 26022 13252
rect 27157 13243 27215 13249
rect 27157 13209 27169 13243
rect 27203 13209 27215 13243
rect 27157 13203 27215 13209
rect 27249 13243 27307 13249
rect 27249 13209 27261 13243
rect 27295 13240 27307 13243
rect 27430 13240 27436 13252
rect 27295 13212 27436 13240
rect 27295 13209 27307 13212
rect 27249 13203 27307 13209
rect 24578 13172 24584 13184
rect 23492 13144 24256 13172
rect 24539 13144 24584 13172
rect 24578 13132 24584 13144
rect 24636 13132 24642 13184
rect 27172 13172 27200 13203
rect 27430 13200 27436 13212
rect 27488 13200 27494 13252
rect 27522 13200 27528 13252
rect 27580 13240 27586 13252
rect 27801 13243 27859 13249
rect 27801 13240 27813 13243
rect 27580 13212 27813 13240
rect 27580 13200 27586 13212
rect 27801 13209 27813 13212
rect 27847 13209 27859 13243
rect 27801 13203 27859 13209
rect 28166 13200 28172 13252
rect 28224 13240 28230 13252
rect 28353 13243 28411 13249
rect 28353 13240 28365 13243
rect 28224 13212 28365 13240
rect 28224 13200 28230 13212
rect 28353 13209 28365 13212
rect 28399 13209 28411 13243
rect 28353 13203 28411 13209
rect 28445 13243 28503 13249
rect 28445 13209 28457 13243
rect 28491 13240 28503 13243
rect 31665 13243 31723 13249
rect 31665 13240 31677 13243
rect 28491 13212 31677 13240
rect 28491 13209 28503 13212
rect 28445 13203 28503 13209
rect 31665 13209 31677 13212
rect 31711 13209 31723 13243
rect 31665 13203 31723 13209
rect 27982 13172 27988 13184
rect 27172 13144 27988 13172
rect 27982 13132 27988 13144
rect 28040 13132 28046 13184
rect 36262 13172 36268 13184
rect 36223 13144 36268 13172
rect 36262 13132 36268 13144
rect 36320 13132 36326 13184
rect 1104 13082 36892 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 36892 13082
rect 1104 13008 36892 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 2409 12971 2467 12977
rect 2409 12968 2421 12971
rect 1912 12940 2421 12968
rect 1912 12928 1918 12940
rect 2409 12937 2421 12940
rect 2455 12937 2467 12971
rect 2409 12931 2467 12937
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 18509 12971 18567 12977
rect 2740 12940 6914 12968
rect 2740 12928 2746 12940
rect 5626 12900 5632 12912
rect 1872 12872 5632 12900
rect 1872 12841 1900 12872
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 6886 12900 6914 12940
rect 17420 12940 18460 12968
rect 17420 12900 17448 12940
rect 18322 12900 18328 12912
rect 6886 12872 17448 12900
rect 17604 12872 18328 12900
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 17405 12835 17463 12841
rect 2547 12804 3096 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 3068 12705 3096 12804
rect 17405 12801 17417 12835
rect 17451 12832 17463 12835
rect 17604 12832 17632 12872
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 18432 12900 18460 12940
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 19426 12968 19432 12980
rect 18555 12940 19432 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 21177 12971 21235 12977
rect 21177 12968 21189 12971
rect 20772 12940 21189 12968
rect 20772 12928 20778 12940
rect 21177 12937 21189 12940
rect 21223 12937 21235 12971
rect 21177 12931 21235 12937
rect 21818 12928 21824 12980
rect 21876 12968 21882 12980
rect 24578 12968 24584 12980
rect 21876 12940 24584 12968
rect 21876 12928 21882 12940
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 28537 12971 28595 12977
rect 28537 12968 28549 12971
rect 25332 12940 28549 12968
rect 18432 12872 19288 12900
rect 17451 12804 17632 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 17736 12804 18061 12832
rect 17736 12792 17742 12804
rect 18049 12801 18061 12804
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 18782 12792 18788 12844
rect 18840 12832 18846 12844
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 18840 12804 18981 12832
rect 18840 12792 18846 12804
rect 18969 12801 18981 12804
rect 19015 12801 19027 12835
rect 19150 12832 19156 12844
rect 19111 12804 19156 12832
rect 18969 12795 19027 12801
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19260 12832 19288 12872
rect 20162 12860 20168 12912
rect 20220 12900 20226 12912
rect 20220 12872 21404 12900
rect 20220 12860 20226 12872
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 19260 12804 20637 12832
rect 20625 12801 20637 12804
rect 20671 12832 20683 12835
rect 21174 12832 21180 12844
rect 20671 12804 21180 12832
rect 20671 12801 20683 12804
rect 20625 12795 20683 12801
rect 21174 12792 21180 12804
rect 21232 12792 21238 12844
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18230 12764 18236 12776
rect 17911 12736 18236 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 20346 12696 20352 12708
rect 3099 12668 20352 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 20346 12656 20352 12668
rect 20404 12656 20410 12708
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12628 17371 12631
rect 19334 12628 19340 12640
rect 17359 12600 19340 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 19613 12631 19671 12637
rect 19613 12597 19625 12631
rect 19659 12628 19671 12631
rect 19978 12628 19984 12640
rect 19659 12600 19984 12628
rect 19659 12597 19671 12600
rect 19613 12591 19671 12597
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20530 12628 20536 12640
rect 20491 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 21284 12628 21312 12795
rect 21376 12764 21404 12872
rect 22186 12860 22192 12912
rect 22244 12900 22250 12912
rect 22557 12903 22615 12909
rect 22557 12900 22569 12903
rect 22244 12872 22569 12900
rect 22244 12860 22250 12872
rect 22557 12869 22569 12872
rect 22603 12869 22615 12903
rect 22557 12863 22615 12869
rect 22649 12903 22707 12909
rect 22649 12869 22661 12903
rect 22695 12900 22707 12903
rect 23474 12900 23480 12912
rect 22695 12872 23480 12900
rect 22695 12869 22707 12872
rect 22649 12863 22707 12869
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 23845 12903 23903 12909
rect 23845 12869 23857 12903
rect 23891 12900 23903 12903
rect 25332 12900 25360 12940
rect 28537 12937 28549 12940
rect 28583 12937 28595 12971
rect 28537 12931 28595 12937
rect 23891 12872 25360 12900
rect 25409 12903 25467 12909
rect 23891 12869 23903 12872
rect 23845 12863 23903 12869
rect 25409 12869 25421 12903
rect 25455 12900 25467 12903
rect 27154 12900 27160 12912
rect 25455 12872 27160 12900
rect 25455 12869 25467 12872
rect 25409 12863 25467 12869
rect 27154 12860 27160 12872
rect 27212 12860 27218 12912
rect 27433 12903 27491 12909
rect 27433 12869 27445 12903
rect 27479 12900 27491 12903
rect 28258 12900 28264 12912
rect 27479 12872 28264 12900
rect 27479 12869 27491 12872
rect 27433 12863 27491 12869
rect 28258 12860 28264 12872
rect 28316 12860 28322 12912
rect 28368 12872 29132 12900
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12801 26111 12835
rect 26053 12795 26111 12801
rect 22373 12767 22431 12773
rect 22373 12764 22385 12767
rect 21376 12736 22385 12764
rect 22373 12733 22385 12736
rect 22419 12733 22431 12767
rect 23750 12764 23756 12776
rect 23711 12736 23756 12764
rect 22373 12727 22431 12733
rect 22388 12696 22416 12727
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 24857 12767 24915 12773
rect 24857 12764 24869 12767
rect 23860 12736 24869 12764
rect 23860 12696 23888 12736
rect 24857 12733 24869 12736
rect 24903 12733 24915 12767
rect 24857 12727 24915 12733
rect 25501 12767 25559 12773
rect 25501 12733 25513 12767
rect 25547 12764 25559 12767
rect 25774 12764 25780 12776
rect 25547 12736 25780 12764
rect 25547 12733 25559 12736
rect 25501 12727 25559 12733
rect 25774 12724 25780 12736
rect 25832 12724 25838 12776
rect 24302 12696 24308 12708
rect 22388 12668 23888 12696
rect 24263 12668 24308 12696
rect 24302 12656 24308 12668
rect 24360 12656 24366 12708
rect 23842 12628 23848 12640
rect 21284 12600 23848 12628
rect 23842 12588 23848 12600
rect 23900 12628 23906 12640
rect 26068 12628 26096 12795
rect 26142 12792 26148 12844
rect 26200 12832 26206 12844
rect 27985 12835 28043 12841
rect 26200 12804 26245 12832
rect 26200 12792 26206 12804
rect 27985 12801 27997 12835
rect 28031 12832 28043 12835
rect 28074 12832 28080 12844
rect 28031 12804 28080 12832
rect 28031 12801 28043 12804
rect 27985 12795 28043 12801
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 26602 12724 26608 12776
rect 26660 12764 26666 12776
rect 27341 12767 27399 12773
rect 27341 12764 27353 12767
rect 26660 12736 27353 12764
rect 26660 12724 26666 12736
rect 27341 12733 27353 12736
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 27430 12724 27436 12776
rect 27488 12764 27494 12776
rect 28368 12764 28396 12872
rect 29104 12841 29132 12872
rect 28629 12835 28687 12841
rect 28629 12801 28641 12835
rect 28675 12801 28687 12835
rect 28629 12795 28687 12801
rect 29089 12835 29147 12841
rect 29089 12801 29101 12835
rect 29135 12801 29147 12835
rect 29089 12795 29147 12801
rect 27488 12736 28396 12764
rect 28644 12764 28672 12795
rect 29178 12764 29184 12776
rect 28644 12736 29184 12764
rect 27488 12724 27494 12736
rect 29178 12724 29184 12736
rect 29236 12724 29242 12776
rect 27706 12656 27712 12708
rect 27764 12696 27770 12708
rect 29086 12696 29092 12708
rect 27764 12668 29092 12696
rect 27764 12656 27770 12668
rect 29086 12656 29092 12668
rect 29144 12696 29150 12708
rect 29733 12699 29791 12705
rect 29733 12696 29745 12699
rect 29144 12668 29745 12696
rect 29144 12656 29150 12668
rect 29733 12665 29745 12668
rect 29779 12665 29791 12699
rect 29733 12659 29791 12665
rect 23900 12600 26096 12628
rect 23900 12588 23906 12600
rect 26142 12588 26148 12640
rect 26200 12628 26206 12640
rect 29181 12631 29239 12637
rect 29181 12628 29193 12631
rect 26200 12600 29193 12628
rect 26200 12588 26206 12600
rect 29181 12597 29193 12600
rect 29227 12597 29239 12631
rect 29181 12591 29239 12597
rect 1104 12538 36892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36892 12538
rect 1104 12464 36892 12486
rect 17678 12424 17684 12436
rect 17639 12396 17684 12424
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 20622 12424 20628 12436
rect 17788 12396 20116 12424
rect 20583 12396 20628 12424
rect 14458 12316 14464 12368
rect 14516 12356 14522 12368
rect 17788 12356 17816 12396
rect 14516 12328 17816 12356
rect 14516 12316 14522 12328
rect 18230 12316 18236 12368
rect 18288 12316 18294 12368
rect 18877 12359 18935 12365
rect 18877 12325 18889 12359
rect 18923 12356 18935 12359
rect 19797 12359 19855 12365
rect 19797 12356 19809 12359
rect 18923 12328 19809 12356
rect 18923 12325 18935 12328
rect 18877 12319 18935 12325
rect 19797 12325 19809 12328
rect 19843 12356 19855 12359
rect 19978 12356 19984 12368
rect 19843 12328 19984 12356
rect 19843 12325 19855 12328
rect 19797 12319 19855 12325
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 20088 12356 20116 12396
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 21174 12424 21180 12436
rect 21135 12396 21180 12424
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 23198 12424 23204 12436
rect 21284 12396 23204 12424
rect 21284 12356 21312 12396
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 24486 12384 24492 12436
rect 24544 12424 24550 12436
rect 27893 12427 27951 12433
rect 24544 12396 27108 12424
rect 24544 12384 24550 12396
rect 20088 12328 21312 12356
rect 21821 12359 21879 12365
rect 21821 12325 21833 12359
rect 21867 12356 21879 12359
rect 22922 12356 22928 12368
rect 21867 12328 22928 12356
rect 21867 12325 21879 12328
rect 21821 12319 21879 12325
rect 22922 12316 22928 12328
rect 22980 12356 22986 12368
rect 27080 12356 27108 12396
rect 27893 12393 27905 12427
rect 27939 12424 27951 12427
rect 27982 12424 27988 12436
rect 27939 12396 27988 12424
rect 27939 12393 27951 12396
rect 27893 12387 27951 12393
rect 27982 12384 27988 12396
rect 28040 12384 28046 12436
rect 28350 12384 28356 12436
rect 28408 12424 28414 12436
rect 28537 12427 28595 12433
rect 28537 12424 28549 12427
rect 28408 12396 28549 12424
rect 28408 12384 28414 12396
rect 28537 12393 28549 12396
rect 28583 12393 28595 12427
rect 29086 12424 29092 12436
rect 29047 12396 29092 12424
rect 28537 12387 28595 12393
rect 29086 12384 29092 12396
rect 29144 12384 29150 12436
rect 36170 12424 36176 12436
rect 31726 12396 36176 12424
rect 29733 12359 29791 12365
rect 29733 12356 29745 12359
rect 22980 12328 25728 12356
rect 27080 12328 29745 12356
rect 22980 12316 22986 12328
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 18046 12288 18052 12300
rect 12759 12260 18052 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18248 12288 18276 12316
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 18248 12260 19441 12288
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 22002 12248 22008 12300
rect 22060 12288 22066 12300
rect 22373 12291 22431 12297
rect 22373 12288 22385 12291
rect 22060 12260 22385 12288
rect 22060 12248 22066 12260
rect 22373 12257 22385 12260
rect 22419 12257 22431 12291
rect 23566 12288 23572 12300
rect 23479 12260 23572 12288
rect 22373 12251 22431 12257
rect 23566 12248 23572 12260
rect 23624 12288 23630 12300
rect 25700 12297 25728 12328
rect 29733 12325 29745 12328
rect 29779 12356 29791 12359
rect 31726 12356 31754 12396
rect 36170 12384 36176 12396
rect 36228 12384 36234 12436
rect 29779 12328 31754 12356
rect 29779 12325 29791 12328
rect 29733 12319 29791 12325
rect 24673 12291 24731 12297
rect 24673 12288 24685 12291
rect 23624 12260 24685 12288
rect 23624 12248 23630 12260
rect 24673 12257 24685 12260
rect 24719 12257 24731 12291
rect 24673 12251 24731 12257
rect 25685 12291 25743 12297
rect 25685 12257 25697 12291
rect 25731 12257 25743 12291
rect 25685 12251 25743 12257
rect 26697 12291 26755 12297
rect 26697 12257 26709 12291
rect 26743 12288 26755 12291
rect 27706 12288 27712 12300
rect 26743 12260 27712 12288
rect 26743 12257 26755 12260
rect 26697 12251 26755 12257
rect 27706 12248 27712 12260
rect 27764 12248 27770 12300
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12220 12679 12223
rect 13262 12220 13268 12232
rect 12667 12192 13268 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 18196 12192 18245 12220
rect 18196 12180 18202 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 17586 12112 17592 12164
rect 17644 12152 17650 12164
rect 18432 12152 18460 12183
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 19668 12192 19713 12220
rect 19668 12180 19674 12192
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20496 12192 20545 12220
rect 20496 12180 20502 12192
rect 20533 12189 20545 12192
rect 20579 12220 20591 12223
rect 21174 12220 21180 12232
rect 20579 12192 21180 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24544 12192 24777 12220
rect 24544 12180 24550 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 27338 12220 27344 12232
rect 27299 12192 27344 12220
rect 24765 12183 24823 12189
rect 27338 12180 27344 12192
rect 27396 12180 27402 12232
rect 27801 12223 27859 12229
rect 27801 12189 27813 12223
rect 27847 12220 27859 12223
rect 27890 12220 27896 12232
rect 27847 12192 27896 12220
rect 27847 12189 27859 12192
rect 27801 12183 27859 12189
rect 27890 12180 27896 12192
rect 27948 12180 27954 12232
rect 28626 12220 28632 12232
rect 28587 12192 28632 12220
rect 28626 12180 28632 12192
rect 28684 12220 28690 12232
rect 30377 12223 30435 12229
rect 30377 12220 30389 12223
rect 28684 12192 30389 12220
rect 28684 12180 28690 12192
rect 30377 12189 30389 12192
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 17644 12124 18460 12152
rect 17644 12112 17650 12124
rect 18506 12112 18512 12164
rect 18564 12152 18570 12164
rect 19058 12152 19064 12164
rect 18564 12124 19064 12152
rect 18564 12112 18570 12124
rect 19058 12112 19064 12124
rect 19116 12152 19122 12164
rect 21450 12152 21456 12164
rect 19116 12124 21456 12152
rect 19116 12112 19122 12124
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 22281 12155 22339 12161
rect 22281 12121 22293 12155
rect 22327 12121 22339 12155
rect 22922 12152 22928 12164
rect 22883 12124 22928 12152
rect 22281 12115 22339 12121
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 1912 12056 7941 12084
rect 1912 12044 1918 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 13262 12084 13268 12096
rect 13223 12056 13268 12084
rect 7929 12047 7987 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 19610 12084 19616 12096
rect 17552 12056 19616 12084
rect 17552 12044 17558 12056
rect 19610 12044 19616 12056
rect 19668 12044 19674 12096
rect 22296 12084 22324 12115
rect 22922 12112 22928 12124
rect 22980 12112 22986 12164
rect 23474 12152 23480 12164
rect 23435 12124 23480 12152
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 25777 12155 25835 12161
rect 25777 12121 25789 12155
rect 25823 12152 25835 12155
rect 29822 12152 29828 12164
rect 25823 12124 29828 12152
rect 25823 12121 25835 12124
rect 25777 12115 25835 12121
rect 29822 12112 29828 12124
rect 29880 12112 29886 12164
rect 27249 12087 27307 12093
rect 27249 12084 27261 12087
rect 22296 12056 27261 12084
rect 27249 12053 27261 12056
rect 27295 12053 27307 12087
rect 27249 12047 27307 12053
rect 27338 12044 27344 12096
rect 27396 12084 27402 12096
rect 28810 12084 28816 12096
rect 27396 12056 28816 12084
rect 27396 12044 27402 12056
rect 28810 12044 28816 12056
rect 28868 12044 28874 12096
rect 1104 11994 36892 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 36892 11994
rect 1104 11920 36892 11942
rect 17586 11880 17592 11892
rect 17547 11852 17592 11880
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 18138 11880 18144 11892
rect 18099 11852 18144 11880
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 21177 11883 21235 11889
rect 18248 11852 21036 11880
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 8168 11784 8309 11812
rect 8168 11772 8174 11784
rect 8297 11781 8309 11784
rect 8343 11812 8355 11815
rect 17034 11812 17040 11824
rect 8343 11784 17040 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 18248 11812 18276 11852
rect 17880 11784 18276 11812
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11744 14335 11747
rect 17681 11747 17739 11753
rect 14323 11716 14872 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14844 11617 14872 11716
rect 17681 11713 17693 11747
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17696 11676 17724 11707
rect 17880 11676 17908 11784
rect 18782 11772 18788 11824
rect 18840 11812 18846 11824
rect 20073 11815 20131 11821
rect 20073 11812 20085 11815
rect 18840 11784 20085 11812
rect 18840 11772 18846 11784
rect 20073 11781 20085 11784
rect 20119 11781 20131 11815
rect 20073 11775 20131 11781
rect 20346 11772 20352 11824
rect 20404 11812 20410 11824
rect 20622 11812 20628 11824
rect 20404 11784 20628 11812
rect 20404 11772 20410 11784
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 21008 11756 21036 11852
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 22186 11880 22192 11892
rect 21223 11852 22192 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 23293 11883 23351 11889
rect 23293 11849 23305 11883
rect 23339 11880 23351 11883
rect 23750 11880 23756 11892
rect 23339 11852 23756 11880
rect 23339 11849 23351 11852
rect 23293 11843 23351 11849
rect 23750 11840 23756 11852
rect 23808 11840 23814 11892
rect 26142 11880 26148 11892
rect 25056 11852 26148 11880
rect 22557 11815 22615 11821
rect 22557 11781 22569 11815
rect 22603 11812 22615 11815
rect 24670 11812 24676 11824
rect 22603 11784 24676 11812
rect 22603 11781 22615 11784
rect 22557 11775 22615 11781
rect 24670 11772 24676 11784
rect 24728 11772 24734 11824
rect 25056 11821 25084 11852
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 27154 11840 27160 11892
rect 27212 11880 27218 11892
rect 27249 11883 27307 11889
rect 27249 11880 27261 11883
rect 27212 11852 27261 11880
rect 27212 11840 27218 11852
rect 27249 11849 27261 11852
rect 27295 11849 27307 11883
rect 27249 11843 27307 11849
rect 27798 11840 27804 11892
rect 27856 11880 27862 11892
rect 28537 11883 28595 11889
rect 28537 11880 28549 11883
rect 27856 11852 28549 11880
rect 27856 11840 27862 11852
rect 28537 11849 28549 11852
rect 28583 11849 28595 11883
rect 29822 11880 29828 11892
rect 29783 11852 29828 11880
rect 28537 11843 28595 11849
rect 29822 11840 29828 11852
rect 29880 11840 29886 11892
rect 25041 11815 25099 11821
rect 25041 11781 25053 11815
rect 25087 11781 25099 11815
rect 25041 11775 25099 11781
rect 25130 11772 25136 11824
rect 25188 11812 25194 11824
rect 25188 11784 25233 11812
rect 25188 11772 25194 11784
rect 26050 11772 26056 11824
rect 26108 11812 26114 11824
rect 26237 11815 26295 11821
rect 26237 11812 26249 11815
rect 26108 11784 26249 11812
rect 26108 11772 26114 11784
rect 26237 11781 26249 11784
rect 26283 11781 26295 11815
rect 26237 11775 26295 11781
rect 27706 11772 27712 11824
rect 27764 11812 27770 11824
rect 27764 11784 31754 11812
rect 27764 11772 27770 11784
rect 18046 11704 18052 11756
rect 18104 11744 18110 11756
rect 18104 11716 19564 11744
rect 18104 11704 18110 11716
rect 17696 11648 17908 11676
rect 18138 11636 18144 11688
rect 18196 11676 18202 11688
rect 19245 11679 19303 11685
rect 19245 11676 19257 11679
rect 18196 11648 19257 11676
rect 18196 11636 18202 11648
rect 19245 11645 19257 11648
rect 19291 11645 19303 11679
rect 19245 11639 19303 11645
rect 19429 11679 19487 11685
rect 19429 11645 19441 11679
rect 19475 11645 19487 11679
rect 19536 11676 19564 11716
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 21048 11716 21097 11744
rect 21048 11704 21054 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 23198 11704 23204 11756
rect 23256 11744 23262 11756
rect 23385 11747 23443 11753
rect 23385 11744 23397 11747
rect 23256 11716 23397 11744
rect 23256 11704 23262 11716
rect 23385 11713 23397 11716
rect 23431 11713 23443 11747
rect 23385 11707 23443 11713
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 25685 11747 25743 11753
rect 25685 11744 25697 11747
rect 23716 11716 24348 11744
rect 23716 11704 23722 11716
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19536 11648 19993 11676
rect 19429 11639 19487 11645
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 19981 11639 20039 11645
rect 20364 11648 20637 11676
rect 14093 11611 14151 11617
rect 14093 11608 14105 11611
rect 6886 11580 14105 11608
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 6886 11540 6914 11580
rect 14093 11577 14105 11580
rect 14139 11577 14151 11611
rect 14093 11571 14151 11577
rect 14829 11611 14887 11617
rect 14829 11577 14841 11611
rect 14875 11608 14887 11611
rect 18874 11608 18880 11620
rect 14875 11580 18880 11608
rect 14875 11577 14887 11580
rect 14829 11571 14887 11577
rect 18874 11568 18880 11580
rect 18932 11568 18938 11620
rect 19444 11608 19472 11639
rect 20254 11608 20260 11620
rect 19444 11580 20260 11608
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 20364 11552 20392 11648
rect 20625 11645 20637 11648
rect 20671 11676 20683 11679
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 20671 11648 22385 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11676 22707 11679
rect 23750 11676 23756 11688
rect 22695 11648 23756 11676
rect 22695 11645 22707 11648
rect 22649 11639 22707 11645
rect 5592 11512 6914 11540
rect 19061 11543 19119 11549
rect 5592 11500 5598 11512
rect 19061 11509 19073 11543
rect 19107 11540 19119 11543
rect 19978 11540 19984 11552
rect 19107 11512 19984 11540
rect 19107 11509 19119 11512
rect 19061 11503 19119 11509
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20346 11500 20352 11552
rect 20404 11500 20410 11552
rect 21082 11500 21088 11552
rect 21140 11540 21146 11552
rect 21818 11540 21824 11552
rect 21140 11512 21824 11540
rect 21140 11500 21146 11512
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 22388 11540 22416 11639
rect 23750 11636 23756 11648
rect 23808 11636 23814 11688
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11645 24179 11679
rect 24320 11676 24348 11716
rect 25332 11716 25697 11744
rect 25332 11676 25360 11716
rect 25685 11713 25697 11716
rect 25731 11713 25743 11747
rect 26878 11744 26884 11756
rect 25685 11707 25743 11713
rect 26528 11716 26884 11744
rect 24320 11648 25360 11676
rect 26329 11679 26387 11685
rect 24121 11639 24179 11645
rect 26329 11645 26341 11679
rect 26375 11676 26387 11679
rect 26528 11676 26556 11716
rect 26878 11704 26884 11716
rect 26936 11704 26942 11756
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 27522 11744 27528 11756
rect 27387 11716 27528 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 27522 11704 27528 11716
rect 27580 11704 27586 11756
rect 27798 11744 27804 11756
rect 27759 11716 27804 11744
rect 27798 11704 27804 11716
rect 27856 11704 27862 11756
rect 28445 11747 28503 11753
rect 28445 11713 28457 11747
rect 28491 11744 28503 11747
rect 28534 11744 28540 11756
rect 28491 11716 28540 11744
rect 28491 11713 28503 11716
rect 28445 11707 28503 11713
rect 28534 11704 28540 11716
rect 28592 11704 28598 11756
rect 29089 11747 29147 11753
rect 29089 11713 29101 11747
rect 29135 11744 29147 11747
rect 29178 11744 29184 11756
rect 29135 11716 29184 11744
rect 29135 11713 29147 11716
rect 29089 11707 29147 11713
rect 29178 11704 29184 11716
rect 29236 11704 29242 11756
rect 29730 11744 29736 11756
rect 29691 11716 29736 11744
rect 29730 11704 29736 11716
rect 29788 11704 29794 11756
rect 26375 11648 26556 11676
rect 26375 11645 26387 11648
rect 26329 11639 26387 11645
rect 22738 11568 22744 11620
rect 22796 11608 22802 11620
rect 24136 11608 24164 11639
rect 27614 11636 27620 11688
rect 27672 11676 27678 11688
rect 27893 11679 27951 11685
rect 27893 11676 27905 11679
rect 27672 11648 27905 11676
rect 27672 11636 27678 11648
rect 27893 11645 27905 11648
rect 27939 11645 27951 11679
rect 31726 11676 31754 11784
rect 35434 11676 35440 11688
rect 27893 11639 27951 11645
rect 28000 11648 28994 11676
rect 31726 11648 35440 11676
rect 22796 11580 24164 11608
rect 22796 11568 22802 11580
rect 25774 11568 25780 11620
rect 25832 11608 25838 11620
rect 28000 11608 28028 11648
rect 25832 11580 28028 11608
rect 28966 11608 28994 11648
rect 35434 11636 35440 11648
rect 35492 11636 35498 11688
rect 29181 11611 29239 11617
rect 29181 11608 29193 11611
rect 28966 11580 29193 11608
rect 25832 11568 25838 11580
rect 29181 11577 29193 11580
rect 29227 11577 29239 11611
rect 29181 11571 29239 11577
rect 24118 11540 24124 11552
rect 22388 11512 24124 11540
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24302 11500 24308 11552
rect 24360 11540 24366 11552
rect 27798 11540 27804 11552
rect 24360 11512 27804 11540
rect 24360 11500 24366 11512
rect 27798 11500 27804 11512
rect 27856 11500 27862 11552
rect 1104 11450 36892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36892 11450
rect 1104 11376 36892 11398
rect 17494 11336 17500 11348
rect 17455 11308 17500 11336
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 18874 11296 18880 11348
rect 18932 11336 18938 11348
rect 24486 11336 24492 11348
rect 18932 11308 24492 11336
rect 18932 11296 18938 11308
rect 24486 11296 24492 11308
rect 24544 11296 24550 11348
rect 24670 11336 24676 11348
rect 24631 11308 24676 11336
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 24762 11296 24768 11348
rect 24820 11336 24826 11348
rect 28902 11336 28908 11348
rect 24820 11308 28908 11336
rect 24820 11296 24826 11308
rect 28902 11296 28908 11308
rect 28960 11296 28966 11348
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 30469 11339 30527 11345
rect 30469 11336 30481 11339
rect 29052 11308 30481 11336
rect 29052 11296 29058 11308
rect 30469 11305 30481 11308
rect 30515 11305 30527 11339
rect 30469 11299 30527 11305
rect 18966 11228 18972 11280
rect 19024 11268 19030 11280
rect 19024 11240 21128 11268
rect 19024 11228 19030 11240
rect 19058 11200 19064 11212
rect 16960 11172 19064 11200
rect 1854 11132 1860 11144
rect 1815 11104 1860 11132
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 16960 11141 16988 11172
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19521 11203 19579 11209
rect 19521 11169 19533 11203
rect 19567 11200 19579 11203
rect 20162 11200 20168 11212
rect 19567 11172 20168 11200
rect 19567 11169 19579 11172
rect 19521 11163 19579 11169
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 21100 11209 21128 11240
rect 21358 11228 21364 11280
rect 21416 11268 21422 11280
rect 22002 11268 22008 11280
rect 21416 11240 22008 11268
rect 21416 11228 21422 11240
rect 21085 11203 21143 11209
rect 21085 11169 21097 11203
rect 21131 11169 21143 11203
rect 21726 11200 21732 11212
rect 21687 11172 21732 11200
rect 21085 11163 21143 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11101 17003 11135
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 16945 11095 17003 11101
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 18046 11132 18052 11144
rect 17959 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11132 18110 11144
rect 18506 11132 18512 11144
rect 18104 11104 18512 11132
rect 18104 11092 18110 11104
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 19334 11132 19340 11144
rect 18923 11104 19340 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 16853 11067 16911 11073
rect 16853 11033 16865 11067
rect 16899 11064 16911 11067
rect 19242 11064 19248 11076
rect 16899 11036 19248 11064
rect 16899 11033 16911 11036
rect 16853 11027 16911 11033
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 19613 11067 19671 11073
rect 19613 11033 19625 11067
rect 19659 11033 19671 11067
rect 20530 11064 20536 11076
rect 20491 11036 20536 11064
rect 19613 11027 19671 11033
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 19628 10996 19656 11027
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 21177 11067 21235 11073
rect 21177 11033 21189 11067
rect 21223 11064 21235 11067
rect 21836 11064 21864 11240
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 25314 11228 25320 11280
rect 25372 11268 25378 11280
rect 25372 11240 27108 11268
rect 25372 11228 25378 11240
rect 22922 11200 22928 11212
rect 22883 11172 22928 11200
rect 22922 11160 22928 11172
rect 22980 11160 22986 11212
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25777 11203 25835 11209
rect 25777 11200 25789 11203
rect 25280 11172 25789 11200
rect 25280 11160 25286 11172
rect 25777 11169 25789 11172
rect 25823 11200 25835 11203
rect 26142 11200 26148 11212
rect 25823 11172 26148 11200
rect 25823 11169 25835 11172
rect 25777 11163 25835 11169
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 27080 11209 27108 11240
rect 27065 11203 27123 11209
rect 27065 11169 27077 11203
rect 27111 11169 27123 11203
rect 27706 11200 27712 11212
rect 27667 11172 27712 11200
rect 27065 11163 27123 11169
rect 27706 11160 27712 11172
rect 27764 11160 27770 11212
rect 29825 11203 29883 11209
rect 29825 11200 29837 11203
rect 28000 11172 29837 11200
rect 23198 11092 23204 11144
rect 23256 11132 23262 11144
rect 23385 11135 23443 11141
rect 23385 11132 23397 11135
rect 23256 11104 23397 11132
rect 23256 11092 23262 11104
rect 23385 11101 23397 11104
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 24762 11132 24768 11144
rect 23808 11104 24768 11132
rect 23808 11092 23814 11104
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 22281 11067 22339 11073
rect 22281 11064 22293 11067
rect 21223 11036 21680 11064
rect 21836 11036 22293 11064
rect 21223 11033 21235 11036
rect 21177 11027 21235 11033
rect 19392 10968 19656 10996
rect 21652 10996 21680 11036
rect 22281 11033 22293 11036
rect 22327 11033 22339 11067
rect 22281 11027 22339 11033
rect 22373 11067 22431 11073
rect 22373 11033 22385 11067
rect 22419 11064 22431 11067
rect 23934 11064 23940 11076
rect 22419 11036 22876 11064
rect 22419 11033 22431 11036
rect 22373 11027 22431 11033
rect 22094 10996 22100 11008
rect 21652 10968 22100 10996
rect 19392 10956 19398 10968
rect 22094 10956 22100 10968
rect 22152 10956 22158 11008
rect 22848 10996 22876 11036
rect 23032 11036 23940 11064
rect 23032 10996 23060 11036
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 24026 11024 24032 11076
rect 24084 11024 24090 11076
rect 25498 11064 25504 11076
rect 25459 11036 25504 11064
rect 25498 11024 25504 11036
rect 25556 11024 25562 11076
rect 25593 11067 25651 11073
rect 25593 11033 25605 11067
rect 25639 11064 25651 11067
rect 25774 11064 25780 11076
rect 25639 11036 25780 11064
rect 25639 11033 25651 11036
rect 25593 11027 25651 11033
rect 25774 11024 25780 11036
rect 25832 11024 25838 11076
rect 27157 11067 27215 11073
rect 27157 11033 27169 11067
rect 27203 11064 27215 11067
rect 28000 11064 28028 11172
rect 29825 11169 29837 11172
rect 29871 11169 29883 11203
rect 29825 11163 29883 11169
rect 28534 11132 28540 11144
rect 28495 11104 28540 11132
rect 28534 11092 28540 11104
rect 28592 11092 28598 11144
rect 29917 11135 29975 11141
rect 29917 11101 29929 11135
rect 29963 11101 29975 11135
rect 29917 11095 29975 11101
rect 27203 11036 28028 11064
rect 29932 11064 29960 11095
rect 30098 11092 30104 11144
rect 30156 11132 30162 11144
rect 30377 11135 30435 11141
rect 30377 11132 30389 11135
rect 30156 11104 30389 11132
rect 30156 11092 30162 11104
rect 30377 11101 30389 11104
rect 30423 11101 30435 11135
rect 36078 11132 36084 11144
rect 36039 11104 36084 11132
rect 30377 11095 30435 11101
rect 36078 11092 36084 11104
rect 36136 11092 36142 11144
rect 31478 11064 31484 11076
rect 29932 11036 31484 11064
rect 27203 11033 27215 11036
rect 27157 11027 27215 11033
rect 31478 11024 31484 11036
rect 31536 11024 31542 11076
rect 35621 11067 35679 11073
rect 35621 11033 35633 11067
rect 35667 11064 35679 11067
rect 36262 11064 36268 11076
rect 35667 11036 36268 11064
rect 35667 11033 35679 11036
rect 35621 11027 35679 11033
rect 36262 11024 36268 11036
rect 36320 11024 36326 11076
rect 22848 10968 23060 10996
rect 23569 10999 23627 11005
rect 23569 10965 23581 10999
rect 23615 10996 23627 10999
rect 24044 10996 24072 11024
rect 23615 10968 24072 10996
rect 23615 10965 23627 10968
rect 23569 10959 23627 10965
rect 27614 10956 27620 11008
rect 27672 10996 27678 11008
rect 28629 10999 28687 11005
rect 28629 10996 28641 10999
rect 27672 10968 28641 10996
rect 27672 10956 27678 10968
rect 28629 10965 28641 10968
rect 28675 10965 28687 10999
rect 28629 10959 28687 10965
rect 1104 10906 36892 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 36892 10906
rect 1104 10832 36892 10854
rect 17405 10795 17463 10801
rect 17405 10761 17417 10795
rect 17451 10792 17463 10795
rect 18046 10792 18052 10804
rect 17451 10764 18052 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19576 10764 20392 10792
rect 19576 10752 19582 10764
rect 18138 10684 18144 10736
rect 18196 10724 18202 10736
rect 18693 10727 18751 10733
rect 18693 10724 18705 10727
rect 18196 10696 18705 10724
rect 18196 10684 18202 10696
rect 18693 10693 18705 10696
rect 18739 10693 18751 10727
rect 18693 10687 18751 10693
rect 19242 10684 19248 10736
rect 19300 10724 19306 10736
rect 20257 10727 20315 10733
rect 20257 10724 20269 10727
rect 19300 10696 20269 10724
rect 19300 10684 19306 10696
rect 20257 10693 20269 10696
rect 20303 10693 20315 10727
rect 20364 10724 20392 10764
rect 21726 10752 21732 10804
rect 21784 10792 21790 10804
rect 28813 10795 28871 10801
rect 28813 10792 28825 10795
rect 21784 10764 25820 10792
rect 21784 10752 21790 10764
rect 22005 10727 22063 10733
rect 22005 10724 22017 10727
rect 20364 10696 22017 10724
rect 20257 10687 20315 10693
rect 22005 10693 22017 10696
rect 22051 10693 22063 10727
rect 22005 10687 22063 10693
rect 22925 10727 22983 10733
rect 22925 10693 22937 10727
rect 22971 10724 22983 10727
rect 23290 10724 23296 10736
rect 22971 10696 23296 10724
rect 22971 10693 22983 10696
rect 22925 10687 22983 10693
rect 23290 10684 23296 10696
rect 23348 10684 23354 10736
rect 24486 10724 24492 10736
rect 24447 10696 24492 10724
rect 24486 10684 24492 10696
rect 24544 10684 24550 10736
rect 25792 10733 25820 10764
rect 25884 10764 28825 10792
rect 25884 10733 25912 10764
rect 28813 10761 28825 10764
rect 28859 10761 28871 10795
rect 28813 10755 28871 10761
rect 30006 10752 30012 10804
rect 30064 10792 30070 10804
rect 30101 10795 30159 10801
rect 30101 10792 30113 10795
rect 30064 10764 30113 10792
rect 30064 10752 30070 10764
rect 30101 10761 30113 10764
rect 30147 10761 30159 10795
rect 30101 10755 30159 10761
rect 25777 10727 25835 10733
rect 25777 10693 25789 10727
rect 25823 10693 25835 10727
rect 25777 10687 25835 10693
rect 25869 10727 25927 10733
rect 25869 10693 25881 10727
rect 25915 10693 25927 10727
rect 25869 10687 25927 10693
rect 26142 10684 26148 10736
rect 26200 10724 26206 10736
rect 27249 10727 27307 10733
rect 27249 10724 27261 10727
rect 26200 10696 27261 10724
rect 26200 10684 26206 10696
rect 27249 10693 27261 10696
rect 27295 10693 27307 10727
rect 27249 10687 27307 10693
rect 27341 10727 27399 10733
rect 27341 10693 27353 10727
rect 27387 10724 27399 10727
rect 27890 10724 27896 10736
rect 27387 10696 27896 10724
rect 27387 10693 27399 10696
rect 27341 10687 27399 10693
rect 27890 10684 27896 10696
rect 27948 10684 27954 10736
rect 28074 10684 28080 10736
rect 28132 10724 28138 10736
rect 29457 10727 29515 10733
rect 29457 10724 29469 10727
rect 28132 10696 29469 10724
rect 28132 10684 28138 10696
rect 29457 10693 29469 10696
rect 29503 10693 29515 10727
rect 29457 10687 29515 10693
rect 17862 10656 17868 10668
rect 17823 10628 17868 10656
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 28626 10616 28632 10668
rect 28684 10656 28690 10668
rect 28905 10659 28963 10665
rect 28905 10656 28917 10659
rect 28684 10628 28917 10656
rect 28684 10616 28690 10628
rect 28905 10625 28917 10628
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 28994 10616 29000 10668
rect 29052 10656 29058 10668
rect 29549 10659 29607 10665
rect 29549 10656 29561 10659
rect 29052 10628 29561 10656
rect 29052 10616 29058 10628
rect 29549 10625 29561 10628
rect 29595 10625 29607 10659
rect 29549 10619 29607 10625
rect 30009 10659 30067 10665
rect 30009 10625 30021 10659
rect 30055 10625 30067 10659
rect 30009 10619 30067 10625
rect 18601 10591 18659 10597
rect 18601 10557 18613 10591
rect 18647 10588 18659 10591
rect 19426 10588 19432 10600
rect 18647 10560 19432 10588
rect 18647 10557 18659 10560
rect 18601 10551 18659 10557
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 19610 10588 19616 10600
rect 19571 10560 19616 10588
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 20036 10560 20177 10588
rect 20036 10548 20042 10560
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 20806 10548 20812 10600
rect 20864 10588 20870 10600
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 20864 10560 21189 10588
rect 20864 10548 20870 10560
rect 21177 10557 21189 10560
rect 21223 10588 21235 10591
rect 22738 10588 22744 10600
rect 21223 10560 22744 10588
rect 21223 10557 21235 10560
rect 21177 10551 21235 10557
rect 22738 10548 22744 10560
rect 22796 10548 22802 10600
rect 23014 10588 23020 10600
rect 22975 10560 23020 10588
rect 23014 10548 23020 10560
rect 23072 10548 23078 10600
rect 23290 10548 23296 10600
rect 23348 10588 23354 10600
rect 23569 10591 23627 10597
rect 23569 10588 23581 10591
rect 23348 10560 23581 10588
rect 23348 10548 23354 10560
rect 23569 10557 23581 10560
rect 23615 10557 23627 10591
rect 23569 10551 23627 10557
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 23716 10560 24593 10588
rect 23716 10548 23722 10560
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 24762 10548 24768 10600
rect 24820 10588 24826 10600
rect 26970 10588 26976 10600
rect 24820 10560 26976 10588
rect 24820 10548 24826 10560
rect 26970 10548 26976 10560
rect 27028 10548 27034 10600
rect 27706 10588 27712 10600
rect 27667 10560 27712 10588
rect 27706 10548 27712 10560
rect 27764 10548 27770 10600
rect 29270 10548 29276 10600
rect 29328 10588 29334 10600
rect 30024 10588 30052 10619
rect 29328 10560 30052 10588
rect 29328 10548 29334 10560
rect 6086 10480 6092 10532
rect 6144 10520 6150 10532
rect 19628 10520 19656 10548
rect 26329 10523 26387 10529
rect 6144 10492 19656 10520
rect 23676 10492 25268 10520
rect 6144 10480 6150 10492
rect 17957 10455 18015 10461
rect 17957 10421 17969 10455
rect 18003 10452 18015 10455
rect 18966 10452 18972 10464
rect 18003 10424 18972 10452
rect 18003 10421 18015 10424
rect 17957 10415 18015 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19242 10412 19248 10464
rect 19300 10452 19306 10464
rect 22830 10452 22836 10464
rect 19300 10424 22836 10452
rect 19300 10412 19306 10424
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 23290 10412 23296 10464
rect 23348 10452 23354 10464
rect 23676 10452 23704 10492
rect 23348 10424 23704 10452
rect 23348 10412 23354 10424
rect 25038 10412 25044 10464
rect 25096 10452 25102 10464
rect 25133 10455 25191 10461
rect 25133 10452 25145 10455
rect 25096 10424 25145 10452
rect 25096 10412 25102 10424
rect 25133 10421 25145 10424
rect 25179 10421 25191 10455
rect 25240 10452 25268 10492
rect 26329 10489 26341 10523
rect 26375 10520 26387 10523
rect 26418 10520 26424 10532
rect 26375 10492 26424 10520
rect 26375 10489 26387 10492
rect 26329 10483 26387 10489
rect 26418 10480 26424 10492
rect 26476 10520 26482 10532
rect 28442 10520 28448 10532
rect 26476 10492 28448 10520
rect 26476 10480 26482 10492
rect 28442 10480 28448 10492
rect 28500 10480 28506 10532
rect 27614 10452 27620 10464
rect 25240 10424 27620 10452
rect 25133 10415 25191 10421
rect 27614 10412 27620 10424
rect 27672 10412 27678 10464
rect 36357 10455 36415 10461
rect 36357 10421 36369 10455
rect 36403 10452 36415 10455
rect 36538 10452 36544 10464
rect 36403 10424 36544 10452
rect 36403 10421 36415 10424
rect 36357 10415 36415 10421
rect 36538 10412 36544 10424
rect 36596 10412 36602 10464
rect 1104 10362 36892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36892 10362
rect 1104 10288 36892 10310
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 5684 10220 7573 10248
rect 5684 10208 5690 10220
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 18138 10248 18144 10260
rect 18099 10220 18144 10248
rect 7561 10211 7619 10217
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 19334 10248 19340 10260
rect 18831 10220 19340 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 21634 10248 21640 10260
rect 19668 10220 21640 10248
rect 19668 10208 19674 10220
rect 21634 10208 21640 10220
rect 21692 10208 21698 10260
rect 23106 10208 23112 10260
rect 23164 10248 23170 10260
rect 24762 10248 24768 10260
rect 23164 10220 24768 10248
rect 23164 10208 23170 10220
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 25317 10251 25375 10257
rect 25317 10217 25329 10251
rect 25363 10248 25375 10251
rect 25498 10248 25504 10260
rect 25363 10220 25504 10248
rect 25363 10217 25375 10220
rect 25317 10211 25375 10217
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 26234 10208 26240 10260
rect 26292 10248 26298 10260
rect 27709 10251 27767 10257
rect 27709 10248 27721 10251
rect 26292 10220 27721 10248
rect 26292 10208 26298 10220
rect 27709 10217 27721 10220
rect 27755 10217 27767 10251
rect 27709 10211 27767 10217
rect 28258 10208 28264 10260
rect 28316 10248 28322 10260
rect 28353 10251 28411 10257
rect 28353 10248 28365 10251
rect 28316 10220 28365 10248
rect 28316 10208 28322 10220
rect 28353 10217 28365 10220
rect 28399 10217 28411 10251
rect 28353 10211 28411 10217
rect 18248 10152 19334 10180
rect 18248 10053 18276 10152
rect 19306 10124 19334 10152
rect 22186 10140 22192 10192
rect 22244 10180 22250 10192
rect 22922 10180 22928 10192
rect 22244 10152 22928 10180
rect 22244 10140 22250 10152
rect 22922 10140 22928 10152
rect 22980 10140 22986 10192
rect 26418 10180 26424 10192
rect 26379 10152 26424 10180
rect 26418 10140 26424 10152
rect 26476 10140 26482 10192
rect 26970 10180 26976 10192
rect 26931 10152 26976 10180
rect 26970 10140 26976 10152
rect 27028 10140 27034 10192
rect 19306 10084 19340 10124
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 22462 10112 22468 10124
rect 19536 10084 22468 10112
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 18233 10047 18291 10053
rect 7699 10016 8248 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 8220 9985 8248 10016
rect 18233 10013 18245 10047
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19536 10044 19564 10084
rect 22462 10072 22468 10084
rect 22520 10072 22526 10124
rect 22830 10112 22836 10124
rect 22791 10084 22836 10112
rect 22830 10072 22836 10084
rect 22888 10072 22894 10124
rect 23014 10072 23020 10124
rect 23072 10112 23078 10124
rect 23109 10115 23167 10121
rect 23109 10112 23121 10115
rect 23072 10084 23121 10112
rect 23072 10072 23078 10084
rect 23109 10081 23121 10084
rect 23155 10081 23167 10115
rect 23109 10075 23167 10081
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23937 10115 23995 10121
rect 23937 10112 23949 10115
rect 23256 10084 23949 10112
rect 23256 10072 23262 10084
rect 23937 10081 23949 10084
rect 23983 10081 23995 10115
rect 36081 10115 36139 10121
rect 36081 10112 36093 10115
rect 23937 10075 23995 10081
rect 25332 10084 36093 10112
rect 25332 10053 25360 10084
rect 27172 10053 27200 10084
rect 36081 10081 36093 10084
rect 36127 10081 36139 10115
rect 36081 10075 36139 10081
rect 18923 10016 19564 10044
rect 25317 10047 25375 10053
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 25317 10013 25329 10047
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10013 27215 10047
rect 27614 10044 27620 10056
rect 27575 10016 27620 10044
rect 27157 10007 27215 10013
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 28350 10004 28356 10056
rect 28408 10044 28414 10056
rect 28445 10047 28503 10053
rect 28445 10044 28457 10047
rect 28408 10016 28457 10044
rect 28408 10004 28414 10016
rect 28445 10013 28457 10016
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 29089 10047 29147 10053
rect 29089 10013 29101 10047
rect 29135 10044 29147 10047
rect 29454 10044 29460 10056
rect 29135 10016 29460 10044
rect 29135 10013 29147 10016
rect 29089 10007 29147 10013
rect 29454 10004 29460 10016
rect 29512 10004 29518 10056
rect 36354 10044 36360 10056
rect 36315 10016 36360 10044
rect 36354 10004 36360 10016
rect 36412 10004 36418 10056
rect 8205 9979 8263 9985
rect 8205 9945 8217 9979
rect 8251 9976 8263 9979
rect 19334 9976 19340 9988
rect 8251 9948 19340 9976
rect 8251 9945 8263 9948
rect 8205 9939 8263 9945
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9945 19763 9979
rect 19705 9939 19763 9945
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 19978 9976 19984 9988
rect 19843 9948 19984 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 17589 9911 17647 9917
rect 17589 9877 17601 9911
rect 17635 9908 17647 9911
rect 17862 9908 17868 9920
rect 17635 9880 17868 9908
rect 17635 9877 17647 9880
rect 17589 9871 17647 9877
rect 17862 9868 17868 9880
rect 17920 9908 17926 9920
rect 19610 9908 19616 9920
rect 17920 9880 19616 9908
rect 17920 9868 17926 9880
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 19720 9908 19748 9939
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 20530 9936 20536 9988
rect 20588 9976 20594 9988
rect 20717 9979 20775 9985
rect 20717 9976 20729 9979
rect 20588 9948 20729 9976
rect 20588 9936 20594 9948
rect 20717 9945 20729 9948
rect 20763 9945 20775 9979
rect 20717 9939 20775 9945
rect 21637 9979 21695 9985
rect 21637 9945 21649 9979
rect 21683 9945 21695 9979
rect 21637 9939 21695 9945
rect 20162 9908 20168 9920
rect 19720 9880 20168 9908
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 20254 9868 20260 9920
rect 20312 9908 20318 9920
rect 21652 9908 21680 9939
rect 21726 9936 21732 9988
rect 21784 9976 21790 9988
rect 22934 9979 22992 9985
rect 21784 9948 21829 9976
rect 21784 9936 21790 9948
rect 22934 9945 22946 9979
rect 22980 9976 22992 9979
rect 22980 9948 23060 9976
rect 22980 9945 22992 9948
rect 22934 9939 22992 9945
rect 20312 9880 21680 9908
rect 23032 9908 23060 9948
rect 24118 9936 24124 9988
rect 24176 9976 24182 9988
rect 25869 9979 25927 9985
rect 25869 9976 25881 9979
rect 24176 9948 25881 9976
rect 24176 9936 24182 9948
rect 25869 9945 25881 9948
rect 25915 9945 25927 9979
rect 25869 9939 25927 9945
rect 25970 9979 26028 9985
rect 25970 9945 25982 9979
rect 26016 9976 26028 9979
rect 28997 9979 29055 9985
rect 28997 9976 29009 9979
rect 26016 9948 29009 9976
rect 26016 9945 26028 9948
rect 25970 9939 26028 9945
rect 28997 9945 29009 9948
rect 29043 9945 29055 9979
rect 28997 9939 29055 9945
rect 24670 9908 24676 9920
rect 23032 9880 24676 9908
rect 20312 9868 20318 9880
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 34977 9911 35035 9917
rect 34977 9877 34989 9911
rect 35023 9908 35035 9911
rect 35618 9908 35624 9920
rect 35023 9880 35624 9908
rect 35023 9877 35035 9880
rect 34977 9871 35035 9877
rect 35618 9868 35624 9880
rect 35676 9868 35682 9920
rect 1104 9818 36892 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 36892 9818
rect 1104 9744 36892 9766
rect 19426 9704 19432 9716
rect 19339 9676 19432 9704
rect 19426 9664 19432 9676
rect 19484 9704 19490 9716
rect 20070 9704 20076 9716
rect 19484 9676 20076 9704
rect 19484 9664 19490 9676
rect 20070 9664 20076 9676
rect 20128 9664 20134 9716
rect 20714 9664 20720 9716
rect 20772 9664 20778 9716
rect 21726 9664 21732 9716
rect 21784 9704 21790 9716
rect 23290 9704 23296 9716
rect 21784 9676 23296 9704
rect 21784 9664 21790 9676
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 23566 9664 23572 9716
rect 23624 9704 23630 9716
rect 23624 9676 25912 9704
rect 23624 9664 23630 9676
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 17589 9639 17647 9645
rect 17589 9636 17601 9639
rect 12860 9608 17601 9636
rect 12860 9596 12866 9608
rect 17589 9605 17601 9608
rect 17635 9636 17647 9639
rect 17635 9608 19104 9636
rect 17635 9605 17647 9608
rect 17589 9599 17647 9605
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 17175 9540 18153 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 18141 9537 18153 9540
rect 18187 9568 18199 9571
rect 18966 9568 18972 9580
rect 18187 9540 18736 9568
rect 18927 9540 18972 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18708 9432 18736 9540
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 19076 9568 19104 9608
rect 19150 9596 19156 9648
rect 19208 9636 19214 9648
rect 20165 9639 20223 9645
rect 20165 9636 20177 9639
rect 19208 9608 20177 9636
rect 19208 9596 19214 9608
rect 20165 9605 20177 9608
rect 20211 9605 20223 9639
rect 20165 9599 20223 9605
rect 20257 9639 20315 9645
rect 20257 9605 20269 9639
rect 20303 9636 20315 9639
rect 20732 9636 20760 9664
rect 20303 9608 20760 9636
rect 20809 9639 20867 9645
rect 20303 9605 20315 9608
rect 20257 9599 20315 9605
rect 20809 9605 20821 9639
rect 20855 9636 20867 9639
rect 22554 9636 22560 9648
rect 20855 9608 22560 9636
rect 20855 9605 20867 9608
rect 20809 9599 20867 9605
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 24762 9636 24768 9648
rect 23506 9608 24768 9636
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 25884 9636 25912 9676
rect 27724 9676 28028 9704
rect 26513 9639 26571 9645
rect 26513 9636 26525 9639
rect 25714 9608 25820 9636
rect 25884 9608 26525 9636
rect 21269 9571 21327 9577
rect 19076 9540 20024 9568
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 19996 9500 20024 9540
rect 21269 9537 21281 9571
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 21284 9500 21312 9531
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 21416 9540 21461 9568
rect 21416 9528 21422 9540
rect 21542 9500 21548 9512
rect 18840 9472 18885 9500
rect 19996 9472 21548 9500
rect 18840 9460 18846 9472
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 22002 9500 22008 9512
rect 21963 9472 22008 9500
rect 22002 9460 22008 9472
rect 22060 9460 22066 9512
rect 22281 9503 22339 9509
rect 22281 9500 22293 9503
rect 22112 9472 22293 9500
rect 21910 9432 21916 9444
rect 18708 9404 21916 9432
rect 21910 9392 21916 9404
rect 21968 9392 21974 9444
rect 18233 9367 18291 9373
rect 18233 9333 18245 9367
rect 18279 9364 18291 9367
rect 18414 9364 18420 9376
rect 18279 9336 18420 9364
rect 18279 9333 18291 9336
rect 18233 9327 18291 9333
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 22112 9364 22140 9472
rect 22281 9469 22293 9472
rect 22327 9500 22339 9503
rect 22646 9500 22652 9512
rect 22327 9472 22652 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 22646 9460 22652 9472
rect 22704 9460 22710 9512
rect 24210 9500 24216 9512
rect 24171 9472 24216 9500
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 24489 9503 24547 9509
rect 24489 9500 24501 9503
rect 24320 9472 24501 9500
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 24320 9432 24348 9472
rect 24489 9469 24501 9472
rect 24535 9469 24547 9503
rect 25792 9500 25820 9608
rect 26513 9605 26525 9608
rect 26559 9605 26571 9639
rect 26513 9599 26571 9605
rect 26786 9596 26792 9648
rect 26844 9636 26850 9648
rect 27724 9636 27752 9676
rect 27890 9636 27896 9648
rect 26844 9608 27752 9636
rect 27851 9608 27896 9636
rect 26844 9596 26850 9608
rect 27890 9596 27896 9608
rect 27948 9596 27954 9648
rect 28000 9636 28028 9676
rect 31018 9636 31024 9648
rect 28000 9608 31024 9636
rect 31018 9596 31024 9608
rect 31076 9596 31082 9648
rect 36354 9636 36360 9648
rect 36315 9608 36360 9636
rect 36354 9596 36360 9608
rect 36412 9596 36418 9648
rect 26613 9571 26671 9577
rect 26613 9537 26625 9571
rect 26659 9568 26671 9571
rect 27062 9568 27068 9580
rect 26659 9540 27068 9568
rect 26659 9537 26671 9540
rect 26613 9531 26671 9537
rect 27062 9528 27068 9540
rect 27120 9528 27126 9580
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 27212 9540 27257 9568
rect 27212 9528 27218 9540
rect 27430 9528 27436 9580
rect 27488 9568 27494 9580
rect 27985 9571 28043 9577
rect 27985 9568 27997 9571
rect 27488 9540 27997 9568
rect 27488 9528 27494 9540
rect 27985 9537 27997 9540
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 32766 9500 32772 9512
rect 25792 9472 32772 9500
rect 24489 9463 24547 9469
rect 32766 9460 32772 9472
rect 32824 9460 32830 9512
rect 27249 9435 27307 9441
rect 27249 9432 27261 9435
rect 23624 9404 24348 9432
rect 23624 9392 23630 9404
rect 24320 9376 24348 9404
rect 25516 9404 27261 9432
rect 23750 9364 23756 9376
rect 19116 9336 22140 9364
rect 23711 9336 23756 9364
rect 19116 9324 19122 9336
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 24302 9324 24308 9376
rect 24360 9324 24366 9376
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 25516 9364 25544 9404
rect 27249 9401 27261 9404
rect 27295 9401 27307 9435
rect 27249 9395 27307 9401
rect 28537 9435 28595 9441
rect 28537 9401 28549 9435
rect 28583 9432 28595 9435
rect 29178 9432 29184 9444
rect 28583 9404 29184 9432
rect 28583 9401 28595 9404
rect 28537 9395 28595 9401
rect 29178 9392 29184 9404
rect 29236 9392 29242 9444
rect 32306 9392 32312 9444
rect 32364 9432 32370 9444
rect 32364 9404 33824 9432
rect 32364 9392 32370 9404
rect 25958 9364 25964 9376
rect 24728 9336 25544 9364
rect 25919 9336 25964 9364
rect 24728 9324 24734 9336
rect 25958 9324 25964 9336
rect 26016 9364 26022 9376
rect 27154 9364 27160 9376
rect 26016 9336 27160 9364
rect 26016 9324 26022 9336
rect 27154 9324 27160 9336
rect 27212 9324 27218 9376
rect 28442 9324 28448 9376
rect 28500 9364 28506 9376
rect 28997 9367 29055 9373
rect 28997 9364 29009 9367
rect 28500 9336 29009 9364
rect 28500 9324 28506 9336
rect 28997 9333 29009 9336
rect 29043 9333 29055 9367
rect 28997 9327 29055 9333
rect 32858 9324 32864 9376
rect 32916 9364 32922 9376
rect 33796 9373 33824 9404
rect 33045 9367 33103 9373
rect 33045 9364 33057 9367
rect 32916 9336 33057 9364
rect 32916 9324 32922 9336
rect 33045 9333 33057 9336
rect 33091 9333 33103 9367
rect 33045 9327 33103 9333
rect 33781 9367 33839 9373
rect 33781 9333 33793 9367
rect 33827 9364 33839 9367
rect 34241 9367 34299 9373
rect 34241 9364 34253 9367
rect 33827 9336 34253 9364
rect 33827 9333 33839 9336
rect 33781 9327 33839 9333
rect 34241 9333 34253 9336
rect 34287 9333 34299 9367
rect 34241 9327 34299 9333
rect 34790 9324 34796 9376
rect 34848 9364 34854 9376
rect 35161 9367 35219 9373
rect 35161 9364 35173 9367
rect 34848 9336 35173 9364
rect 34848 9324 34854 9336
rect 35161 9333 35173 9336
rect 35207 9333 35219 9367
rect 35161 9327 35219 9333
rect 35805 9367 35863 9373
rect 35805 9333 35817 9367
rect 35851 9364 35863 9367
rect 36170 9364 36176 9376
rect 35851 9336 36176 9364
rect 35851 9333 35863 9336
rect 35805 9327 35863 9333
rect 36170 9324 36176 9336
rect 36228 9324 36234 9376
rect 1104 9274 36892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36892 9274
rect 1104 9200 36892 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 6546 9160 6552 9172
rect 2455 9132 6552 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 2424 8956 2452 9123
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19426 9160 19432 9172
rect 18923 9132 19432 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 20254 9120 20260 9172
rect 20312 9160 20318 9172
rect 20438 9160 20444 9172
rect 20312 9132 20444 9160
rect 20312 9120 20318 9132
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 22186 9160 22192 9172
rect 21560 9132 22192 9160
rect 17586 9052 17592 9104
rect 17644 9092 17650 9104
rect 21450 9092 21456 9104
rect 17644 9064 21456 9092
rect 17644 9052 17650 9064
rect 21450 9052 21456 9064
rect 21508 9052 21514 9104
rect 18414 9024 18420 9036
rect 18375 8996 18420 9024
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 19392 8996 19441 9024
rect 19392 8984 19398 8996
rect 19429 8993 19441 8996
rect 19475 9024 19487 9027
rect 20070 9024 20076 9036
rect 19475 8996 20076 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 20441 9027 20499 9033
rect 20441 8993 20453 9027
rect 20487 9024 20499 9027
rect 21560 9024 21588 9132
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 24026 9120 24032 9172
rect 24084 9160 24090 9172
rect 25958 9160 25964 9172
rect 24084 9132 25964 9160
rect 24084 9120 24090 9132
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26329 9163 26387 9169
rect 26329 9129 26341 9163
rect 26375 9160 26387 9163
rect 27614 9160 27620 9172
rect 26375 9132 27620 9160
rect 26375 9129 26387 9132
rect 26329 9123 26387 9129
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 28166 9120 28172 9172
rect 28224 9160 28230 9172
rect 29362 9160 29368 9172
rect 28224 9132 29368 9160
rect 28224 9120 28230 9132
rect 29362 9120 29368 9132
rect 29420 9160 29426 9172
rect 32306 9160 32312 9172
rect 29420 9132 31754 9160
rect 32267 9132 32312 9160
rect 29420 9120 29426 9132
rect 22922 9052 22928 9104
rect 22980 9092 22986 9104
rect 23382 9092 23388 9104
rect 22980 9064 23388 9092
rect 22980 9052 22986 9064
rect 23382 9052 23388 9064
rect 23440 9052 23446 9104
rect 23750 9052 23756 9104
rect 23808 9092 23814 9104
rect 23808 9064 24716 9092
rect 23808 9052 23814 9064
rect 20487 8996 21588 9024
rect 20487 8993 20499 8996
rect 20441 8987 20499 8993
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22833 9027 22891 9033
rect 22833 9024 22845 9027
rect 22060 8996 22845 9024
rect 22060 8984 22066 8996
rect 22833 8993 22845 8996
rect 22879 9024 22891 9027
rect 24210 9024 24216 9036
rect 22879 8996 24216 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 24210 8984 24216 8996
rect 24268 9024 24274 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 24268 8996 24593 9024
rect 24268 8984 24274 8996
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24688 9024 24716 9064
rect 28258 9052 28264 9104
rect 28316 9092 28322 9104
rect 31386 9092 31392 9104
rect 28316 9064 31392 9092
rect 28316 9052 28322 9064
rect 31386 9052 31392 9064
rect 31444 9052 31450 9104
rect 31726 9092 31754 9132
rect 32306 9120 32312 9132
rect 32364 9120 32370 9172
rect 32858 9160 32864 9172
rect 32819 9132 32864 9160
rect 32858 9120 32864 9132
rect 32916 9120 32922 9172
rect 33134 9092 33140 9104
rect 31726 9064 33140 9092
rect 33134 9052 33140 9064
rect 33192 9052 33198 9104
rect 24857 9027 24915 9033
rect 24857 9024 24869 9027
rect 24688 8996 24869 9024
rect 24581 8987 24639 8993
rect 24857 8993 24869 8996
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 25222 8984 25228 9036
rect 25280 9024 25286 9036
rect 26789 9027 26847 9033
rect 25280 8996 26096 9024
rect 25280 8984 25286 8996
rect 1903 8928 2452 8956
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 17276 8928 17785 8956
rect 17276 8916 17282 8928
rect 17773 8925 17785 8928
rect 17819 8925 17831 8959
rect 17773 8919 17831 8925
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18012 8928 18245 8956
rect 18012 8916 18018 8928
rect 18233 8925 18245 8928
rect 18279 8956 18291 8959
rect 19242 8956 19248 8968
rect 18279 8928 19248 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 25958 8916 25964 8968
rect 26016 8916 26022 8968
rect 26068 8956 26096 8996
rect 26789 8993 26801 9027
rect 26835 9024 26847 9027
rect 29178 9024 29184 9036
rect 26835 8996 29184 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 29178 8984 29184 8996
rect 29236 8984 29242 9036
rect 33689 8959 33747 8965
rect 26068 8928 26188 8956
rect 17681 8891 17739 8897
rect 17681 8857 17693 8891
rect 17727 8888 17739 8891
rect 20349 8891 20407 8897
rect 17727 8860 19380 8888
rect 17727 8857 17739 8860
rect 17681 8851 17739 8857
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 19352 8820 19380 8860
rect 20349 8857 20361 8891
rect 20395 8857 20407 8891
rect 20349 8851 20407 8857
rect 20364 8820 20392 8851
rect 21818 8848 21824 8900
rect 21876 8848 21882 8900
rect 22462 8848 22468 8900
rect 22520 8888 22526 8900
rect 22557 8891 22615 8897
rect 22557 8888 22569 8891
rect 22520 8860 22569 8888
rect 22520 8848 22526 8860
rect 22557 8857 22569 8860
rect 22603 8857 22615 8891
rect 22557 8851 22615 8857
rect 23293 8891 23351 8897
rect 23293 8857 23305 8891
rect 23339 8857 23351 8891
rect 23842 8888 23848 8900
rect 23803 8860 23848 8888
rect 23293 8851 23351 8857
rect 19352 8792 20392 8820
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 20990 8820 20996 8832
rect 20864 8792 20996 8820
rect 20864 8780 20870 8792
rect 20990 8780 20996 8792
rect 21048 8820 21054 8832
rect 21085 8823 21143 8829
rect 21085 8820 21097 8823
rect 21048 8792 21097 8820
rect 21048 8780 21054 8792
rect 21085 8789 21097 8792
rect 21131 8789 21143 8823
rect 21085 8783 21143 8789
rect 21726 8780 21732 8832
rect 21784 8820 21790 8832
rect 23308 8820 23336 8851
rect 23842 8848 23848 8860
rect 23900 8848 23906 8900
rect 23937 8891 23995 8897
rect 23937 8857 23949 8891
rect 23983 8888 23995 8891
rect 24118 8888 24124 8900
rect 23983 8860 24124 8888
rect 23983 8857 23995 8860
rect 23937 8851 23995 8857
rect 24118 8848 24124 8860
rect 24176 8848 24182 8900
rect 25130 8888 25136 8900
rect 24780 8860 25136 8888
rect 21784 8792 23336 8820
rect 21784 8780 21790 8792
rect 23382 8780 23388 8832
rect 23440 8820 23446 8832
rect 24780 8820 24808 8860
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 26160 8888 26188 8928
rect 33689 8925 33701 8959
rect 33735 8956 33747 8959
rect 34241 8959 34299 8965
rect 34241 8956 34253 8959
rect 33735 8928 34253 8956
rect 33735 8925 33747 8928
rect 33689 8919 33747 8925
rect 34241 8925 34253 8928
rect 34287 8956 34299 8959
rect 34514 8956 34520 8968
rect 34287 8928 34520 8956
rect 34287 8925 34299 8928
rect 34241 8919 34299 8925
rect 34514 8916 34520 8928
rect 34572 8916 34578 8968
rect 27065 8891 27123 8897
rect 27065 8888 27077 8891
rect 26160 8860 27077 8888
rect 27065 8857 27077 8860
rect 27111 8888 27123 8891
rect 30466 8888 30472 8900
rect 27111 8860 27476 8888
rect 28290 8860 30472 8888
rect 27111 8857 27123 8860
rect 27065 8851 27123 8857
rect 23440 8792 24808 8820
rect 27448 8820 27476 8860
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 35894 8848 35900 8900
rect 35952 8888 35958 8900
rect 35952 8860 35997 8888
rect 35952 8848 35958 8860
rect 28442 8820 28448 8832
rect 27448 8792 28448 8820
rect 23440 8780 23446 8792
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 28537 8823 28595 8829
rect 28537 8789 28549 8823
rect 28583 8820 28595 8823
rect 28626 8820 28632 8832
rect 28583 8792 28632 8820
rect 28583 8789 28595 8792
rect 28537 8783 28595 8789
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 29089 8823 29147 8829
rect 29089 8789 29101 8823
rect 29135 8820 29147 8823
rect 29178 8820 29184 8832
rect 29135 8792 29184 8820
rect 29135 8789 29147 8792
rect 29089 8783 29147 8789
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 34238 8780 34244 8832
rect 34296 8820 34302 8832
rect 34885 8823 34943 8829
rect 34885 8820 34897 8823
rect 34296 8792 34897 8820
rect 34296 8780 34302 8792
rect 34885 8789 34897 8792
rect 34931 8789 34943 8823
rect 34885 8783 34943 8789
rect 1104 8730 36892 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 36892 8730
rect 1104 8656 36892 8678
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 19518 8616 19524 8628
rect 17828 8588 19524 8616
rect 17828 8576 17834 8588
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 20898 8616 20904 8628
rect 19628 8588 20904 8616
rect 17865 8551 17923 8557
rect 17865 8517 17877 8551
rect 17911 8548 17923 8551
rect 18601 8551 18659 8557
rect 18601 8548 18613 8551
rect 17911 8520 18613 8548
rect 17911 8517 17923 8520
rect 17865 8511 17923 8517
rect 18601 8517 18613 8520
rect 18647 8517 18659 8551
rect 18601 8511 18659 8517
rect 17770 8480 17776 8492
rect 17731 8452 17776 8480
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 19628 8489 19656 8588
rect 20898 8576 20904 8588
rect 20956 8616 20962 8628
rect 20956 8588 21220 8616
rect 20956 8576 20962 8588
rect 19886 8548 19892 8560
rect 19847 8520 19892 8548
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 20990 8440 20996 8492
rect 21048 8440 21054 8492
rect 21192 8480 21220 8588
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 36078 8616 36084 8628
rect 21600 8588 36084 8616
rect 21600 8576 21606 8588
rect 36078 8576 36084 8588
rect 36136 8576 36142 8628
rect 23290 8548 23296 8560
rect 23138 8520 23296 8548
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 28258 8548 28264 8560
rect 25806 8520 28264 8548
rect 28258 8508 28264 8520
rect 28316 8508 28322 8560
rect 31570 8548 31576 8560
rect 29210 8520 31576 8548
rect 31570 8508 31576 8520
rect 31628 8508 31634 8560
rect 31757 8551 31815 8557
rect 31757 8517 31769 8551
rect 31803 8548 31815 8551
rect 31846 8548 31852 8560
rect 31803 8520 31852 8548
rect 31803 8517 31815 8520
rect 31757 8511 31815 8517
rect 31846 8508 31852 8520
rect 31904 8548 31910 8560
rect 32306 8548 32312 8560
rect 31904 8520 32312 8548
rect 31904 8508 31910 8520
rect 32306 8508 32312 8520
rect 32364 8548 32370 8560
rect 32493 8551 32551 8557
rect 32493 8548 32505 8551
rect 32364 8520 32505 8548
rect 32364 8508 32370 8520
rect 32493 8517 32505 8520
rect 32539 8517 32551 8551
rect 32493 8511 32551 8517
rect 22094 8480 22100 8492
rect 21192 8452 22100 8480
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8480 23903 8483
rect 24210 8480 24216 8492
rect 23891 8452 24216 8480
rect 23891 8449 23903 8452
rect 23845 8443 23903 8449
rect 24210 8440 24216 8452
rect 24268 8480 24274 8492
rect 24305 8483 24363 8489
rect 24305 8480 24317 8483
rect 24268 8452 24317 8480
rect 24268 8440 24274 8452
rect 24305 8449 24317 8452
rect 24351 8449 24363 8483
rect 24305 8443 24363 8449
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8480 27399 8483
rect 28166 8480 28172 8492
rect 27387 8452 28172 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 28166 8440 28172 8452
rect 28224 8440 28230 8492
rect 33229 8483 33287 8489
rect 33229 8449 33241 8483
rect 33275 8480 33287 8483
rect 33275 8452 33824 8480
rect 33275 8449 33287 8452
rect 33229 8443 33287 8449
rect 18506 8412 18512 8424
rect 18467 8384 18512 8412
rect 18506 8372 18512 8384
rect 18564 8412 18570 8424
rect 19334 8412 19340 8424
rect 18564 8384 19340 8412
rect 18564 8372 18570 8384
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 24578 8412 24584 8424
rect 24539 8384 24584 8412
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 27249 8415 27307 8421
rect 27249 8412 27261 8415
rect 24728 8384 27261 8412
rect 24728 8372 24734 8384
rect 27249 8381 27261 8384
rect 27295 8381 27307 8415
rect 27522 8412 27528 8424
rect 27249 8375 27307 8381
rect 27356 8384 27528 8412
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8313 19119 8347
rect 21726 8344 21732 8356
rect 19061 8307 19119 8313
rect 20916 8316 21732 8344
rect 19076 8276 19104 8307
rect 19426 8276 19432 8288
rect 19076 8248 19432 8276
rect 19426 8236 19432 8248
rect 19484 8276 19490 8288
rect 20916 8276 20944 8316
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 22094 8304 22100 8356
rect 22152 8344 22158 8356
rect 27356 8344 27384 8384
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 27893 8415 27951 8421
rect 27893 8412 27905 8415
rect 27580 8384 27905 8412
rect 27580 8372 27586 8384
rect 27893 8381 27905 8384
rect 27939 8381 27951 8415
rect 29641 8415 29699 8421
rect 29641 8412 29653 8415
rect 27893 8375 27951 8381
rect 28368 8384 29653 8412
rect 22152 8316 22197 8344
rect 25884 8316 27384 8344
rect 22152 8304 22158 8316
rect 19484 8248 20944 8276
rect 19484 8236 19490 8248
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 21361 8279 21419 8285
rect 21361 8276 21373 8279
rect 21232 8248 21373 8276
rect 21232 8236 21238 8248
rect 21361 8245 21373 8248
rect 21407 8245 21419 8279
rect 21361 8239 21419 8245
rect 21450 8236 21456 8288
rect 21508 8276 21514 8288
rect 23581 8279 23639 8285
rect 23581 8276 23593 8279
rect 21508 8248 23593 8276
rect 21508 8236 21514 8248
rect 23581 8245 23593 8248
rect 23627 8276 23639 8279
rect 25884 8276 25912 8316
rect 27430 8304 27436 8356
rect 27488 8344 27494 8356
rect 28368 8344 28396 8384
rect 29641 8381 29653 8384
rect 29687 8381 29699 8415
rect 29641 8375 29699 8381
rect 29917 8415 29975 8421
rect 29917 8381 29929 8415
rect 29963 8381 29975 8415
rect 29917 8375 29975 8381
rect 27488 8316 28396 8344
rect 29932 8344 29960 8375
rect 30282 8344 30288 8356
rect 29932 8316 30288 8344
rect 27488 8304 27494 8316
rect 30282 8304 30288 8316
rect 30340 8344 30346 8356
rect 30377 8347 30435 8353
rect 30377 8344 30389 8347
rect 30340 8316 30389 8344
rect 30340 8304 30346 8316
rect 30377 8313 30389 8316
rect 30423 8313 30435 8347
rect 30377 8307 30435 8313
rect 31754 8304 31760 8356
rect 31812 8344 31818 8356
rect 33796 8353 33824 8452
rect 33137 8347 33195 8353
rect 33137 8344 33149 8347
rect 31812 8316 33149 8344
rect 31812 8304 31818 8316
rect 33137 8313 33149 8316
rect 33183 8313 33195 8347
rect 33137 8307 33195 8313
rect 33781 8347 33839 8353
rect 33781 8313 33793 8347
rect 33827 8344 33839 8347
rect 34514 8344 34520 8356
rect 33827 8316 34520 8344
rect 33827 8313 33839 8316
rect 33781 8307 33839 8313
rect 34514 8304 34520 8316
rect 34572 8344 34578 8356
rect 34977 8347 35035 8353
rect 34977 8344 34989 8347
rect 34572 8316 34989 8344
rect 34572 8304 34578 8316
rect 34977 8313 34989 8316
rect 35023 8344 35035 8347
rect 35342 8344 35348 8356
rect 35023 8316 35348 8344
rect 35023 8313 35035 8316
rect 34977 8307 35035 8313
rect 35342 8304 35348 8316
rect 35400 8304 35406 8356
rect 36262 8344 36268 8356
rect 36223 8316 36268 8344
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 26050 8276 26056 8288
rect 23627 8248 25912 8276
rect 26011 8248 26056 8276
rect 23627 8245 23639 8248
rect 23581 8239 23639 8245
rect 26050 8236 26056 8248
rect 26108 8236 26114 8288
rect 34146 8236 34152 8288
rect 34204 8276 34210 8288
rect 34241 8279 34299 8285
rect 34241 8276 34253 8279
rect 34204 8248 34253 8276
rect 34204 8236 34210 8248
rect 34241 8245 34253 8248
rect 34287 8245 34299 8279
rect 35434 8276 35440 8288
rect 35395 8248 35440 8276
rect 34241 8239 34299 8245
rect 35434 8236 35440 8248
rect 35492 8236 35498 8288
rect 1104 8186 36892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36892 8186
rect 1104 8112 36892 8134
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 23293 8075 23351 8081
rect 23293 8072 23305 8075
rect 22244 8044 23305 8072
rect 22244 8032 22250 8044
rect 23293 8041 23305 8044
rect 23339 8041 23351 8075
rect 23934 8072 23940 8084
rect 23895 8044 23940 8072
rect 23293 8035 23351 8041
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 24486 8032 24492 8084
rect 24544 8072 24550 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 24544 8044 24685 8072
rect 24544 8032 24550 8044
rect 24673 8041 24685 8044
rect 24719 8041 24731 8075
rect 24673 8035 24731 8041
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 26586 8075 26644 8081
rect 26586 8072 26598 8075
rect 26108 8044 26598 8072
rect 26108 8032 26114 8044
rect 26586 8041 26598 8044
rect 26632 8072 26644 8075
rect 29086 8072 29092 8084
rect 26632 8044 29092 8072
rect 26632 8041 26644 8044
rect 26586 8035 26644 8041
rect 29086 8032 29092 8044
rect 29144 8032 29150 8084
rect 31202 8032 31208 8084
rect 31260 8072 31266 8084
rect 31757 8075 31815 8081
rect 31757 8072 31769 8075
rect 31260 8044 31769 8072
rect 31260 8032 31266 8044
rect 31757 8041 31769 8044
rect 31803 8072 31815 8075
rect 31846 8072 31852 8084
rect 31803 8044 31852 8072
rect 31803 8041 31815 8044
rect 31757 8035 31815 8041
rect 31846 8032 31852 8044
rect 31904 8032 31910 8084
rect 22649 8007 22707 8013
rect 20088 7976 21036 8004
rect 20088 7945 20116 7976
rect 20073 7939 20131 7945
rect 18708 7908 20024 7936
rect 18708 7877 18736 7908
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 19889 7871 19947 7877
rect 19889 7868 19901 7871
rect 18831 7840 19901 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 19889 7837 19901 7840
rect 19935 7837 19947 7871
rect 19996 7868 20024 7908
rect 20073 7905 20085 7939
rect 20119 7905 20131 7939
rect 20898 7936 20904 7948
rect 20859 7908 20904 7936
rect 20073 7899 20131 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 21008 7936 21036 7976
rect 22649 7973 22661 8007
rect 22695 8004 22707 8007
rect 23014 8004 23020 8016
rect 22695 7976 23020 8004
rect 22695 7973 22707 7976
rect 22649 7967 22707 7973
rect 23014 7964 23020 7976
rect 23072 7964 23078 8016
rect 28077 8007 28135 8013
rect 28077 7973 28089 8007
rect 28123 8004 28135 8007
rect 28718 8004 28724 8016
rect 28123 7976 28724 8004
rect 28123 7973 28135 7976
rect 28077 7967 28135 7973
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 33410 7964 33416 8016
rect 33468 8004 33474 8016
rect 33468 7976 35894 8004
rect 33468 7964 33474 7976
rect 24118 7936 24124 7948
rect 21008 7908 24124 7936
rect 24118 7896 24124 7908
rect 24176 7936 24182 7948
rect 24670 7936 24676 7948
rect 24176 7908 24676 7936
rect 24176 7896 24182 7908
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7936 25375 7939
rect 25869 7939 25927 7945
rect 25869 7936 25881 7939
rect 25363 7908 25881 7936
rect 25363 7905 25375 7908
rect 25317 7899 25375 7905
rect 25869 7905 25881 7908
rect 25915 7936 25927 7939
rect 26142 7936 26148 7948
rect 25915 7908 26148 7936
rect 25915 7905 25927 7908
rect 25869 7899 25927 7905
rect 26142 7896 26148 7908
rect 26200 7936 26206 7948
rect 26329 7939 26387 7945
rect 26329 7936 26341 7939
rect 26200 7908 26341 7936
rect 26200 7896 26206 7908
rect 26329 7905 26341 7908
rect 26375 7936 26387 7939
rect 29178 7936 29184 7948
rect 26375 7908 29184 7936
rect 26375 7905 26387 7908
rect 26329 7899 26387 7905
rect 29178 7896 29184 7908
rect 29236 7896 29242 7948
rect 32858 7896 32864 7948
rect 32916 7936 32922 7948
rect 33597 7939 33655 7945
rect 33597 7936 33609 7939
rect 32916 7908 33609 7936
rect 32916 7896 32922 7908
rect 20806 7868 20812 7880
rect 19996 7840 20812 7868
rect 19889 7831 19947 7837
rect 17589 7803 17647 7809
rect 17589 7769 17601 7803
rect 17635 7800 17647 7803
rect 18064 7800 18092 7831
rect 20806 7828 20812 7840
rect 20864 7828 20870 7880
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 23658 7868 23664 7880
rect 23431 7840 23664 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 24026 7868 24032 7880
rect 23987 7840 24032 7868
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 24762 7868 24768 7880
rect 24723 7840 24768 7868
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 29638 7868 29644 7880
rect 27738 7840 29644 7868
rect 29638 7828 29644 7840
rect 29696 7828 29702 7880
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 33152 7877 33180 7908
rect 33597 7905 33609 7908
rect 33643 7936 33655 7939
rect 34514 7936 34520 7948
rect 33643 7908 34520 7936
rect 33643 7905 33655 7908
rect 33597 7899 33655 7905
rect 34514 7896 34520 7908
rect 34572 7936 34578 7948
rect 34885 7939 34943 7945
rect 34885 7936 34897 7939
rect 34572 7908 34897 7936
rect 34572 7896 34578 7908
rect 34885 7905 34897 7908
rect 34931 7936 34943 7939
rect 35434 7936 35440 7948
rect 34931 7908 35440 7936
rect 34931 7905 34943 7908
rect 34885 7899 34943 7905
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 35866 7936 35894 7976
rect 36081 7939 36139 7945
rect 36081 7936 36093 7939
rect 35866 7908 36093 7936
rect 36081 7905 36093 7908
rect 36127 7905 36139 7939
rect 36081 7899 36139 7905
rect 33045 7871 33103 7877
rect 33045 7868 33057 7871
rect 29972 7840 33057 7868
rect 29972 7828 29978 7840
rect 33045 7837 33057 7840
rect 33091 7837 33103 7871
rect 33045 7831 33103 7837
rect 33137 7871 33195 7877
rect 33137 7837 33149 7871
rect 33183 7837 33195 7871
rect 36354 7868 36360 7880
rect 36315 7840 36360 7868
rect 33137 7831 33195 7837
rect 36354 7828 36360 7840
rect 36412 7828 36418 7880
rect 21174 7800 21180 7812
rect 17635 7772 19564 7800
rect 21135 7772 21180 7800
rect 17635 7769 17647 7772
rect 17589 7763 17647 7769
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 19058 7732 19064 7744
rect 18187 7704 19064 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 19242 7692 19248 7744
rect 19300 7732 19306 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19300 7704 19441 7732
rect 19300 7692 19306 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19536 7732 19564 7772
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 31205 7803 31263 7809
rect 22402 7772 26556 7800
rect 22738 7732 22744 7744
rect 19536 7704 22744 7732
rect 19429 7695 19487 7701
rect 22738 7692 22744 7704
rect 22796 7692 22802 7744
rect 22830 7692 22836 7744
rect 22888 7732 22894 7744
rect 24026 7732 24032 7744
rect 22888 7704 24032 7732
rect 22888 7692 22894 7704
rect 24026 7692 24032 7704
rect 24084 7692 24090 7744
rect 26528 7732 26556 7772
rect 28000 7772 30420 7800
rect 28000 7732 28028 7772
rect 26528 7704 28028 7732
rect 28721 7735 28779 7741
rect 28721 7701 28733 7735
rect 28767 7732 28779 7735
rect 29178 7732 29184 7744
rect 28767 7704 29184 7732
rect 28767 7701 28779 7704
rect 28721 7695 28779 7701
rect 29178 7692 29184 7704
rect 29236 7732 29242 7744
rect 29733 7735 29791 7741
rect 29733 7732 29745 7735
rect 29236 7704 29745 7732
rect 29236 7692 29242 7704
rect 29733 7701 29745 7704
rect 29779 7732 29791 7735
rect 30282 7732 30288 7744
rect 29779 7704 30288 7732
rect 29779 7701 29791 7704
rect 29733 7695 29791 7701
rect 30282 7692 30288 7704
rect 30340 7692 30346 7744
rect 30392 7732 30420 7772
rect 31205 7769 31217 7803
rect 31251 7800 31263 7803
rect 32122 7800 32128 7812
rect 31251 7772 32128 7800
rect 31251 7769 31263 7772
rect 31205 7763 31263 7769
rect 32122 7760 32128 7772
rect 32180 7760 32186 7812
rect 32030 7732 32036 7744
rect 30392 7704 32036 7732
rect 32030 7692 32036 7704
rect 32088 7692 32094 7744
rect 32306 7732 32312 7744
rect 32267 7704 32312 7732
rect 32306 7692 32312 7704
rect 32364 7692 32370 7744
rect 34146 7732 34152 7744
rect 34107 7704 34152 7732
rect 34146 7692 34152 7704
rect 34204 7692 34210 7744
rect 1104 7642 36892 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 36892 7642
rect 1104 7568 36892 7590
rect 20530 7528 20536 7540
rect 17328 7500 20536 7528
rect 17328 7469 17356 7500
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 22097 7531 22155 7537
rect 22097 7497 22109 7531
rect 22143 7528 22155 7531
rect 22186 7528 22192 7540
rect 22143 7500 22192 7528
rect 22143 7497 22155 7500
rect 22097 7491 22155 7497
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 22741 7531 22799 7537
rect 22741 7497 22753 7531
rect 22787 7528 22799 7531
rect 23842 7528 23848 7540
rect 22787 7500 23848 7528
rect 22787 7497 22799 7500
rect 22741 7491 22799 7497
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 25777 7531 25835 7537
rect 25777 7497 25789 7531
rect 25823 7497 25835 7531
rect 25777 7491 25835 7497
rect 17313 7463 17371 7469
rect 17313 7429 17325 7463
rect 17359 7429 17371 7463
rect 18230 7460 18236 7472
rect 18191 7432 18236 7460
rect 17313 7423 17371 7429
rect 18230 7420 18236 7432
rect 18288 7420 18294 7472
rect 19058 7460 19064 7472
rect 19019 7432 19064 7460
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 19334 7420 19340 7472
rect 19392 7460 19398 7472
rect 23750 7460 23756 7472
rect 19392 7432 20484 7460
rect 19392 7420 19398 7432
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 20456 7401 20484 7432
rect 22204 7432 23756 7460
rect 22204 7401 22232 7432
rect 23750 7420 23756 7432
rect 23808 7420 23814 7472
rect 24302 7460 24308 7472
rect 24044 7432 24308 7460
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7392 22707 7395
rect 23014 7392 23020 7404
rect 22695 7364 23020 7392
rect 22695 7361 22707 7364
rect 22649 7355 22707 7361
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 24044 7392 24072 7432
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 25792 7460 25820 7491
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 26421 7531 26479 7537
rect 26421 7528 26433 7531
rect 26200 7500 26433 7528
rect 26200 7488 26206 7500
rect 26421 7497 26433 7500
rect 26467 7497 26479 7531
rect 26421 7491 26479 7497
rect 28902 7488 28908 7540
rect 28960 7528 28966 7540
rect 29733 7531 29791 7537
rect 29733 7528 29745 7531
rect 28960 7500 29745 7528
rect 28960 7488 28966 7500
rect 29733 7497 29745 7500
rect 29779 7528 29791 7531
rect 36354 7528 36360 7540
rect 29779 7500 35894 7528
rect 36315 7500 36360 7528
rect 29779 7497 29791 7500
rect 29733 7491 29791 7497
rect 26510 7460 26516 7472
rect 25792 7432 26516 7460
rect 26510 7420 26516 7432
rect 26568 7420 26574 7472
rect 27157 7463 27215 7469
rect 27157 7429 27169 7463
rect 27203 7460 27215 7463
rect 27246 7460 27252 7472
rect 27203 7432 27252 7460
rect 27203 7429 27215 7432
rect 27157 7423 27215 7429
rect 27246 7420 27252 7432
rect 27304 7420 27310 7472
rect 31754 7460 31760 7472
rect 28474 7432 31760 7460
rect 31754 7420 31760 7432
rect 31812 7420 31818 7472
rect 33781 7463 33839 7469
rect 33781 7460 33793 7463
rect 31864 7432 33793 7460
rect 23523 7364 24072 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 25406 7352 25412 7404
rect 25464 7352 25470 7404
rect 25958 7352 25964 7404
rect 26016 7392 26022 7404
rect 27338 7392 27344 7404
rect 26016 7364 27344 7392
rect 26016 7352 26022 7364
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 30653 7395 30711 7401
rect 30653 7361 30665 7395
rect 30699 7392 30711 7395
rect 31202 7392 31208 7404
rect 30699 7364 31208 7392
rect 30699 7361 30711 7364
rect 30653 7355 30711 7361
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 31864 7392 31892 7432
rect 33781 7429 33793 7432
rect 33827 7429 33839 7463
rect 33781 7423 33839 7429
rect 34698 7420 34704 7472
rect 34756 7460 34762 7472
rect 35342 7460 35348 7472
rect 34756 7432 35348 7460
rect 34756 7420 34762 7432
rect 35342 7420 35348 7432
rect 35400 7460 35406 7472
rect 35437 7463 35495 7469
rect 35437 7460 35449 7463
rect 35400 7432 35449 7460
rect 35400 7420 35406 7432
rect 35437 7429 35449 7432
rect 35483 7429 35495 7463
rect 35866 7460 35894 7500
rect 36354 7488 36360 7500
rect 36412 7488 36418 7540
rect 36446 7460 36452 7472
rect 35866 7432 36452 7460
rect 35437 7423 35495 7429
rect 36446 7420 36452 7432
rect 36504 7420 36510 7472
rect 31726 7364 31892 7392
rect 18325 7327 18383 7333
rect 18325 7293 18337 7327
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7324 19027 7327
rect 19426 7324 19432 7336
rect 19015 7296 19432 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 18340 7256 18368 7287
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7324 20039 7327
rect 20254 7324 20260 7336
rect 20027 7296 20260 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20622 7324 20628 7336
rect 20583 7296 20628 7324
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 23385 7327 23443 7333
rect 23385 7324 23397 7327
rect 20772 7296 23397 7324
rect 20772 7284 20778 7296
rect 23385 7293 23397 7296
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 24026 7284 24032 7336
rect 24084 7324 24090 7336
rect 24302 7324 24308 7336
rect 24084 7296 24129 7324
rect 24215 7296 24308 7324
rect 24084 7284 24090 7296
rect 24302 7284 24308 7296
rect 24360 7324 24366 7336
rect 27890 7324 27896 7336
rect 24360 7296 27896 7324
rect 24360 7284 24366 7296
rect 27890 7284 27896 7296
rect 27948 7284 27954 7336
rect 28902 7324 28908 7336
rect 28863 7296 28908 7324
rect 28902 7284 28908 7296
rect 28960 7284 28966 7336
rect 29178 7324 29184 7336
rect 29139 7296 29184 7324
rect 29178 7284 29184 7296
rect 29236 7284 29242 7336
rect 31726 7324 31754 7364
rect 32306 7352 32312 7404
rect 32364 7392 32370 7404
rect 32585 7395 32643 7401
rect 32585 7392 32597 7395
rect 32364 7364 32597 7392
rect 32364 7352 32370 7364
rect 32585 7361 32597 7364
rect 32631 7361 32643 7395
rect 32585 7355 32643 7361
rect 30852 7296 31754 7324
rect 18598 7256 18604 7268
rect 18340 7228 18604 7256
rect 18598 7216 18604 7228
rect 18656 7256 18662 7268
rect 19242 7256 19248 7268
rect 18656 7228 19248 7256
rect 18656 7216 18662 7228
rect 19242 7216 19248 7228
rect 19300 7256 19306 7268
rect 20809 7259 20867 7265
rect 20809 7256 20821 7259
rect 19300 7228 20821 7256
rect 19300 7216 19306 7228
rect 20809 7225 20821 7228
rect 20855 7225 20867 7259
rect 20809 7219 20867 7225
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 21174 7188 21180 7200
rect 19392 7160 21180 7188
rect 19392 7148 19398 7160
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 22738 7148 22744 7200
rect 22796 7188 22802 7200
rect 25498 7188 25504 7200
rect 22796 7160 25504 7188
rect 22796 7148 22802 7160
rect 25498 7148 25504 7160
rect 25556 7148 25562 7200
rect 28442 7148 28448 7200
rect 28500 7188 28506 7200
rect 30852 7188 30880 7296
rect 30926 7216 30932 7268
rect 30984 7256 30990 7268
rect 32493 7259 32551 7265
rect 32493 7256 32505 7259
rect 30984 7228 32505 7256
rect 30984 7216 30990 7228
rect 32493 7225 32505 7228
rect 32539 7225 32551 7259
rect 32600 7256 32628 7355
rect 32766 7352 32772 7404
rect 32824 7392 32830 7404
rect 33229 7395 33287 7401
rect 33229 7392 33241 7395
rect 32824 7364 33241 7392
rect 32824 7352 32830 7364
rect 33229 7361 33241 7364
rect 33275 7392 33287 7395
rect 33873 7395 33931 7401
rect 33873 7392 33885 7395
rect 33275 7364 33885 7392
rect 33275 7361 33287 7364
rect 33229 7355 33287 7361
rect 33873 7361 33885 7364
rect 33919 7392 33931 7395
rect 34146 7392 34152 7404
rect 33919 7364 34152 7392
rect 33919 7361 33931 7364
rect 33873 7355 33931 7361
rect 34146 7352 34152 7364
rect 34204 7392 34210 7404
rect 34333 7395 34391 7401
rect 34333 7392 34345 7395
rect 34204 7364 34345 7392
rect 34204 7352 34210 7364
rect 34333 7361 34345 7364
rect 34379 7392 34391 7395
rect 34885 7395 34943 7401
rect 34885 7392 34897 7395
rect 34379 7364 34897 7392
rect 34379 7361 34391 7364
rect 34333 7355 34391 7361
rect 34885 7361 34897 7364
rect 34931 7392 34943 7395
rect 35526 7392 35532 7404
rect 34931 7364 35532 7392
rect 34931 7361 34943 7364
rect 34885 7355 34943 7361
rect 35526 7352 35532 7364
rect 35584 7352 35590 7404
rect 34698 7256 34704 7268
rect 32600 7228 34704 7256
rect 32493 7219 32551 7225
rect 34698 7216 34704 7228
rect 34756 7216 34762 7268
rect 28500 7160 30880 7188
rect 31757 7191 31815 7197
rect 28500 7148 28506 7160
rect 31757 7157 31769 7191
rect 31803 7188 31815 7191
rect 31846 7188 31852 7200
rect 31803 7160 31852 7188
rect 31803 7157 31815 7160
rect 31757 7151 31815 7157
rect 31846 7148 31852 7160
rect 31904 7148 31910 7200
rect 31938 7148 31944 7200
rect 31996 7188 32002 7200
rect 33137 7191 33195 7197
rect 33137 7188 33149 7191
rect 31996 7160 33149 7188
rect 31996 7148 32002 7160
rect 33137 7157 33149 7160
rect 33183 7157 33195 7191
rect 33137 7151 33195 7157
rect 1104 7098 36892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36892 7098
rect 1104 7024 36892 7046
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19484 6956 20116 6984
rect 19484 6944 19490 6956
rect 20088 6925 20116 6956
rect 25406 6944 25412 6996
rect 25464 6984 25470 6996
rect 32950 6984 32956 6996
rect 25464 6956 32956 6984
rect 25464 6944 25470 6956
rect 32950 6944 32956 6956
rect 33008 6944 33014 6996
rect 35526 6984 35532 6996
rect 35487 6956 35532 6984
rect 35526 6944 35532 6956
rect 35584 6944 35590 6996
rect 20073 6919 20131 6925
rect 18708 6888 19012 6916
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 18230 6848 18236 6860
rect 17451 6820 18236 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 1946 6740 1952 6792
rect 2004 6780 2010 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 2004 6752 9137 6780
rect 2004 6740 2010 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 17494 6780 17500 6792
rect 17455 6752 17500 6780
rect 9125 6743 9183 6749
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17957 6783 18015 6789
rect 17957 6780 17969 6783
rect 17644 6752 17969 6780
rect 17644 6740 17650 6752
rect 17957 6749 17969 6752
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18708 6780 18736 6888
rect 18984 6848 19012 6888
rect 19306 6888 19472 6916
rect 19306 6848 19334 6888
rect 18984 6820 19334 6848
rect 19444 6848 19472 6888
rect 20073 6885 20085 6919
rect 20119 6885 20131 6919
rect 29362 6916 29368 6928
rect 20073 6879 20131 6885
rect 26988 6888 29368 6916
rect 20622 6848 20628 6860
rect 19444 6820 20628 6848
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 20806 6848 20812 6860
rect 20767 6820 20812 6848
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 21634 6808 21640 6860
rect 21692 6848 21698 6860
rect 22833 6851 22891 6857
rect 22833 6848 22845 6851
rect 21692 6820 22845 6848
rect 21692 6808 21698 6820
rect 22833 6817 22845 6820
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 23198 6808 23204 6860
rect 23256 6848 23262 6860
rect 23293 6851 23351 6857
rect 23293 6848 23305 6851
rect 23256 6820 23305 6848
rect 23256 6808 23262 6820
rect 23293 6817 23305 6820
rect 23339 6817 23351 6851
rect 23293 6811 23351 6817
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24026 6848 24032 6860
rect 23983 6820 24032 6848
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24026 6808 24032 6820
rect 24084 6848 24090 6860
rect 24673 6851 24731 6857
rect 24673 6848 24685 6851
rect 24084 6820 24685 6848
rect 24084 6808 24090 6820
rect 24673 6817 24685 6820
rect 24719 6848 24731 6851
rect 25225 6851 25283 6857
rect 25225 6848 25237 6851
rect 24719 6820 25237 6848
rect 24719 6817 24731 6820
rect 24673 6811 24731 6817
rect 25225 6817 25237 6820
rect 25271 6848 25283 6851
rect 25685 6851 25743 6857
rect 25685 6848 25697 6851
rect 25271 6820 25697 6848
rect 25271 6817 25283 6820
rect 25225 6811 25283 6817
rect 25685 6817 25697 6820
rect 25731 6848 25743 6851
rect 26050 6848 26056 6860
rect 25731 6820 26056 6848
rect 25731 6817 25743 6820
rect 25685 6811 25743 6817
rect 26050 6808 26056 6820
rect 26108 6808 26114 6860
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 26988 6848 27016 6888
rect 29362 6876 29368 6888
rect 29420 6916 29426 6928
rect 29546 6916 29552 6928
rect 29420 6888 29552 6916
rect 29420 6876 29426 6888
rect 29546 6876 29552 6888
rect 29604 6876 29610 6928
rect 26384 6820 27016 6848
rect 26384 6808 26390 6820
rect 27338 6808 27344 6860
rect 27396 6848 27402 6860
rect 32582 6848 32588 6860
rect 27396 6820 32588 6848
rect 27396 6808 27402 6820
rect 32582 6808 32588 6820
rect 32640 6808 32646 6860
rect 32858 6848 32864 6860
rect 32819 6820 32864 6848
rect 32858 6808 32864 6820
rect 32916 6808 32922 6860
rect 33042 6808 33048 6860
rect 33100 6848 33106 6860
rect 34149 6851 34207 6857
rect 34149 6848 34161 6851
rect 33100 6820 34161 6848
rect 33100 6808 33106 6820
rect 34149 6817 34161 6820
rect 34195 6817 34207 6851
rect 34149 6811 34207 6817
rect 34514 6808 34520 6860
rect 34572 6848 34578 6860
rect 34572 6820 35112 6848
rect 34572 6808 34578 6820
rect 35084 6792 35112 6820
rect 18095 6752 18736 6780
rect 18785 6783 18843 6789
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 18785 6749 18797 6783
rect 18831 6782 18843 6783
rect 18831 6780 18920 6782
rect 19334 6780 19340 6792
rect 18831 6754 19340 6780
rect 18831 6749 18843 6754
rect 18892 6752 19340 6754
rect 18785 6743 18843 6749
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 31481 6783 31539 6789
rect 28966 6752 29132 6780
rect 18966 6672 18972 6724
rect 19024 6712 19030 6724
rect 19521 6715 19579 6721
rect 19521 6712 19533 6715
rect 19024 6684 19533 6712
rect 19024 6672 19030 6684
rect 19521 6681 19533 6684
rect 19567 6681 19579 6715
rect 19521 6675 19579 6681
rect 19613 6715 19671 6721
rect 19613 6681 19625 6715
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 21085 6715 21143 6721
rect 21085 6681 21097 6715
rect 21131 6712 21143 6715
rect 21174 6712 21180 6724
rect 21131 6684 21180 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 18506 6644 18512 6656
rect 9263 6616 18512 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 18693 6647 18751 6653
rect 18693 6613 18705 6647
rect 18739 6644 18751 6647
rect 19628 6644 19656 6675
rect 21174 6672 21180 6684
rect 21232 6712 21238 6724
rect 21358 6712 21364 6724
rect 21232 6684 21364 6712
rect 21232 6672 21238 6684
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 25682 6712 25688 6724
rect 22310 6684 25688 6712
rect 25682 6672 25688 6684
rect 25740 6672 25746 6724
rect 25961 6715 26019 6721
rect 25961 6681 25973 6715
rect 26007 6712 26019 6715
rect 26234 6712 26240 6724
rect 26007 6684 26240 6712
rect 26007 6681 26019 6684
rect 25961 6675 26019 6681
rect 26234 6672 26240 6684
rect 26292 6672 26298 6724
rect 28966 6712 28994 6752
rect 27186 6684 28994 6712
rect 29104 6712 29132 6752
rect 31481 6749 31493 6783
rect 31527 6780 31539 6783
rect 31846 6780 31852 6792
rect 31527 6752 31852 6780
rect 31527 6749 31539 6752
rect 31481 6743 31539 6749
rect 31846 6740 31852 6752
rect 31904 6780 31910 6792
rect 32309 6783 32367 6789
rect 32309 6780 32321 6783
rect 31904 6752 32321 6780
rect 31904 6740 31910 6752
rect 32309 6749 32321 6752
rect 32355 6780 32367 6783
rect 32766 6780 32772 6792
rect 32355 6752 32772 6780
rect 32355 6749 32367 6752
rect 32309 6743 32367 6749
rect 32766 6740 32772 6752
rect 32824 6740 32830 6792
rect 32953 6783 33011 6789
rect 32953 6749 32965 6783
rect 32999 6780 33011 6783
rect 33226 6780 33232 6792
rect 32999 6752 33232 6780
rect 32999 6749 33011 6752
rect 32953 6743 33011 6749
rect 33226 6740 33232 6752
rect 33284 6740 33290 6792
rect 33597 6783 33655 6789
rect 33597 6749 33609 6783
rect 33643 6780 33655 6783
rect 33686 6780 33692 6792
rect 33643 6752 33692 6780
rect 33643 6749 33655 6752
rect 33597 6743 33655 6749
rect 33686 6740 33692 6752
rect 33744 6740 33750 6792
rect 34241 6783 34299 6789
rect 34241 6749 34253 6783
rect 34287 6780 34299 6783
rect 34698 6780 34704 6792
rect 34287 6752 34704 6780
rect 34287 6749 34299 6752
rect 34241 6743 34299 6749
rect 34698 6740 34704 6752
rect 34756 6740 34762 6792
rect 35066 6780 35072 6792
rect 35027 6752 35072 6780
rect 35066 6740 35072 6752
rect 35124 6780 35130 6792
rect 36081 6783 36139 6789
rect 36081 6780 36093 6783
rect 35124 6752 36093 6780
rect 35124 6740 35130 6752
rect 36081 6749 36093 6752
rect 36127 6749 36139 6783
rect 36081 6743 36139 6749
rect 34514 6712 34520 6724
rect 29104 6684 34520 6712
rect 34514 6672 34520 6684
rect 34572 6672 34578 6724
rect 18739 6616 19656 6644
rect 18739 6613 18751 6616
rect 18693 6607 18751 6613
rect 20254 6604 20260 6656
rect 20312 6644 20318 6656
rect 23014 6644 23020 6656
rect 20312 6616 23020 6644
rect 20312 6604 20318 6616
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 24394 6604 24400 6656
rect 24452 6644 24458 6656
rect 24762 6644 24768 6656
rect 24452 6616 24768 6644
rect 24452 6604 24458 6616
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25774 6644 25780 6656
rect 25004 6616 25780 6644
rect 25004 6604 25010 6616
rect 25774 6604 25780 6616
rect 25832 6604 25838 6656
rect 27433 6647 27491 6653
rect 27433 6613 27445 6647
rect 27479 6644 27491 6647
rect 27982 6644 27988 6656
rect 27479 6616 27988 6644
rect 27479 6613 27491 6616
rect 27433 6607 27491 6613
rect 27982 6604 27988 6616
rect 28040 6604 28046 6656
rect 28074 6604 28080 6656
rect 28132 6644 28138 6656
rect 28629 6647 28687 6653
rect 28629 6644 28641 6647
rect 28132 6616 28641 6644
rect 28132 6604 28138 6616
rect 28629 6613 28641 6616
rect 28675 6644 28687 6647
rect 29178 6644 29184 6656
rect 28675 6616 29184 6644
rect 28675 6613 28687 6616
rect 28629 6607 28687 6613
rect 29178 6604 29184 6616
rect 29236 6644 29242 6656
rect 29546 6644 29552 6656
rect 29236 6616 29552 6644
rect 29236 6604 29242 6616
rect 29546 6604 29552 6616
rect 29604 6644 29610 6656
rect 29733 6647 29791 6653
rect 29733 6644 29745 6647
rect 29604 6616 29745 6644
rect 29604 6604 29610 6616
rect 29733 6613 29745 6616
rect 29779 6613 29791 6647
rect 30742 6644 30748 6656
rect 30703 6616 30748 6644
rect 29733 6607 29791 6613
rect 30742 6604 30748 6616
rect 30800 6604 30806 6656
rect 31110 6604 31116 6656
rect 31168 6644 31174 6656
rect 32217 6647 32275 6653
rect 32217 6644 32229 6647
rect 31168 6616 32229 6644
rect 31168 6604 31174 6616
rect 32217 6613 32229 6616
rect 32263 6613 32275 6647
rect 32217 6607 32275 6613
rect 32398 6604 32404 6656
rect 32456 6644 32462 6656
rect 33226 6644 33232 6656
rect 32456 6616 33232 6644
rect 32456 6604 32462 6616
rect 33226 6604 33232 6616
rect 33284 6604 33290 6656
rect 33502 6644 33508 6656
rect 33463 6616 33508 6644
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 33594 6604 33600 6656
rect 33652 6644 33658 6656
rect 34977 6647 35035 6653
rect 34977 6644 34989 6647
rect 33652 6616 34989 6644
rect 33652 6604 33658 6616
rect 34977 6613 34989 6616
rect 35023 6613 35035 6647
rect 34977 6607 35035 6613
rect 1104 6554 36892 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 36892 6554
rect 1104 6480 36892 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 1854 6440 1860 6452
rect 1811 6412 1860 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 18598 6440 18604 6452
rect 18559 6412 18604 6440
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 20806 6440 20812 6452
rect 19812 6412 20812 6440
rect 17494 6332 17500 6384
rect 17552 6372 17558 6384
rect 19812 6372 19840 6412
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 22186 6400 22192 6452
rect 22244 6440 22250 6452
rect 24394 6440 24400 6452
rect 22244 6412 24400 6440
rect 22244 6400 22250 6412
rect 24394 6400 24400 6412
rect 24452 6400 24458 6452
rect 30374 6440 30380 6452
rect 24504 6412 30380 6440
rect 17552 6344 19656 6372
rect 17552 6332 17558 6344
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 17405 6307 17463 6313
rect 17405 6273 17417 6307
rect 17451 6304 17463 6307
rect 17957 6307 18015 6313
rect 17957 6304 17969 6307
rect 17451 6276 17969 6304
rect 17451 6273 17463 6276
rect 17405 6267 17463 6273
rect 17957 6273 17969 6276
rect 18003 6304 18015 6307
rect 18690 6304 18696 6316
rect 18003 6276 18696 6304
rect 18003 6273 18015 6276
rect 17957 6267 18015 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19024 6276 19257 6304
rect 19024 6264 19030 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18656 6208 19073 6236
rect 18656 6196 18662 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19628 6236 19656 6344
rect 19720 6344 19840 6372
rect 19981 6375 20039 6381
rect 19720 6313 19748 6344
rect 19981 6341 19993 6375
rect 20027 6372 20039 6375
rect 20254 6372 20260 6384
rect 20027 6344 20260 6372
rect 20027 6341 20039 6344
rect 19981 6335 20039 6341
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 24504 6372 24532 6412
rect 30374 6400 30380 6412
rect 30432 6400 30438 6452
rect 31386 6400 31392 6452
rect 31444 6440 31450 6452
rect 31665 6443 31723 6449
rect 31665 6440 31677 6443
rect 31444 6412 31677 6440
rect 31444 6400 31450 6412
rect 31665 6409 31677 6412
rect 31711 6409 31723 6443
rect 32582 6440 32588 6452
rect 32543 6412 32588 6440
rect 31665 6403 31723 6409
rect 32582 6400 32588 6412
rect 32640 6400 32646 6452
rect 32766 6400 32772 6452
rect 32824 6440 32830 6452
rect 33594 6440 33600 6452
rect 32824 6412 33600 6440
rect 32824 6400 32830 6412
rect 33594 6400 33600 6412
rect 33652 6400 33658 6452
rect 34514 6440 34520 6452
rect 34475 6412 34520 6440
rect 34514 6400 34520 6412
rect 34572 6400 34578 6452
rect 35526 6400 35532 6452
rect 35584 6440 35590 6452
rect 36265 6443 36323 6449
rect 36265 6440 36277 6443
rect 35584 6412 36277 6440
rect 35584 6400 35590 6412
rect 36265 6409 36277 6412
rect 36311 6409 36323 6443
rect 36265 6403 36323 6409
rect 21206 6344 22324 6372
rect 23138 6344 24532 6372
rect 24857 6375 24915 6381
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 22002 6304 22008 6316
rect 19705 6267 19763 6273
rect 21928 6276 22008 6304
rect 21928 6236 21956 6276
rect 22002 6264 22008 6276
rect 22060 6264 22066 6316
rect 22097 6239 22155 6245
rect 22097 6236 22109 6239
rect 19628 6208 21956 6236
rect 22020 6208 22109 6236
rect 19061 6199 19119 6205
rect 18049 6171 18107 6177
rect 18049 6137 18061 6171
rect 18095 6168 18107 6171
rect 19610 6168 19616 6180
rect 18095 6140 19616 6168
rect 18095 6137 18107 6140
rect 18049 6131 18107 6137
rect 19610 6128 19616 6140
rect 19668 6128 19674 6180
rect 22020 6168 22048 6208
rect 22097 6205 22109 6208
rect 22143 6205 22155 6239
rect 22097 6199 22155 6205
rect 21376 6140 22048 6168
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 21376 6100 21404 6140
rect 20496 6072 21404 6100
rect 21453 6103 21511 6109
rect 20496 6060 20502 6072
rect 21453 6069 21465 6103
rect 21499 6100 21511 6103
rect 22186 6100 22192 6112
rect 21499 6072 22192 6100
rect 21499 6069 21511 6072
rect 21453 6063 21511 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22296 6100 22324 6344
rect 24857 6341 24869 6375
rect 24903 6372 24915 6375
rect 24946 6372 24952 6384
rect 24903 6344 24952 6372
rect 24903 6341 24915 6344
rect 24857 6335 24915 6341
rect 24946 6332 24952 6344
rect 25004 6332 25010 6384
rect 27522 6372 27528 6384
rect 26082 6344 27528 6372
rect 27522 6332 27528 6344
rect 27580 6332 27586 6384
rect 33502 6372 33508 6384
rect 28842 6344 33508 6372
rect 33502 6332 33508 6344
rect 33560 6332 33566 6384
rect 35066 6372 35072 6384
rect 34624 6344 35072 6372
rect 23845 6307 23903 6313
rect 23845 6273 23857 6307
rect 23891 6304 23903 6307
rect 24026 6304 24032 6316
rect 23891 6276 24032 6304
rect 23891 6273 23903 6276
rect 23845 6267 23903 6273
rect 24026 6264 24032 6276
rect 24084 6304 24090 6316
rect 24581 6307 24639 6313
rect 24581 6304 24593 6307
rect 24084 6276 24593 6304
rect 24084 6264 24090 6276
rect 24581 6273 24593 6276
rect 24627 6273 24639 6307
rect 24581 6267 24639 6273
rect 26068 6276 27844 6304
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6236 23627 6239
rect 26068 6236 26096 6276
rect 26602 6236 26608 6248
rect 23615 6208 23888 6236
rect 23615 6205 23627 6208
rect 23569 6199 23627 6205
rect 23860 6180 23888 6208
rect 24596 6208 26096 6236
rect 26563 6208 26608 6236
rect 24596 6180 24624 6208
rect 26602 6196 26608 6208
rect 26660 6196 26666 6248
rect 27816 6245 27844 6276
rect 30558 6264 30564 6316
rect 30616 6304 30622 6316
rect 31757 6307 31815 6313
rect 31757 6304 31769 6307
rect 30616 6276 31769 6304
rect 30616 6264 30622 6276
rect 31757 6273 31769 6276
rect 31803 6304 31815 6307
rect 31846 6304 31852 6316
rect 31803 6276 31852 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 31846 6264 31852 6276
rect 31904 6264 31910 6316
rect 32674 6304 32680 6316
rect 32635 6276 32680 6304
rect 32674 6264 32680 6276
rect 32732 6264 32738 6316
rect 32858 6264 32864 6316
rect 32916 6304 32922 6316
rect 33321 6307 33379 6313
rect 33321 6304 33333 6307
rect 32916 6276 33333 6304
rect 32916 6264 32922 6276
rect 33321 6273 33333 6276
rect 33367 6304 33379 6307
rect 33686 6304 33692 6316
rect 33367 6276 33692 6304
rect 33367 6273 33379 6276
rect 33321 6267 33379 6273
rect 33686 6264 33692 6276
rect 33744 6304 33750 6316
rect 34624 6313 34652 6344
rect 35066 6332 35072 6344
rect 35124 6372 35130 6384
rect 35434 6372 35440 6384
rect 35124 6344 35440 6372
rect 35124 6332 35130 6344
rect 35434 6332 35440 6344
rect 35492 6372 35498 6384
rect 35713 6375 35771 6381
rect 35713 6372 35725 6375
rect 35492 6344 35725 6372
rect 35492 6332 35498 6344
rect 35713 6341 35725 6344
rect 35759 6341 35771 6375
rect 35713 6335 35771 6341
rect 33965 6307 34023 6313
rect 33965 6304 33977 6307
rect 33744 6276 33977 6304
rect 33744 6264 33750 6276
rect 33965 6273 33977 6276
rect 34011 6273 34023 6307
rect 34609 6307 34667 6313
rect 34609 6304 34621 6307
rect 33965 6267 34023 6273
rect 34072 6276 34621 6304
rect 27801 6239 27859 6245
rect 27801 6205 27813 6239
rect 27847 6205 27859 6239
rect 29270 6236 29276 6248
rect 29231 6208 29276 6236
rect 27801 6199 27859 6205
rect 29270 6196 29276 6208
rect 29328 6196 29334 6248
rect 29549 6239 29607 6245
rect 29549 6205 29561 6239
rect 29595 6205 29607 6239
rect 29549 6199 29607 6205
rect 23842 6128 23848 6180
rect 23900 6128 23906 6180
rect 24578 6128 24584 6180
rect 24636 6128 24642 6180
rect 26988 6140 28120 6168
rect 26988 6100 27016 6140
rect 27154 6100 27160 6112
rect 22296 6072 27016 6100
rect 27115 6072 27160 6100
rect 27154 6060 27160 6072
rect 27212 6060 27218 6112
rect 28092 6100 28120 6140
rect 29564 6112 29592 6199
rect 30466 6196 30472 6248
rect 30524 6236 30530 6248
rect 33229 6239 33287 6245
rect 33229 6236 33241 6239
rect 30524 6208 33241 6236
rect 30524 6196 30530 6208
rect 33229 6205 33241 6208
rect 33275 6205 33287 6239
rect 33229 6199 33287 6205
rect 29638 6128 29644 6180
rect 29696 6168 29702 6180
rect 33873 6171 33931 6177
rect 33873 6168 33885 6171
rect 29696 6140 33885 6168
rect 29696 6128 29702 6140
rect 33873 6137 33885 6140
rect 33919 6137 33931 6171
rect 33873 6131 33931 6137
rect 29178 6100 29184 6112
rect 28092 6072 29184 6100
rect 29178 6060 29184 6072
rect 29236 6060 29242 6112
rect 29546 6060 29552 6112
rect 29604 6100 29610 6112
rect 30009 6103 30067 6109
rect 30009 6100 30021 6103
rect 29604 6072 30021 6100
rect 29604 6060 29610 6072
rect 30009 6069 30021 6072
rect 30055 6069 30067 6103
rect 30009 6063 30067 6069
rect 30466 6060 30472 6112
rect 30524 6100 30530 6112
rect 30561 6103 30619 6109
rect 30561 6100 30573 6103
rect 30524 6072 30573 6100
rect 30524 6060 30530 6072
rect 30561 6069 30573 6072
rect 30607 6069 30619 6103
rect 30561 6063 30619 6069
rect 31570 6060 31576 6112
rect 31628 6100 31634 6112
rect 32582 6100 32588 6112
rect 31628 6072 32588 6100
rect 31628 6060 31634 6072
rect 32582 6060 32588 6072
rect 32640 6060 32646 6112
rect 32674 6060 32680 6112
rect 32732 6100 32738 6112
rect 34072 6100 34100 6276
rect 34609 6273 34621 6276
rect 34655 6273 34667 6307
rect 34609 6267 34667 6273
rect 35253 6307 35311 6313
rect 35253 6273 35265 6307
rect 35299 6273 35311 6307
rect 35253 6267 35311 6273
rect 34514 6196 34520 6248
rect 34572 6236 34578 6248
rect 34698 6236 34704 6248
rect 34572 6208 34704 6236
rect 34572 6196 34578 6208
rect 34698 6196 34704 6208
rect 34756 6236 34762 6248
rect 35268 6236 35296 6267
rect 34756 6208 35296 6236
rect 34756 6196 34762 6208
rect 32732 6072 34100 6100
rect 32732 6060 32738 6072
rect 34698 6060 34704 6112
rect 34756 6100 34762 6112
rect 35161 6103 35219 6109
rect 35161 6100 35173 6103
rect 34756 6072 35173 6100
rect 34756 6060 34762 6072
rect 35161 6069 35173 6072
rect 35207 6069 35219 6103
rect 35161 6063 35219 6069
rect 1104 6010 36892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36892 6010
rect 1104 5936 36892 5958
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 17313 5899 17371 5905
rect 17313 5865 17325 5899
rect 17359 5896 17371 5899
rect 17954 5896 17960 5908
rect 17359 5868 17960 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 18598 5896 18604 5908
rect 18559 5868 18604 5896
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 22094 5896 22100 5908
rect 20272 5868 22100 5896
rect 20272 5828 20300 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 23308 5868 28672 5896
rect 18524 5800 20300 5828
rect 20364 5800 20944 5828
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2314 5692 2320 5704
rect 1903 5664 2320 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 16684 5664 17233 5692
rect 16684 5568 16712 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 18524 5701 18552 5800
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 20364 5760 20392 5800
rect 20806 5760 20812 5772
rect 18748 5732 20392 5760
rect 20767 5732 20812 5760
rect 18748 5720 18754 5732
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 20916 5760 20944 5800
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 20916 5732 22845 5760
rect 22833 5729 22845 5732
rect 22879 5760 22891 5763
rect 22922 5760 22928 5772
rect 22879 5732 22928 5760
rect 22879 5729 22891 5732
rect 22833 5723 22891 5729
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17828 5664 17877 5692
rect 17828 5652 17834 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20346 5692 20352 5704
rect 20211 5664 20352 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 23308 5692 23336 5868
rect 23385 5831 23443 5837
rect 23385 5797 23397 5831
rect 23431 5828 23443 5831
rect 26602 5828 26608 5840
rect 23431 5800 26608 5828
rect 23431 5797 23443 5800
rect 23385 5791 23443 5797
rect 22218 5664 23336 5692
rect 19521 5627 19579 5633
rect 19521 5624 19533 5627
rect 17880 5596 19533 5624
rect 17880 5568 17908 5596
rect 19521 5593 19533 5596
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 19610 5584 19616 5636
rect 19668 5624 19674 5636
rect 19668 5596 19713 5624
rect 19668 5584 19674 5596
rect 20438 5584 20444 5636
rect 20496 5624 20502 5636
rect 21085 5627 21143 5633
rect 21085 5624 21097 5627
rect 20496 5596 21097 5624
rect 20496 5584 20502 5596
rect 21085 5593 21097 5596
rect 21131 5593 21143 5627
rect 21085 5587 21143 5593
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 16666 5556 16672 5568
rect 16627 5528 16672 5556
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 17862 5516 17868 5568
rect 17920 5516 17926 5568
rect 17957 5559 18015 5565
rect 17957 5525 17969 5559
rect 18003 5556 18015 5559
rect 18782 5556 18788 5568
rect 18003 5528 18788 5556
rect 18003 5525 18015 5528
rect 17957 5519 18015 5525
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 21174 5516 21180 5568
rect 21232 5556 21238 5568
rect 23400 5556 23428 5791
rect 26602 5788 26608 5800
rect 26660 5788 26666 5840
rect 27246 5828 27252 5840
rect 26712 5800 27252 5828
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 26712 5760 26740 5800
rect 27246 5788 27252 5800
rect 27304 5788 27310 5840
rect 23900 5732 26740 5760
rect 23900 5720 23906 5732
rect 27154 5720 27160 5772
rect 27212 5760 27218 5772
rect 27341 5763 27399 5769
rect 27341 5760 27353 5763
rect 27212 5732 27353 5760
rect 27212 5720 27218 5732
rect 27341 5729 27353 5732
rect 27387 5760 27399 5763
rect 28074 5760 28080 5772
rect 27387 5732 28080 5760
rect 27387 5729 27399 5732
rect 27341 5723 27399 5729
rect 28074 5720 28080 5732
rect 28132 5720 28138 5772
rect 28644 5760 28672 5868
rect 29086 5856 29092 5908
rect 29144 5896 29150 5908
rect 29990 5899 30048 5905
rect 29990 5896 30002 5899
rect 29144 5868 29189 5896
rect 29288 5868 30002 5896
rect 29144 5856 29150 5868
rect 28718 5788 28724 5840
rect 28776 5828 28782 5840
rect 29288 5828 29316 5868
rect 29990 5865 30002 5868
rect 30036 5865 30048 5899
rect 31478 5896 31484 5908
rect 31439 5868 31484 5896
rect 29990 5859 30048 5865
rect 31478 5856 31484 5868
rect 31536 5856 31542 5908
rect 32030 5896 32036 5908
rect 31991 5868 32036 5896
rect 32030 5856 32036 5868
rect 32088 5856 32094 5908
rect 32582 5856 32588 5908
rect 32640 5896 32646 5908
rect 32640 5868 32812 5896
rect 32640 5856 32646 5868
rect 28776 5800 29316 5828
rect 28776 5788 28782 5800
rect 31018 5788 31024 5840
rect 31076 5828 31082 5840
rect 32677 5831 32735 5837
rect 32677 5828 32689 5831
rect 31076 5800 32689 5828
rect 31076 5788 31082 5800
rect 32677 5797 32689 5800
rect 32723 5797 32735 5831
rect 32784 5828 32812 5868
rect 32950 5856 32956 5908
rect 33008 5896 33014 5908
rect 33321 5899 33379 5905
rect 33321 5896 33333 5899
rect 33008 5868 33333 5896
rect 33008 5856 33014 5868
rect 33321 5865 33333 5868
rect 33367 5865 33379 5899
rect 33321 5859 33379 5865
rect 33965 5831 34023 5837
rect 33965 5828 33977 5831
rect 32784 5800 33977 5828
rect 32677 5791 32735 5797
rect 33965 5797 33977 5800
rect 34011 5797 34023 5831
rect 33965 5791 34023 5797
rect 32306 5760 32312 5772
rect 28644 5732 32312 5760
rect 32306 5720 32312 5732
rect 32364 5720 32370 5772
rect 32692 5732 32996 5760
rect 25682 5652 25688 5704
rect 25740 5692 25746 5704
rect 25740 5664 27384 5692
rect 25740 5652 25746 5664
rect 23937 5627 23995 5633
rect 23937 5593 23949 5627
rect 23983 5624 23995 5627
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 23983 5596 24685 5624
rect 23983 5593 23995 5596
rect 23937 5587 23995 5593
rect 24673 5593 24685 5596
rect 24719 5624 24731 5627
rect 24719 5596 26096 5624
rect 24719 5593 24731 5596
rect 24673 5587 24731 5593
rect 26068 5568 26096 5596
rect 26142 5584 26148 5636
rect 26200 5624 26206 5636
rect 26697 5627 26755 5633
rect 26697 5624 26709 5627
rect 26200 5596 26709 5624
rect 26200 5584 26206 5596
rect 26697 5593 26709 5596
rect 26743 5593 26755 5627
rect 26697 5587 26755 5593
rect 25498 5556 25504 5568
rect 21232 5528 23428 5556
rect 25459 5528 25504 5556
rect 21232 5516 21238 5528
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 26050 5556 26056 5568
rect 26011 5528 26056 5556
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 27356 5556 27384 5664
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 29733 5695 29791 5701
rect 29733 5692 29745 5695
rect 29696 5664 29745 5692
rect 29696 5652 29702 5664
rect 29733 5661 29745 5664
rect 29779 5661 29791 5695
rect 29733 5655 29791 5661
rect 31110 5652 31116 5704
rect 31168 5652 31174 5704
rect 31662 5652 31668 5704
rect 31720 5692 31726 5704
rect 32125 5695 32183 5701
rect 32125 5692 32137 5695
rect 31720 5664 32137 5692
rect 31720 5652 31726 5664
rect 32125 5661 32137 5664
rect 32171 5692 32183 5695
rect 32692 5692 32720 5732
rect 32171 5664 32720 5692
rect 32769 5695 32827 5701
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 32769 5661 32781 5695
rect 32815 5661 32827 5695
rect 32968 5692 32996 5732
rect 33134 5720 33140 5772
rect 33192 5760 33198 5772
rect 36081 5763 36139 5769
rect 36081 5760 36093 5763
rect 33192 5732 36093 5760
rect 33192 5720 33198 5732
rect 36081 5729 36093 5732
rect 36127 5729 36139 5763
rect 36081 5723 36139 5729
rect 33413 5695 33471 5701
rect 33413 5692 33425 5695
rect 32968 5664 33425 5692
rect 32769 5655 32827 5661
rect 33413 5661 33425 5664
rect 33459 5692 33471 5695
rect 33778 5692 33784 5704
rect 33459 5664 33784 5692
rect 33459 5661 33471 5664
rect 33413 5655 33471 5661
rect 27614 5624 27620 5636
rect 27575 5596 27620 5624
rect 27614 5584 27620 5596
rect 27672 5584 27678 5636
rect 28842 5596 29960 5624
rect 29822 5556 29828 5568
rect 27356 5528 29828 5556
rect 29822 5516 29828 5528
rect 29880 5516 29886 5568
rect 29932 5556 29960 5596
rect 31312 5596 31754 5624
rect 31312 5556 31340 5596
rect 29932 5528 31340 5556
rect 31726 5568 31754 5596
rect 32674 5584 32680 5636
rect 32732 5624 32738 5636
rect 32784 5624 32812 5655
rect 33778 5652 33784 5664
rect 33836 5652 33842 5704
rect 34054 5692 34060 5704
rect 34015 5664 34060 5692
rect 34054 5652 34060 5664
rect 34112 5652 34118 5704
rect 35069 5695 35127 5701
rect 35069 5661 35081 5695
rect 35115 5692 35127 5695
rect 35434 5692 35440 5704
rect 35115 5664 35440 5692
rect 35115 5661 35127 5664
rect 35069 5655 35127 5661
rect 35434 5652 35440 5664
rect 35492 5652 35498 5704
rect 36354 5692 36360 5704
rect 36315 5664 36360 5692
rect 36354 5652 36360 5664
rect 36412 5652 36418 5704
rect 32732 5596 32812 5624
rect 32732 5584 32738 5596
rect 31726 5528 31760 5568
rect 31754 5516 31760 5528
rect 31812 5516 31818 5568
rect 33134 5516 33140 5568
rect 33192 5556 33198 5568
rect 34977 5559 35035 5565
rect 34977 5556 34989 5559
rect 33192 5528 34989 5556
rect 33192 5516 33198 5528
rect 34977 5525 34989 5528
rect 35023 5525 35035 5559
rect 34977 5519 35035 5525
rect 1104 5466 36892 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 36892 5466
rect 1104 5392 36892 5414
rect 19061 5355 19119 5361
rect 19061 5321 19073 5355
rect 19107 5352 19119 5355
rect 19150 5352 19156 5364
rect 19107 5324 19156 5352
rect 19107 5321 19119 5324
rect 19061 5315 19119 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 19978 5352 19984 5364
rect 19751 5324 19984 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 22002 5312 22008 5364
rect 22060 5352 22066 5364
rect 28905 5355 28963 5361
rect 22060 5324 23060 5352
rect 22060 5312 22066 5324
rect 16758 5244 16764 5296
rect 16816 5284 16822 5296
rect 17405 5287 17463 5293
rect 17405 5284 17417 5287
rect 16816 5256 17417 5284
rect 16816 5244 16822 5256
rect 17405 5253 17417 5256
rect 17451 5253 17463 5287
rect 17405 5247 17463 5253
rect 18325 5287 18383 5293
rect 18325 5253 18337 5287
rect 18371 5284 18383 5287
rect 20070 5284 20076 5296
rect 18371 5256 20076 5284
rect 18371 5253 18383 5256
rect 18325 5247 18383 5253
rect 20070 5244 20076 5256
rect 20128 5244 20134 5296
rect 13538 5176 13544 5228
rect 13596 5216 13602 5228
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 13596 5188 14565 5216
rect 13596 5176 13602 5188
rect 14553 5185 14565 5188
rect 14599 5216 14611 5219
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 14599 5188 15209 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 15197 5179 15255 5185
rect 18156 5188 18981 5216
rect 17310 5148 17316 5160
rect 17271 5120 17316 5148
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 18156 5148 18184 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5185 19671 5219
rect 19613 5179 19671 5185
rect 18012 5120 18184 5148
rect 19628 5148 19656 5179
rect 22922 5148 22928 5160
rect 19628 5120 22928 5148
rect 18012 5108 18018 5120
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 15286 5080 15292 5092
rect 14691 5052 15292 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 15286 5040 15292 5052
rect 15344 5040 15350 5092
rect 17586 5040 17592 5092
rect 17644 5080 17650 5092
rect 19628 5080 19656 5120
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 17644 5052 19656 5080
rect 17644 5040 17650 5052
rect 20806 5040 20812 5092
rect 20864 5080 20870 5092
rect 22002 5080 22008 5092
rect 20864 5052 22008 5080
rect 20864 5040 20870 5052
rect 22002 5040 22008 5052
rect 22060 5040 22066 5092
rect 23032 5021 23060 5324
rect 28905 5321 28917 5355
rect 28951 5352 28963 5355
rect 28994 5352 29000 5364
rect 28951 5324 29000 5352
rect 28951 5321 28963 5324
rect 28905 5315 28963 5321
rect 28994 5312 29000 5324
rect 29052 5312 29058 5364
rect 33042 5352 33048 5364
rect 30116 5324 33048 5352
rect 30116 5284 30144 5324
rect 33042 5312 33048 5324
rect 33100 5312 33106 5364
rect 33778 5312 33784 5364
rect 33836 5352 33842 5364
rect 34241 5355 34299 5361
rect 34241 5352 34253 5355
rect 33836 5324 34253 5352
rect 33836 5312 33842 5324
rect 34241 5321 34253 5324
rect 34287 5352 34299 5355
rect 34422 5352 34428 5364
rect 34287 5324 34428 5352
rect 34287 5321 34299 5324
rect 34241 5315 34299 5321
rect 34422 5312 34428 5324
rect 34480 5312 34486 5364
rect 34885 5355 34943 5361
rect 34885 5321 34897 5355
rect 34931 5352 34943 5355
rect 35434 5352 35440 5364
rect 34931 5324 35440 5352
rect 34931 5321 34943 5324
rect 34885 5315 34943 5321
rect 35434 5312 35440 5324
rect 35492 5312 35498 5364
rect 28828 5256 30144 5284
rect 27154 5216 27160 5228
rect 27115 5188 27160 5216
rect 27154 5176 27160 5188
rect 27212 5176 27218 5228
rect 28828 5216 28856 5256
rect 30374 5244 30380 5296
rect 30432 5284 30438 5296
rect 30432 5256 30477 5284
rect 30432 5244 30438 5256
rect 30558 5244 30564 5296
rect 30616 5284 30622 5296
rect 30742 5284 30748 5296
rect 30616 5256 30748 5284
rect 30616 5244 30622 5256
rect 30742 5244 30748 5256
rect 30800 5284 30806 5296
rect 31662 5284 31668 5296
rect 30800 5256 31668 5284
rect 30800 5244 30806 5256
rect 28566 5188 28856 5216
rect 29086 5176 29092 5228
rect 29144 5216 29150 5228
rect 30098 5216 30104 5228
rect 29144 5188 30104 5216
rect 29144 5176 29150 5188
rect 30098 5176 30104 5188
rect 30156 5176 30162 5228
rect 30466 5216 30472 5228
rect 30427 5188 30472 5216
rect 30466 5176 30472 5188
rect 30524 5176 30530 5228
rect 31128 5225 31156 5256
rect 31662 5244 31668 5256
rect 31720 5284 31726 5296
rect 31720 5256 32536 5284
rect 31720 5244 31726 5256
rect 31021 5219 31079 5225
rect 31021 5216 31033 5219
rect 30576 5188 31033 5216
rect 27522 5108 27528 5160
rect 27580 5148 27586 5160
rect 27580 5120 28856 5148
rect 27580 5108 27586 5120
rect 24949 5083 25007 5089
rect 24949 5049 24961 5083
rect 24995 5080 25007 5083
rect 26418 5080 26424 5092
rect 24995 5052 26424 5080
rect 24995 5049 25007 5052
rect 24949 5043 25007 5049
rect 26418 5040 26424 5052
rect 26476 5040 26482 5092
rect 28828 5080 28856 5120
rect 29178 5108 29184 5160
rect 29236 5148 29242 5160
rect 30576 5148 30604 5188
rect 31021 5185 31033 5188
rect 31067 5185 31079 5219
rect 31021 5179 31079 5185
rect 31113 5219 31171 5225
rect 31113 5185 31125 5219
rect 31159 5185 31171 5219
rect 31754 5216 31760 5228
rect 31715 5188 31760 5216
rect 31113 5179 31171 5185
rect 31754 5176 31760 5188
rect 31812 5176 31818 5228
rect 32398 5216 32404 5228
rect 32359 5188 32404 5216
rect 32398 5176 32404 5188
rect 32456 5176 32462 5228
rect 32508 5225 32536 5256
rect 32858 5244 32864 5296
rect 32916 5284 32922 5296
rect 32916 5256 33824 5284
rect 32916 5244 32922 5256
rect 32493 5219 32551 5225
rect 32493 5185 32505 5219
rect 32539 5185 32551 5219
rect 32493 5179 32551 5185
rect 33137 5219 33195 5225
rect 33137 5185 33149 5219
rect 33183 5216 33195 5219
rect 33226 5216 33232 5228
rect 33183 5188 33232 5216
rect 33183 5185 33195 5188
rect 33137 5179 33195 5185
rect 33226 5176 33232 5188
rect 33284 5216 33290 5228
rect 33502 5216 33508 5228
rect 33284 5188 33508 5216
rect 33284 5176 33290 5188
rect 33502 5176 33508 5188
rect 33560 5176 33566 5228
rect 33796 5225 33824 5256
rect 33781 5219 33839 5225
rect 33781 5185 33793 5219
rect 33827 5185 33839 5219
rect 33781 5179 33839 5185
rect 34054 5176 34060 5228
rect 34112 5216 34118 5228
rect 35897 5219 35955 5225
rect 35897 5216 35909 5219
rect 34112 5188 35909 5216
rect 34112 5176 34118 5188
rect 35897 5185 35909 5188
rect 35943 5185 35955 5219
rect 35897 5179 35955 5185
rect 29236 5120 30604 5148
rect 29236 5108 29242 5120
rect 30742 5108 30748 5160
rect 30800 5148 30806 5160
rect 33689 5151 33747 5157
rect 33689 5148 33701 5151
rect 30800 5120 33701 5148
rect 30800 5108 30806 5120
rect 33689 5117 33701 5120
rect 33735 5117 33747 5151
rect 33689 5111 33747 5117
rect 32582 5080 32588 5092
rect 28828 5052 32588 5080
rect 32582 5040 32588 5052
rect 32640 5040 32646 5092
rect 33042 5080 33048 5092
rect 33003 5052 33048 5080
rect 33042 5040 33048 5052
rect 33100 5040 33106 5092
rect 33502 5040 33508 5092
rect 33560 5080 33566 5092
rect 34054 5080 34060 5092
rect 33560 5052 34060 5080
rect 33560 5040 33566 5052
rect 34054 5040 34060 5052
rect 34112 5040 34118 5092
rect 23017 5015 23075 5021
rect 23017 4981 23029 5015
rect 23063 5012 23075 5015
rect 23658 5012 23664 5024
rect 23063 4984 23664 5012
rect 23063 4981 23075 4984
rect 23017 4975 23075 4981
rect 23658 4972 23664 4984
rect 23716 4972 23722 5024
rect 24118 5012 24124 5024
rect 24079 4984 24124 5012
rect 24118 4972 24124 4984
rect 24176 4972 24182 5024
rect 25501 5015 25559 5021
rect 25501 4981 25513 5015
rect 25547 5012 25559 5015
rect 26050 5012 26056 5024
rect 25547 4984 26056 5012
rect 25547 4981 25559 4984
rect 25501 4975 25559 4981
rect 26050 4972 26056 4984
rect 26108 5012 26114 5024
rect 26513 5015 26571 5021
rect 26513 5012 26525 5015
rect 26108 4984 26525 5012
rect 26108 4972 26114 4984
rect 26513 4981 26525 4984
rect 26559 4981 26571 5015
rect 26513 4975 26571 4981
rect 27420 5015 27478 5021
rect 27420 4981 27432 5015
rect 27466 5012 27478 5015
rect 29086 5012 29092 5024
rect 27466 4984 29092 5012
rect 27466 4981 27478 4984
rect 27420 4975 27478 4981
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 29638 5012 29644 5024
rect 29599 4984 29644 5012
rect 29638 4972 29644 4984
rect 29696 4972 29702 5024
rect 29822 4972 29828 5024
rect 29880 5012 29886 5024
rect 31665 5015 31723 5021
rect 31665 5012 31677 5015
rect 29880 4984 31677 5012
rect 29880 4972 29886 4984
rect 31665 4981 31677 4984
rect 31711 4981 31723 5015
rect 31665 4975 31723 4981
rect 1104 4922 36892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36892 4922
rect 1104 4848 36892 4870
rect 16758 4808 16764 4820
rect 16719 4780 16764 4808
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 22646 4808 22652 4820
rect 17144 4780 22508 4808
rect 22607 4780 22652 4808
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 17144 4672 17172 4780
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 18141 4743 18199 4749
rect 18141 4740 18153 4743
rect 17828 4712 18153 4740
rect 17828 4700 17834 4712
rect 18141 4709 18153 4712
rect 18187 4709 18199 4743
rect 22480 4740 22508 4780
rect 22646 4768 22652 4780
rect 22704 4768 22710 4820
rect 22756 4780 24164 4808
rect 22756 4740 22784 4780
rect 22480 4712 22784 4740
rect 24136 4740 24164 4780
rect 25222 4768 25228 4820
rect 25280 4808 25286 4820
rect 33042 4808 33048 4820
rect 25280 4780 33048 4808
rect 25280 4768 25286 4780
rect 33042 4768 33048 4780
rect 33100 4768 33106 4820
rect 35434 4808 35440 4820
rect 35395 4780 35440 4808
rect 35434 4768 35440 4780
rect 35492 4768 35498 4820
rect 24136 4712 27463 4740
rect 18141 4703 18199 4709
rect 17310 4672 17316 4684
rect 15151 4644 17172 4672
rect 17271 4644 17316 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20864 4644 20913 4672
rect 20864 4632 20870 4644
rect 20901 4641 20913 4644
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 21177 4675 21235 4681
rect 21177 4641 21189 4675
rect 21223 4672 21235 4675
rect 21634 4672 21640 4684
rect 21223 4644 21640 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 21634 4632 21640 4644
rect 21692 4672 21698 4684
rect 23109 4675 23167 4681
rect 23109 4672 23121 4675
rect 21692 4644 23121 4672
rect 21692 4632 21698 4644
rect 23109 4641 23121 4644
rect 23155 4641 23167 4675
rect 23109 4635 23167 4641
rect 23658 4632 23664 4684
rect 23716 4672 23722 4684
rect 23753 4675 23811 4681
rect 23753 4672 23765 4675
rect 23716 4644 23765 4672
rect 23716 4632 23722 4644
rect 23753 4641 23765 4644
rect 23799 4672 23811 4675
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 23799 4644 24685 4672
rect 23799 4641 23811 4644
rect 23753 4635 23811 4641
rect 24673 4641 24685 4644
rect 24719 4672 24731 4675
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 24719 4644 25237 4672
rect 24719 4641 24731 4644
rect 24673 4635 24731 4641
rect 25225 4641 25237 4644
rect 25271 4672 25283 4675
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 25271 4644 25789 4672
rect 25271 4641 25283 4644
rect 25225 4635 25283 4641
rect 25777 4641 25789 4644
rect 25823 4672 25835 4675
rect 26050 4672 26056 4684
rect 25823 4644 26056 4672
rect 25823 4641 25835 4644
rect 25777 4635 25835 4641
rect 26050 4632 26056 4644
rect 26108 4672 26114 4684
rect 26329 4675 26387 4681
rect 26329 4672 26341 4675
rect 26108 4644 26341 4672
rect 26108 4632 26114 4644
rect 26329 4641 26341 4644
rect 26375 4672 26387 4675
rect 26881 4675 26939 4681
rect 26881 4672 26893 4675
rect 26375 4644 26893 4672
rect 26375 4641 26387 4644
rect 26329 4635 26387 4641
rect 26881 4641 26893 4644
rect 26927 4672 26939 4675
rect 27154 4672 27160 4684
rect 26927 4644 27160 4672
rect 26927 4641 26939 4644
rect 26881 4635 26939 4641
rect 27154 4632 27160 4644
rect 27212 4672 27218 4684
rect 27341 4675 27399 4681
rect 27341 4672 27353 4675
rect 27212 4644 27353 4672
rect 27212 4632 27218 4644
rect 27341 4641 27353 4644
rect 27387 4641 27399 4675
rect 27435 4672 27463 4712
rect 29086 4700 29092 4752
rect 29144 4740 29150 4752
rect 29730 4740 29736 4752
rect 29144 4712 29736 4740
rect 29144 4700 29150 4712
rect 29730 4700 29736 4712
rect 29788 4700 29794 4752
rect 31478 4700 31484 4752
rect 31536 4700 31542 4752
rect 30466 4672 30472 4684
rect 27435 4644 30472 4672
rect 27341 4635 27399 4641
rect 30466 4632 30472 4644
rect 30524 4632 30530 4684
rect 31205 4675 31263 4681
rect 31205 4641 31217 4675
rect 31251 4672 31263 4675
rect 31496 4672 31524 4700
rect 32582 4672 32588 4684
rect 31251 4644 31524 4672
rect 32543 4644 32588 4672
rect 31251 4641 31263 4644
rect 31205 4635 31263 4641
rect 32582 4632 32588 4644
rect 32640 4632 32646 4684
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13538 4604 13544 4616
rect 13127 4576 13544 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13538 4564 13544 4576
rect 13596 4604 13602 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13596 4576 14289 4604
rect 13596 4564 13602 4576
rect 14277 4573 14289 4576
rect 14323 4604 14335 4607
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 14323 4576 14841 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 19242 4604 19248 4616
rect 16899 4576 19248 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 29914 4604 29920 4616
rect 28750 4576 29920 4604
rect 29914 4564 29920 4576
rect 29972 4564 29978 4616
rect 31481 4607 31539 4613
rect 31481 4573 31493 4607
rect 31527 4573 31539 4607
rect 31481 4567 31539 4573
rect 13633 4539 13691 4545
rect 13633 4505 13645 4539
rect 13679 4536 13691 4539
rect 25222 4536 25228 4548
rect 13679 4508 21128 4536
rect 22402 4508 25228 4536
rect 13679 4505 13691 4508
rect 13633 4499 13691 4505
rect 21100 4468 21128 4508
rect 25222 4496 25228 4508
rect 25280 4496 25286 4548
rect 26326 4496 26332 4548
rect 26384 4536 26390 4548
rect 27614 4536 27620 4548
rect 26384 4508 27620 4536
rect 26384 4496 26390 4508
rect 27614 4496 27620 4508
rect 27672 4496 27678 4548
rect 29012 4508 29960 4536
rect 21450 4468 21456 4480
rect 21100 4440 21456 4468
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 25314 4428 25320 4480
rect 25372 4468 25378 4480
rect 29012 4468 29040 4508
rect 25372 4440 29040 4468
rect 29089 4471 29147 4477
rect 25372 4428 25378 4440
rect 29089 4437 29101 4471
rect 29135 4468 29147 4471
rect 29362 4468 29368 4480
rect 29135 4440 29368 4468
rect 29135 4437 29147 4440
rect 29089 4431 29147 4437
rect 29362 4428 29368 4440
rect 29420 4428 29426 4480
rect 29932 4468 29960 4508
rect 30742 4496 30748 4548
rect 30800 4496 30806 4548
rect 31496 4536 31524 4567
rect 31754 4564 31760 4616
rect 31812 4604 31818 4616
rect 32674 4604 32680 4616
rect 31812 4576 32680 4604
rect 31812 4564 31818 4576
rect 32674 4564 32680 4576
rect 32732 4564 32738 4616
rect 33321 4607 33379 4613
rect 33321 4573 33333 4607
rect 33367 4604 33379 4607
rect 33502 4604 33508 4616
rect 33367 4576 33508 4604
rect 33367 4573 33379 4576
rect 33321 4567 33379 4573
rect 33502 4564 33508 4576
rect 33560 4564 33566 4616
rect 33778 4564 33784 4616
rect 33836 4604 33842 4616
rect 33965 4607 34023 4613
rect 33965 4604 33977 4607
rect 33836 4576 33977 4604
rect 33836 4564 33842 4576
rect 33965 4573 33977 4576
rect 34011 4604 34023 4607
rect 34885 4607 34943 4613
rect 34885 4604 34897 4607
rect 34011 4576 34897 4604
rect 34011 4573 34023 4576
rect 33965 4567 34023 4573
rect 34885 4573 34897 4576
rect 34931 4573 34943 4607
rect 34885 4567 34943 4573
rect 35894 4564 35900 4616
rect 35952 4604 35958 4616
rect 36081 4607 36139 4613
rect 36081 4604 36093 4607
rect 35952 4576 36093 4604
rect 35952 4564 35958 4576
rect 36081 4573 36093 4576
rect 36127 4573 36139 4607
rect 36081 4567 36139 4573
rect 31496 4508 32076 4536
rect 32048 4480 32076 4508
rect 31478 4468 31484 4480
rect 29932 4440 31484 4468
rect 31478 4428 31484 4440
rect 31536 4428 31542 4480
rect 32030 4468 32036 4480
rect 31991 4440 32036 4468
rect 32030 4428 32036 4440
rect 32088 4428 32094 4480
rect 32692 4468 32720 4564
rect 33226 4536 33232 4548
rect 33187 4508 33232 4536
rect 33226 4496 33232 4508
rect 33284 4496 33290 4548
rect 33318 4468 33324 4480
rect 32692 4440 33324 4468
rect 33318 4428 33324 4440
rect 33376 4428 33382 4480
rect 33870 4468 33876 4480
rect 33831 4440 33876 4468
rect 33870 4428 33876 4440
rect 33928 4428 33934 4480
rect 36262 4468 36268 4480
rect 36223 4440 36268 4468
rect 36262 4428 36268 4440
rect 36320 4428 36326 4480
rect 1104 4378 36892 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 36892 4378
rect 1104 4304 36892 4326
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 13538 4264 13544 4276
rect 13495 4236 13544 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 21361 4267 21419 4273
rect 21361 4264 21373 4267
rect 20864 4236 21373 4264
rect 20864 4224 20870 4236
rect 21361 4233 21373 4236
rect 21407 4233 21419 4267
rect 32674 4264 32680 4276
rect 21361 4227 21419 4233
rect 24504 4236 32680 4264
rect 13556 4128 13584 4224
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13556 4100 13921 4128
rect 13909 4097 13921 4100
rect 13955 4128 13967 4131
rect 14829 4131 14887 4137
rect 14829 4128 14841 4131
rect 13955 4100 14841 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 14829 4097 14841 4100
rect 14875 4128 14887 4131
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 14875 4100 15761 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17736 4100 17785 4128
rect 17736 4088 17742 4100
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18966 4128 18972 4140
rect 17920 4100 17965 4128
rect 18927 4100 18972 4128
rect 17920 4088 17926 4100
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 21376 4128 21404 4227
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 22370 4196 22376 4208
rect 21508 4168 22376 4196
rect 21508 4156 21514 4168
rect 22370 4156 22376 4168
rect 22428 4156 22434 4208
rect 24504 4196 24532 4236
rect 32674 4224 32680 4236
rect 32732 4224 32738 4276
rect 32858 4224 32864 4276
rect 32916 4264 32922 4276
rect 32916 4236 34836 4264
rect 32916 4224 32922 4236
rect 23598 4168 24532 4196
rect 25314 4156 25320 4208
rect 25372 4156 25378 4208
rect 28442 4156 28448 4208
rect 28500 4156 28506 4208
rect 28994 4156 29000 4208
rect 29052 4196 29058 4208
rect 29917 4199 29975 4205
rect 29917 4196 29929 4199
rect 29052 4168 29929 4196
rect 29052 4156 29058 4168
rect 29917 4165 29929 4168
rect 29963 4165 29975 4199
rect 34698 4196 34704 4208
rect 31142 4168 34704 4196
rect 29917 4159 29975 4165
rect 34698 4156 34704 4168
rect 34756 4156 34762 4208
rect 22097 4131 22155 4137
rect 22097 4128 22109 4131
rect 19116 4100 19161 4128
rect 21376 4100 22109 4128
rect 19116 4088 19122 4100
rect 22097 4097 22109 4100
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 26050 4088 26056 4140
rect 26108 4128 26114 4140
rect 26513 4131 26571 4137
rect 26513 4128 26525 4131
rect 26108 4100 26525 4128
rect 26108 4088 26114 4100
rect 26513 4097 26525 4100
rect 26559 4097 26571 4131
rect 26513 4091 26571 4097
rect 26602 4088 26608 4140
rect 26660 4128 26666 4140
rect 26660 4100 27752 4128
rect 26660 4088 26666 4100
rect 14182 4060 14188 4072
rect 14143 4032 14188 4060
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 22373 4063 22431 4069
rect 15151 4032 22094 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 21634 3924 21640 3936
rect 18012 3896 21640 3924
rect 18012 3884 18018 3896
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 22066 3924 22094 4032
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 22830 4060 22836 4072
rect 22419 4032 22836 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22830 4020 22836 4032
rect 22888 4020 22894 4072
rect 22922 4020 22928 4072
rect 22980 4060 22986 4072
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 22980 4032 24317 4060
rect 22980 4020 22986 4032
rect 24305 4029 24317 4032
rect 24351 4029 24363 4063
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 24305 4023 24363 4029
rect 24780 4032 25789 4060
rect 23474 3952 23480 4004
rect 23532 3992 23538 4004
rect 24780 3992 24808 4032
rect 25777 4029 25789 4032
rect 25823 4060 25835 4063
rect 26234 4060 26240 4072
rect 25823 4032 26240 4060
rect 25823 4029 25835 4032
rect 25777 4023 25835 4029
rect 26234 4020 26240 4032
rect 26292 4020 26298 4072
rect 27430 4060 27436 4072
rect 27391 4032 27436 4060
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 27724 4060 27752 4100
rect 31202 4088 31208 4140
rect 31260 4128 31266 4140
rect 31260 4100 31754 4128
rect 31260 4088 31266 4100
rect 28442 4060 28448 4072
rect 27724 4032 28448 4060
rect 28442 4020 28448 4032
rect 28500 4020 28506 4072
rect 28902 4060 28908 4072
rect 28863 4032 28908 4060
rect 28902 4020 28908 4032
rect 28960 4020 28966 4072
rect 29178 4060 29184 4072
rect 29091 4032 29184 4060
rect 29178 4020 29184 4032
rect 29236 4060 29242 4072
rect 29638 4060 29644 4072
rect 29236 4032 29644 4060
rect 29236 4020 29242 4032
rect 29638 4020 29644 4032
rect 29696 4020 29702 4072
rect 31570 4060 31576 4072
rect 29748 4032 31576 4060
rect 29748 3992 29776 4032
rect 31570 4020 31576 4032
rect 31628 4020 31634 4072
rect 31726 4060 31754 4100
rect 32306 4088 32312 4140
rect 32364 4128 32370 4140
rect 32401 4131 32459 4137
rect 32401 4128 32413 4131
rect 32364 4100 32413 4128
rect 32364 4088 32370 4100
rect 32401 4097 32413 4100
rect 32447 4097 32459 4131
rect 32401 4091 32459 4097
rect 32493 4131 32551 4137
rect 32493 4097 32505 4131
rect 32539 4128 32551 4131
rect 32858 4128 32864 4140
rect 32539 4100 32864 4128
rect 32539 4097 32551 4100
rect 32493 4091 32551 4097
rect 32858 4088 32864 4100
rect 32916 4088 32922 4140
rect 33042 4128 33048 4140
rect 33003 4100 33048 4128
rect 33042 4088 33048 4100
rect 33100 4088 33106 4140
rect 33137 4131 33195 4137
rect 33137 4097 33149 4131
rect 33183 4128 33195 4131
rect 33318 4128 33324 4140
rect 33183 4100 33324 4128
rect 33183 4097 33195 4100
rect 33137 4091 33195 4097
rect 33318 4088 33324 4100
rect 33376 4088 33382 4140
rect 33778 4128 33784 4140
rect 33739 4100 33784 4128
rect 33778 4088 33784 4100
rect 33836 4088 33842 4140
rect 34808 4128 34836 4236
rect 35897 4131 35955 4137
rect 35897 4128 35909 4131
rect 34808 4100 35909 4128
rect 35897 4097 35909 4100
rect 35943 4097 35955 4131
rect 35897 4091 35955 4097
rect 34698 4060 34704 4072
rect 31726 4032 34704 4060
rect 34698 4020 34704 4032
rect 34756 4020 34762 4072
rect 32030 3992 32036 4004
rect 23532 3964 24808 3992
rect 27356 3964 27936 3992
rect 23532 3952 23538 3964
rect 23750 3924 23756 3936
rect 22066 3896 23756 3924
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3924 23903 3927
rect 24302 3924 24308 3936
rect 23891 3896 24308 3924
rect 23891 3893 23903 3896
rect 23845 3887 23903 3893
rect 24302 3884 24308 3896
rect 24360 3884 24366 3936
rect 24394 3884 24400 3936
rect 24452 3924 24458 3936
rect 27356 3924 27384 3964
rect 24452 3896 27384 3924
rect 27908 3924 27936 3964
rect 29564 3964 29776 3992
rect 30944 3964 32036 3992
rect 29564 3924 29592 3964
rect 27908 3896 29592 3924
rect 24452 3884 24458 3896
rect 29638 3884 29644 3936
rect 29696 3924 29702 3936
rect 30944 3924 30972 3964
rect 32030 3952 32036 3964
rect 32088 3992 32094 4004
rect 34333 3995 34391 4001
rect 34333 3992 34345 3995
rect 32088 3964 34345 3992
rect 32088 3952 32094 3964
rect 34333 3961 34345 3964
rect 34379 3992 34391 3995
rect 35986 3992 35992 4004
rect 34379 3964 35992 3992
rect 34379 3961 34391 3964
rect 34333 3955 34391 3961
rect 35986 3952 35992 3964
rect 36044 3952 36050 4004
rect 29696 3896 30972 3924
rect 29696 3884 29702 3896
rect 31202 3884 31208 3936
rect 31260 3924 31266 3936
rect 31389 3927 31447 3933
rect 31389 3924 31401 3927
rect 31260 3896 31401 3924
rect 31260 3884 31266 3896
rect 31389 3893 31401 3896
rect 31435 3893 31447 3927
rect 33686 3924 33692 3936
rect 33647 3896 33692 3924
rect 31389 3887 31447 3893
rect 33686 3884 33692 3896
rect 33744 3884 33750 3936
rect 33778 3884 33784 3936
rect 33836 3924 33842 3936
rect 34793 3927 34851 3933
rect 34793 3924 34805 3927
rect 33836 3896 34805 3924
rect 33836 3884 33842 3896
rect 34793 3893 34805 3896
rect 34839 3893 34851 3927
rect 35434 3924 35440 3936
rect 35395 3896 35440 3924
rect 34793 3887 34851 3893
rect 35434 3884 35440 3896
rect 35492 3884 35498 3936
rect 1104 3834 36892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36892 3834
rect 1104 3760 36892 3782
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 13596 3692 14289 3720
rect 13596 3680 13602 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 20441 3723 20499 3729
rect 20441 3689 20453 3723
rect 20487 3720 20499 3723
rect 20806 3720 20812 3732
rect 20487 3692 20812 3720
rect 20487 3689 20499 3692
rect 20441 3683 20499 3689
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 6886 3624 10333 3652
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 6886 3516 6914 3624
rect 10321 3621 10333 3624
rect 10367 3621 10379 3655
rect 10321 3615 10379 3621
rect 1903 3488 6914 3516
rect 10505 3519 10563 3525
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 14292 3516 14320 3683
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 29089 3723 29147 3729
rect 20916 3692 28120 3720
rect 20916 3652 20944 3692
rect 15120 3624 20944 3652
rect 15120 3593 15148 3624
rect 22554 3612 22560 3664
rect 22612 3652 22618 3664
rect 22649 3655 22707 3661
rect 22649 3652 22661 3655
rect 22612 3624 22661 3652
rect 22612 3612 22618 3624
rect 22649 3621 22661 3624
rect 22695 3652 22707 3655
rect 28092 3652 28120 3692
rect 29089 3689 29101 3723
rect 29135 3720 29147 3723
rect 29178 3720 29184 3732
rect 29135 3692 29184 3720
rect 29135 3689 29147 3692
rect 29089 3683 29147 3689
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 31386 3720 31392 3732
rect 29288 3692 31392 3720
rect 29288 3652 29316 3692
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 32490 3720 32496 3732
rect 31496 3692 32496 3720
rect 22695 3624 24256 3652
rect 22695 3621 22707 3624
rect 22649 3615 22707 3621
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3553 15163 3587
rect 15105 3547 15163 3553
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 17678 3584 17684 3596
rect 15252 3556 17684 3584
rect 15252 3544 15258 3556
rect 17678 3544 17684 3556
rect 17736 3584 17742 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17736 3556 18061 3584
rect 17736 3544 17742 3556
rect 18049 3553 18061 3556
rect 18095 3584 18107 3587
rect 20530 3584 20536 3596
rect 18095 3556 20536 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 20530 3544 20536 3556
rect 20588 3544 20594 3596
rect 20806 3544 20812 3596
rect 20864 3544 20870 3596
rect 21634 3544 21640 3596
rect 21692 3584 21698 3596
rect 23753 3587 23811 3593
rect 23753 3584 23765 3587
rect 21692 3556 23765 3584
rect 21692 3544 21698 3556
rect 23753 3553 23765 3556
rect 23799 3553 23811 3587
rect 23753 3547 23811 3553
rect 23842 3544 23848 3596
rect 23900 3584 23906 3596
rect 24029 3587 24087 3593
rect 24029 3584 24041 3587
rect 23900 3556 24041 3584
rect 23900 3544 23906 3556
rect 24029 3553 24041 3556
rect 24075 3584 24087 3587
rect 24118 3584 24124 3596
rect 24075 3556 24124 3584
rect 24075 3553 24087 3556
rect 24029 3547 24087 3553
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 24228 3584 24256 3624
rect 25976 3624 26924 3652
rect 28092 3624 29316 3652
rect 29733 3655 29791 3661
rect 24581 3587 24639 3593
rect 24228 3556 24532 3584
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 14292 3488 14841 3516
rect 10505 3479 10563 3485
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 20824 3516 20852 3544
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20824 3488 20913 3516
rect 14829 3479 14887 3485
rect 20901 3485 20913 3488
rect 20947 3485 20959 3519
rect 24394 3516 24400 3528
rect 22310 3488 24400 3516
rect 20901 3479 20959 3485
rect 10520 3448 10548 3479
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 10520 3420 12434 3448
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 12406 3380 12434 3420
rect 14182 3408 14188 3460
rect 14240 3448 14246 3460
rect 14240 3420 18184 3448
rect 14240 3408 14246 3420
rect 17954 3380 17960 3392
rect 12406 3352 17960 3380
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18156 3380 18184 3420
rect 20714 3408 20720 3460
rect 20772 3448 20778 3460
rect 21177 3451 21235 3457
rect 21177 3448 21189 3451
rect 20772 3420 21189 3448
rect 20772 3408 20778 3420
rect 21177 3417 21189 3420
rect 21223 3417 21235 3451
rect 24504 3448 24532 3556
rect 24581 3553 24593 3587
rect 24627 3584 24639 3587
rect 24854 3584 24860 3596
rect 24627 3556 24860 3584
rect 24627 3553 24639 3556
rect 24581 3547 24639 3553
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 25976 3502 26004 3624
rect 26050 3544 26056 3596
rect 26108 3584 26114 3596
rect 26786 3584 26792 3596
rect 26108 3556 26792 3584
rect 26108 3544 26114 3556
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 26896 3584 26924 3624
rect 29733 3621 29745 3655
rect 29779 3652 29791 3655
rect 30098 3652 30104 3664
rect 29779 3624 30104 3652
rect 29779 3621 29791 3624
rect 29733 3615 29791 3621
rect 30098 3612 30104 3624
rect 30156 3612 30162 3664
rect 31496 3652 31524 3692
rect 32490 3680 32496 3692
rect 32548 3680 32554 3732
rect 32674 3720 32680 3732
rect 32635 3692 32680 3720
rect 32674 3680 32680 3692
rect 32732 3680 32738 3732
rect 34698 3680 34704 3732
rect 34756 3720 34762 3732
rect 34885 3723 34943 3729
rect 34885 3720 34897 3723
rect 34756 3692 34897 3720
rect 34756 3680 34762 3692
rect 34885 3689 34897 3692
rect 34931 3689 34943 3723
rect 34885 3683 34943 3689
rect 31404 3624 31524 3652
rect 31404 3584 31432 3624
rect 31570 3612 31576 3664
rect 31628 3652 31634 3664
rect 33321 3655 33379 3661
rect 33321 3652 33333 3655
rect 31628 3624 33333 3652
rect 31628 3612 31634 3624
rect 33321 3621 33333 3624
rect 33367 3621 33379 3655
rect 33321 3615 33379 3621
rect 35342 3612 35348 3664
rect 35400 3652 35406 3664
rect 36081 3655 36139 3661
rect 36081 3652 36093 3655
rect 35400 3624 36093 3652
rect 35400 3612 35406 3624
rect 36081 3621 36093 3624
rect 36127 3621 36139 3655
rect 36081 3615 36139 3621
rect 26896 3556 31432 3584
rect 31481 3587 31539 3593
rect 31481 3553 31493 3587
rect 31527 3584 31539 3587
rect 32030 3584 32036 3596
rect 31527 3556 32036 3584
rect 31527 3553 31539 3556
rect 31481 3547 31539 3553
rect 32030 3544 32036 3556
rect 32088 3544 32094 3596
rect 33502 3584 33508 3596
rect 33244 3556 33508 3584
rect 33244 3528 33272 3556
rect 33502 3544 33508 3556
rect 33560 3584 33566 3596
rect 35434 3584 35440 3596
rect 33560 3556 35440 3584
rect 33560 3544 33566 3556
rect 28442 3476 28448 3528
rect 28500 3516 28506 3528
rect 29914 3516 29920 3528
rect 28500 3488 29920 3516
rect 28500 3476 28506 3488
rect 29914 3476 29920 3488
rect 29972 3476 29978 3528
rect 31754 3476 31760 3528
rect 31812 3516 31818 3528
rect 32125 3519 32183 3525
rect 32125 3516 32137 3519
rect 31812 3488 32137 3516
rect 31812 3476 31818 3488
rect 32125 3485 32137 3488
rect 32171 3516 32183 3519
rect 32769 3519 32827 3525
rect 32769 3516 32781 3519
rect 32171 3488 32781 3516
rect 32171 3485 32183 3488
rect 32125 3479 32183 3485
rect 32769 3485 32781 3488
rect 32815 3516 32827 3519
rect 33226 3516 33232 3528
rect 32815 3488 33232 3516
rect 32815 3485 32827 3488
rect 32769 3479 32827 3485
rect 33226 3476 33232 3488
rect 33284 3476 33290 3528
rect 33318 3476 33324 3528
rect 33376 3516 33382 3528
rect 34072 3525 34100 3556
rect 35434 3544 35440 3556
rect 35492 3544 35498 3596
rect 33413 3519 33471 3525
rect 33413 3516 33425 3519
rect 33376 3488 33425 3516
rect 33376 3476 33382 3488
rect 33413 3485 33425 3488
rect 33459 3485 33471 3519
rect 33413 3479 33471 3485
rect 34057 3519 34115 3525
rect 34057 3485 34069 3519
rect 34103 3485 34115 3519
rect 34057 3479 34115 3485
rect 36170 3476 36176 3528
rect 36228 3516 36234 3528
rect 36265 3519 36323 3525
rect 36265 3516 36277 3519
rect 36228 3488 36277 3516
rect 36228 3476 36234 3488
rect 36265 3485 36277 3488
rect 36311 3485 36323 3519
rect 36265 3479 36323 3485
rect 24857 3451 24915 3457
rect 24857 3448 24869 3451
rect 24504 3420 24869 3448
rect 21177 3411 21235 3417
rect 24857 3417 24869 3420
rect 24903 3417 24915 3451
rect 27062 3448 27068 3460
rect 27023 3420 27068 3448
rect 24857 3411 24915 3417
rect 27062 3408 27068 3420
rect 27120 3408 27126 3460
rect 30926 3448 30932 3460
rect 28290 3420 29868 3448
rect 30774 3420 30932 3448
rect 26142 3380 26148 3392
rect 18156 3352 26148 3380
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 26329 3383 26387 3389
rect 26329 3380 26341 3383
rect 26292 3352 26341 3380
rect 26292 3340 26298 3352
rect 26329 3349 26341 3352
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 26418 3340 26424 3392
rect 26476 3380 26482 3392
rect 27706 3380 27712 3392
rect 26476 3352 27712 3380
rect 26476 3340 26482 3352
rect 27706 3340 27712 3352
rect 27764 3340 27770 3392
rect 28534 3380 28540 3392
rect 28495 3352 28540 3380
rect 28534 3340 28540 3352
rect 28592 3380 28598 3392
rect 28902 3380 28908 3392
rect 28592 3352 28908 3380
rect 28592 3340 28598 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 29840 3380 29868 3420
rect 30926 3408 30932 3420
rect 30984 3408 30990 3460
rect 31110 3408 31116 3460
rect 31168 3448 31174 3460
rect 31205 3451 31263 3457
rect 31205 3448 31217 3451
rect 31168 3420 31217 3448
rect 31168 3408 31174 3420
rect 31205 3417 31217 3420
rect 31251 3417 31263 3451
rect 33965 3451 34023 3457
rect 33965 3448 33977 3451
rect 31205 3411 31263 3417
rect 31726 3420 33977 3448
rect 31726 3380 31754 3420
rect 33965 3417 33977 3420
rect 34011 3417 34023 3451
rect 33965 3411 34023 3417
rect 32030 3380 32036 3392
rect 29840 3352 31754 3380
rect 31991 3352 32036 3380
rect 32030 3340 32036 3352
rect 32088 3340 32094 3392
rect 35529 3383 35587 3389
rect 35529 3349 35541 3383
rect 35575 3380 35587 3383
rect 35986 3380 35992 3392
rect 35575 3352 35992 3380
rect 35575 3349 35587 3352
rect 35529 3343 35587 3349
rect 35986 3340 35992 3352
rect 36044 3340 36050 3392
rect 1104 3290 36892 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 36892 3290
rect 1104 3216 36892 3238
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 6886 3148 12541 3176
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 6886 3040 6914 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 12529 3139 12587 3145
rect 13265 3179 13323 3185
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 15194 3176 15200 3188
rect 13311 3148 15200 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 1903 3012 6914 3040
rect 11885 3043 11943 3049
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 13280 3040 13308 3139
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16942 3176 16948 3188
rect 16855 3148 16948 3176
rect 16942 3136 16948 3148
rect 17000 3176 17006 3188
rect 17770 3176 17776 3188
rect 17000 3148 17776 3176
rect 17000 3136 17006 3148
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 19705 3179 19763 3185
rect 19705 3145 19717 3179
rect 19751 3176 19763 3179
rect 23566 3176 23572 3188
rect 19751 3148 23572 3176
rect 19751 3145 19763 3148
rect 19705 3139 19763 3145
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 24854 3176 24860 3188
rect 23952 3148 24860 3176
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15344 3080 20010 3108
rect 15344 3068 15350 3080
rect 20898 3068 20904 3120
rect 20956 3108 20962 3120
rect 22005 3111 22063 3117
rect 22005 3108 22017 3111
rect 20956 3080 22017 3108
rect 20956 3068 20962 3080
rect 12759 3012 13308 3040
rect 14277 3043 14335 3049
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 14277 3009 14289 3043
rect 14323 3040 14335 3043
rect 14826 3040 14832 3052
rect 14323 3012 14832 3040
rect 14323 3009 14335 3012
rect 14277 3003 14335 3009
rect 11900 2972 11928 3003
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16942 3040 16948 3052
rect 16163 3012 16948 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 21468 3049 21496 3080
rect 22005 3077 22017 3080
rect 22051 3108 22063 3111
rect 23952 3108 23980 3148
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 26142 3136 26148 3188
rect 26200 3176 26206 3188
rect 31570 3176 31576 3188
rect 26200 3148 31576 3176
rect 26200 3136 26206 3148
rect 31570 3136 31576 3148
rect 31628 3136 31634 3188
rect 31662 3136 31668 3188
rect 31720 3176 31726 3188
rect 32030 3176 32036 3188
rect 31720 3148 32036 3176
rect 31720 3136 31726 3148
rect 32030 3136 32036 3148
rect 32088 3136 32094 3188
rect 32490 3136 32496 3188
rect 32548 3176 32554 3188
rect 33137 3179 33195 3185
rect 33137 3176 33149 3179
rect 32548 3148 33149 3176
rect 32548 3136 32554 3148
rect 33137 3145 33149 3148
rect 33183 3145 33195 3179
rect 33137 3139 33195 3145
rect 25866 3108 25872 3120
rect 22051 3080 23980 3108
rect 25827 3080 25872 3108
rect 22051 3077 22063 3080
rect 22005 3071 22063 3077
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 22925 3043 22983 3049
rect 22925 3009 22937 3043
rect 22971 3040 22983 3043
rect 23106 3040 23112 3052
rect 22971 3012 23112 3040
rect 22971 3009 22983 3012
rect 22925 3003 22983 3009
rect 23106 3000 23112 3012
rect 23164 3000 23170 3052
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 23860 3049 23888 3080
rect 25866 3068 25872 3080
rect 25924 3068 25930 3120
rect 26418 3108 26424 3120
rect 26379 3080 26424 3108
rect 26418 3068 26424 3080
rect 26476 3068 26482 3120
rect 26605 3111 26663 3117
rect 26605 3077 26617 3111
rect 26651 3108 26663 3111
rect 26694 3108 26700 3120
rect 26651 3080 26700 3108
rect 26651 3077 26663 3080
rect 26605 3071 26663 3077
rect 26694 3068 26700 3080
rect 26752 3068 26758 3120
rect 29730 3108 29736 3120
rect 28198 3080 29736 3108
rect 29730 3068 29736 3080
rect 29788 3068 29794 3120
rect 33686 3108 33692 3120
rect 30866 3080 33692 3108
rect 33686 3068 33692 3080
rect 33744 3068 33750 3120
rect 34790 3068 34796 3120
rect 34848 3108 34854 3120
rect 34977 3111 35035 3117
rect 34977 3108 34989 3111
rect 34848 3080 34989 3108
rect 34848 3068 34854 3080
rect 34977 3077 34989 3080
rect 35023 3108 35035 3111
rect 35342 3108 35348 3120
rect 35023 3080 35348 3108
rect 35023 3077 35035 3080
rect 34977 3071 35035 3077
rect 35342 3068 35348 3080
rect 35400 3068 35406 3120
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23808 3012 23857 3040
rect 23808 3000 23814 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 28905 3043 28963 3049
rect 23845 3003 23903 3009
rect 19058 2972 19064 2984
rect 11900 2944 19064 2972
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 21174 2972 21180 2984
rect 21135 2944 21180 2972
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 21376 2944 24133 2972
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 15933 2907 15991 2913
rect 15933 2904 15945 2907
rect 12492 2876 15945 2904
rect 12492 2864 12498 2876
rect 15933 2873 15945 2876
rect 15979 2873 15991 2907
rect 15933 2867 15991 2873
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 4672 2808 11713 2836
rect 4672 2796 4678 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 14090 2836 14096 2848
rect 14051 2808 14096 2836
rect 11701 2799 11759 2805
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 21376 2836 21404 2944
rect 24121 2941 24133 2944
rect 24167 2972 24179 2975
rect 25240 2972 25268 3026
rect 28905 3009 28917 3043
rect 28951 3040 28963 3043
rect 29178 3040 29184 3052
rect 28951 3012 29184 3040
rect 28951 3009 28963 3012
rect 28905 3003 28963 3009
rect 29178 3000 29184 3012
rect 29236 3040 29242 3052
rect 29362 3040 29368 3052
rect 29236 3012 29368 3040
rect 29236 3000 29242 3012
rect 29362 3000 29368 3012
rect 29420 3000 29426 3052
rect 31478 3000 31484 3052
rect 31536 3040 31542 3052
rect 31665 3043 31723 3049
rect 31665 3040 31677 3043
rect 31536 3012 31677 3040
rect 31536 3000 31542 3012
rect 31665 3009 31677 3012
rect 31711 3009 31723 3043
rect 31665 3003 31723 3009
rect 31754 3000 31760 3052
rect 31812 3040 31818 3052
rect 32306 3040 32312 3052
rect 31812 3012 31857 3040
rect 32267 3012 32312 3040
rect 31812 3000 31818 3012
rect 32306 3000 32312 3012
rect 32364 3000 32370 3052
rect 33226 3040 33232 3052
rect 33187 3012 33232 3040
rect 33226 3000 33232 3012
rect 33284 3040 33290 3052
rect 33873 3043 33931 3049
rect 33873 3040 33885 3043
rect 33284 3012 33885 3040
rect 33284 3000 33290 3012
rect 33873 3009 33885 3012
rect 33919 3009 33931 3043
rect 36078 3040 36084 3052
rect 36039 3012 36084 3040
rect 33873 3003 33931 3009
rect 36078 3000 36084 3012
rect 36136 3000 36142 3052
rect 28629 2975 28687 2981
rect 24167 2944 25176 2972
rect 25240 2944 27568 2972
rect 24167 2941 24179 2944
rect 24121 2935 24179 2941
rect 25148 2904 25176 2944
rect 27157 2907 27215 2913
rect 27157 2904 27169 2907
rect 25148 2876 27169 2904
rect 27157 2873 27169 2876
rect 27203 2873 27215 2907
rect 27157 2867 27215 2873
rect 19300 2808 21404 2836
rect 19300 2796 19306 2808
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 22612 2808 22753 2836
rect 22612 2796 22618 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 27540 2836 27568 2944
rect 28629 2941 28641 2975
rect 28675 2972 28687 2975
rect 28675 2944 28856 2972
rect 28675 2941 28687 2944
rect 28629 2935 28687 2941
rect 28828 2904 28856 2944
rect 28994 2932 29000 2984
rect 29052 2972 29058 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 29052 2944 29653 2972
rect 29052 2932 29058 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 29730 2932 29736 2984
rect 29788 2972 29794 2984
rect 33781 2975 33839 2981
rect 33781 2972 33793 2975
rect 29788 2944 33793 2972
rect 29788 2932 29794 2944
rect 33781 2941 33793 2944
rect 33827 2941 33839 2975
rect 36354 2972 36360 2984
rect 36315 2944 36360 2972
rect 33781 2935 33839 2941
rect 36354 2932 36360 2944
rect 36412 2932 36418 2984
rect 28902 2904 28908 2916
rect 28828 2876 28908 2904
rect 28902 2864 28908 2876
rect 28960 2864 28966 2916
rect 32493 2907 32551 2913
rect 32493 2904 32505 2907
rect 30668 2876 32505 2904
rect 29086 2836 29092 2848
rect 27540 2808 29092 2836
rect 22741 2799 22799 2805
rect 29086 2796 29092 2808
rect 29144 2796 29150 2848
rect 29638 2796 29644 2848
rect 29696 2836 29702 2848
rect 30668 2836 30696 2876
rect 32493 2873 32505 2876
rect 32539 2873 32551 2907
rect 34790 2904 34796 2916
rect 34751 2876 34796 2904
rect 32493 2867 32551 2873
rect 34790 2864 34796 2876
rect 34848 2864 34854 2916
rect 31110 2836 31116 2848
rect 29696 2808 30696 2836
rect 31071 2808 31116 2836
rect 29696 2796 29702 2808
rect 31110 2796 31116 2808
rect 31168 2796 31174 2848
rect 1104 2746 36892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36892 2746
rect 1104 2672 36892 2694
rect 1946 2592 1952 2644
rect 2004 2632 2010 2644
rect 2501 2635 2559 2641
rect 2501 2632 2513 2635
rect 2004 2604 2513 2632
rect 2004 2592 2010 2604
rect 2501 2601 2513 2604
rect 2547 2601 2559 2635
rect 4706 2632 4712 2644
rect 4667 2604 4712 2632
rect 2501 2595 2559 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 19429 2635 19487 2641
rect 19429 2632 19441 2635
rect 19116 2604 19441 2632
rect 19116 2592 19122 2604
rect 19429 2601 19441 2604
rect 19475 2601 19487 2635
rect 19429 2595 19487 2601
rect 21266 2592 21272 2644
rect 21324 2632 21330 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21324 2604 22017 2632
rect 21324 2592 21330 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 25958 2592 25964 2644
rect 26016 2632 26022 2644
rect 26786 2632 26792 2644
rect 26016 2604 26792 2632
rect 26016 2592 26022 2604
rect 26786 2592 26792 2604
rect 26844 2592 26850 2644
rect 28350 2632 28356 2644
rect 27448 2604 28356 2632
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 13262 2564 13268 2576
rect 9447 2536 13268 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 16942 2524 16948 2576
rect 17000 2564 17006 2576
rect 27448 2564 27476 2604
rect 28350 2592 28356 2604
rect 28408 2592 28414 2644
rect 29089 2635 29147 2641
rect 29089 2601 29101 2635
rect 29135 2632 29147 2635
rect 29270 2632 29276 2644
rect 29135 2604 29276 2632
rect 29135 2601 29147 2604
rect 29089 2595 29147 2601
rect 29270 2592 29276 2604
rect 29328 2592 29334 2644
rect 29546 2592 29552 2644
rect 29604 2632 29610 2644
rect 31481 2635 31539 2641
rect 31481 2632 31493 2635
rect 29604 2604 31493 2632
rect 29604 2592 29610 2604
rect 31481 2601 31493 2604
rect 31527 2601 31539 2635
rect 31481 2595 31539 2601
rect 33689 2635 33747 2641
rect 33689 2601 33701 2635
rect 33735 2632 33747 2635
rect 34606 2632 34612 2644
rect 33735 2604 34612 2632
rect 33735 2601 33747 2604
rect 33689 2595 33747 2601
rect 34606 2592 34612 2604
rect 34664 2592 34670 2644
rect 35986 2592 35992 2644
rect 36044 2632 36050 2644
rect 36173 2635 36231 2641
rect 36173 2632 36185 2635
rect 36044 2604 36185 2632
rect 36044 2592 36050 2604
rect 36173 2601 36185 2604
rect 36219 2601 36231 2635
rect 36173 2595 36231 2601
rect 17000 2536 22094 2564
rect 17000 2524 17006 2536
rect 4614 2496 4620 2508
rect 1872 2468 4620 2496
rect 1872 2437 1900 2468
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 14090 2496 14096 2508
rect 10520 2468 14096 2496
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4706 2428 4712 2440
rect 4295 2400 4712 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 2332 2360 2360 2391
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 5534 2428 5540 2440
rect 5495 2400 5540 2428
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 10520 2428 10548 2468
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 17678 2496 17684 2508
rect 14568 2468 17684 2496
rect 6871 2400 10548 2428
rect 11977 2431 12035 2437
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12434 2428 12440 2440
rect 12023 2400 12440 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 14568 2437 14596 2468
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 17402 2428 17408 2440
rect 15887 2400 17408 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 17819 2400 18368 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 2961 2363 3019 2369
rect 2961 2360 2973 2363
rect 72 2332 2973 2360
rect 72 2320 78 2332
rect 2961 2329 2973 2332
rect 3007 2329 3019 2363
rect 2961 2323 3019 2329
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 9953 2363 10011 2369
rect 9953 2329 9965 2363
rect 9999 2360 10011 2363
rect 10318 2360 10324 2372
rect 9999 2332 10324 2360
rect 9999 2329 10011 2332
rect 9953 2323 10011 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3292 2264 4077 2292
rect 3292 2252 3298 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5224 2264 5365 2292
rect 5224 2252 5230 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2292 8539 2295
rect 9232 2292 9260 2323
rect 10318 2320 10324 2332
rect 10376 2360 10382 2372
rect 10505 2363 10563 2369
rect 10505 2360 10517 2363
rect 10376 2332 10517 2360
rect 10376 2320 10382 2332
rect 10505 2329 10517 2332
rect 10551 2329 10563 2363
rect 10505 2323 10563 2329
rect 18340 2304 18368 2400
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 18748 2400 19625 2428
rect 18748 2388 18754 2400
rect 19613 2397 19625 2400
rect 19659 2428 19671 2431
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19659 2400 20085 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20990 2428 20996 2440
rect 20951 2400 20996 2428
rect 20073 2391 20131 2397
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 10594 2292 10600 2304
rect 8527 2264 9260 2292
rect 10555 2264 10600 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 13596 2264 14381 2292
rect 13596 2252 13602 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15528 2264 15669 2292
rect 15528 2252 15534 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17460 2264 17601 2292
rect 17460 2252 17466 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 17589 2255 17647 2261
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20680 2264 20821 2292
rect 20680 2252 20686 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 22066 2292 22094 2536
rect 26252 2536 27476 2564
rect 22278 2456 22284 2508
rect 22336 2456 22342 2508
rect 23750 2496 23756 2508
rect 23711 2468 23756 2496
rect 23750 2456 23756 2468
rect 23808 2496 23814 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23808 2468 24593 2496
rect 23808 2456 23814 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24854 2496 24860 2508
rect 24815 2468 24860 2496
rect 24581 2459 24639 2465
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 24946 2456 24952 2508
rect 25004 2496 25010 2508
rect 26252 2496 26280 2536
rect 28626 2524 28632 2576
rect 28684 2564 28690 2576
rect 32766 2564 32772 2576
rect 28684 2536 29868 2564
rect 28684 2524 28690 2536
rect 25004 2468 26280 2496
rect 25004 2456 25010 2468
rect 26326 2456 26332 2508
rect 26384 2496 26390 2508
rect 26384 2468 26429 2496
rect 26384 2456 26390 2468
rect 26786 2456 26792 2508
rect 26844 2496 26850 2508
rect 27341 2499 27399 2505
rect 27341 2496 27353 2499
rect 26844 2468 27353 2496
rect 26844 2456 26850 2468
rect 27341 2465 27353 2468
rect 27387 2465 27399 2499
rect 27341 2459 27399 2465
rect 27617 2499 27675 2505
rect 27617 2465 27629 2499
rect 27663 2496 27675 2499
rect 27663 2468 29408 2496
rect 27663 2465 27675 2468
rect 27617 2459 27675 2465
rect 22296 2428 22324 2456
rect 29380 2428 29408 2468
rect 29454 2456 29460 2508
rect 29512 2496 29518 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29512 2468 29745 2496
rect 29512 2456 29518 2468
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 29840 2496 29868 2536
rect 31128 2536 32772 2564
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 29840 2468 30021 2496
rect 29733 2459 29791 2465
rect 30009 2465 30021 2468
rect 30055 2465 30067 2499
rect 30009 2459 30067 2465
rect 29546 2428 29552 2440
rect 22296 2400 22402 2428
rect 29380 2400 29552 2428
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 31128 2414 31156 2536
rect 32766 2524 32772 2536
rect 32824 2524 32830 2576
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 31312 2468 35173 2496
rect 23477 2363 23535 2369
rect 23477 2329 23489 2363
rect 23523 2360 23535 2363
rect 24946 2360 24952 2372
rect 23523 2332 24952 2360
rect 23523 2329 23535 2332
rect 23477 2323 23535 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 25866 2320 25872 2372
rect 25924 2320 25930 2372
rect 29914 2360 29920 2372
rect 26160 2332 26556 2360
rect 28842 2332 29920 2360
rect 26160 2292 26188 2332
rect 22066 2264 26188 2292
rect 26528 2292 26556 2332
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 31312 2292 31340 2468
rect 35161 2465 35173 2468
rect 35207 2465 35219 2499
rect 35161 2459 35219 2465
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 32122 2428 32128 2440
rect 31444 2400 32128 2428
rect 31444 2388 31450 2400
rect 32122 2388 32128 2400
rect 32180 2428 32186 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32180 2400 32321 2428
rect 32180 2388 32186 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32585 2431 32643 2437
rect 32585 2397 32597 2431
rect 32631 2397 32643 2431
rect 32585 2391 32643 2397
rect 31478 2320 31484 2372
rect 31536 2360 31542 2372
rect 32600 2360 32628 2391
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 32916 2400 33793 2428
rect 32916 2388 32922 2400
rect 33781 2397 33793 2400
rect 33827 2428 33839 2431
rect 34238 2428 34244 2440
rect 33827 2400 34244 2428
rect 33827 2397 33839 2400
rect 33781 2391 33839 2397
rect 34238 2388 34244 2400
rect 34296 2388 34302 2440
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2428 34943 2431
rect 35618 2428 35624 2440
rect 34931 2400 35624 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 35618 2388 35624 2400
rect 35676 2388 35682 2440
rect 31536 2332 32628 2360
rect 31536 2320 31542 2332
rect 26528 2264 31340 2292
rect 20809 2255 20867 2261
rect 1104 2202 36892 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 36892 2202
rect 1104 2128 36892 2150
rect 18322 2048 18328 2100
rect 18380 2088 18386 2100
rect 25590 2088 25596 2100
rect 18380 2060 25596 2088
rect 18380 2048 18386 2060
rect 25590 2048 25596 2060
rect 25648 2048 25654 2100
rect 31478 2088 31484 2100
rect 28966 2060 31484 2088
rect 20530 1980 20536 2032
rect 20588 2020 20594 2032
rect 28966 2020 28994 2060
rect 31478 2048 31484 2060
rect 31536 2048 31542 2100
rect 20588 1992 28994 2020
rect 20588 1980 20594 1992
rect 29914 1980 29920 2032
rect 29972 2020 29978 2032
rect 33134 2020 33140 2032
rect 29972 1992 33140 2020
rect 29972 1980 29978 1992
rect 33134 1980 33140 1992
rect 33192 1980 33198 2032
rect 10594 1912 10600 1964
rect 10652 1952 10658 1964
rect 25038 1952 25044 1964
rect 10652 1924 25044 1952
rect 10652 1912 10658 1924
rect 25038 1912 25044 1924
rect 25096 1912 25102 1964
rect 25866 1912 25872 1964
rect 25924 1952 25930 1964
rect 33870 1952 33876 1964
rect 25924 1924 33876 1952
rect 25924 1912 25930 1924
rect 33870 1912 33876 1924
rect 33928 1912 33934 1964
rect 28350 1844 28356 1896
rect 28408 1884 28414 1896
rect 31202 1884 31208 1896
rect 28408 1856 31208 1884
rect 28408 1844 28414 1856
rect 31202 1844 31208 1856
rect 31260 1844 31266 1896
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20 37408 72 37460
rect 13544 37408 13596 37460
rect 16120 37408 16172 37460
rect 21272 37408 21324 37460
rect 5540 37315 5592 37324
rect 5540 37281 5549 37315
rect 5549 37281 5583 37315
rect 5583 37281 5592 37315
rect 5540 37272 5592 37281
rect 7104 37272 7156 37324
rect 10324 37272 10376 37324
rect 16120 37272 16172 37324
rect 1952 37204 2004 37256
rect 3056 37247 3108 37256
rect 3056 37213 3065 37247
rect 3065 37213 3099 37247
rect 3099 37213 3108 37247
rect 3056 37204 3108 37213
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 5172 37204 5224 37256
rect 7472 37247 7524 37256
rect 7472 37213 7481 37247
rect 7481 37213 7515 37247
rect 7515 37213 7524 37247
rect 7472 37204 7524 37213
rect 9036 37204 9088 37256
rect 10876 37247 10928 37256
rect 10876 37213 10885 37247
rect 10885 37213 10919 37247
rect 10919 37213 10928 37247
rect 10876 37204 10928 37213
rect 12440 37204 12492 37256
rect 14188 37204 14240 37256
rect 17040 37272 17092 37324
rect 17408 37204 17460 37256
rect 18880 37204 18932 37256
rect 8944 37136 8996 37188
rect 25504 37340 25556 37392
rect 22652 37272 22704 37324
rect 22560 37204 22612 37256
rect 24860 37315 24912 37324
rect 24860 37281 24869 37315
rect 24869 37281 24903 37315
rect 24903 37281 24912 37315
rect 24860 37272 24912 37281
rect 35532 37315 35584 37324
rect 35532 37281 35541 37315
rect 35541 37281 35575 37315
rect 35575 37281 35584 37315
rect 35532 37272 35584 37281
rect 24492 37204 24544 37256
rect 26792 37204 26844 37256
rect 28816 37204 28868 37256
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 3884 37068 3936 37120
rect 23204 37136 23256 37188
rect 28632 37136 28684 37188
rect 33600 37204 33652 37256
rect 35808 37247 35860 37256
rect 35808 37213 35817 37247
rect 35817 37213 35851 37247
rect 35851 37213 35860 37247
rect 35808 37204 35860 37213
rect 14464 37111 14516 37120
rect 14464 37077 14473 37111
rect 14473 37077 14507 37111
rect 14507 37077 14516 37111
rect 14464 37068 14516 37077
rect 19248 37068 19300 37120
rect 19340 37068 19392 37120
rect 26424 37068 26476 37120
rect 28356 37068 28408 37120
rect 29644 37068 29696 37120
rect 31760 37068 31812 37120
rect 33508 37068 33560 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1676 36907 1728 36916
rect 1676 36873 1685 36907
rect 1685 36873 1719 36907
rect 1719 36873 1728 36907
rect 1676 36864 1728 36873
rect 1952 36864 2004 36916
rect 3056 36864 3108 36916
rect 18880 36907 18932 36916
rect 18880 36873 18889 36907
rect 18889 36873 18923 36907
rect 18923 36873 18932 36907
rect 18880 36864 18932 36873
rect 24492 36907 24544 36916
rect 24492 36873 24501 36907
rect 24501 36873 24535 36907
rect 24535 36873 24544 36907
rect 24492 36864 24544 36873
rect 34796 36864 34848 36916
rect 36268 36907 36320 36916
rect 36268 36873 36277 36907
rect 36277 36873 36311 36907
rect 36311 36873 36320 36907
rect 36268 36864 36320 36873
rect 10876 36796 10928 36848
rect 1768 36728 1820 36780
rect 7472 36728 7524 36780
rect 11060 36728 11112 36780
rect 17592 36771 17644 36780
rect 17592 36737 17601 36771
rect 17601 36737 17635 36771
rect 17635 36737 17644 36771
rect 17592 36728 17644 36737
rect 19248 36796 19300 36848
rect 19432 36728 19484 36780
rect 23204 36771 23256 36780
rect 23204 36737 23213 36771
rect 23213 36737 23247 36771
rect 23247 36737 23256 36771
rect 23204 36728 23256 36737
rect 23388 36728 23440 36780
rect 35992 36728 36044 36780
rect 29736 36592 29788 36644
rect 28632 36524 28684 36576
rect 28816 36567 28868 36576
rect 28816 36533 28825 36567
rect 28825 36533 28859 36567
rect 28859 36533 28868 36567
rect 28816 36524 28868 36533
rect 33600 36524 33652 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2780 36320 2832 36372
rect 36728 36320 36780 36372
rect 32312 36116 32364 36168
rect 17592 36048 17644 36100
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 36084 35683 36136 35692
rect 36084 35649 36093 35683
rect 36093 35649 36127 35683
rect 36127 35649 36136 35683
rect 36084 35640 36136 35649
rect 36268 35479 36320 35488
rect 36268 35445 36277 35479
rect 36277 35445 36311 35479
rect 36311 35445 36320 35479
rect 36268 35436 36320 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 36084 35232 36136 35284
rect 2688 35028 2740 35080
rect 1676 34935 1728 34944
rect 1676 34901 1685 34935
rect 1685 34901 1719 34935
rect 1719 34901 1728 34935
rect 1676 34892 1728 34901
rect 35440 34935 35492 34944
rect 35440 34901 35449 34935
rect 35449 34901 35483 34935
rect 35483 34901 35492 34935
rect 35440 34892 35492 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 35532 33464 35584 33516
rect 36268 33371 36320 33380
rect 36268 33337 36277 33371
rect 36277 33337 36311 33371
rect 36311 33337 36320 33371
rect 36268 33328 36320 33337
rect 35532 33303 35584 33312
rect 35532 33269 35541 33303
rect 35541 33269 35575 33303
rect 35575 33269 35584 33303
rect 35532 33260 35584 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1676 32827 1728 32836
rect 1676 32793 1685 32827
rect 1685 32793 1719 32827
rect 1719 32793 1728 32827
rect 1676 32784 1728 32793
rect 17868 32716 17920 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1676 32555 1728 32564
rect 1676 32521 1685 32555
rect 1685 32521 1719 32555
rect 1719 32521 1728 32555
rect 1676 32512 1728 32521
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3976 32011 4028 32020
rect 3976 31977 3985 32011
rect 3985 31977 4019 32011
rect 4019 31977 4028 32011
rect 3976 31968 4028 31977
rect 36452 31832 36504 31884
rect 1860 31807 1912 31816
rect 1860 31773 1869 31807
rect 1869 31773 1903 31807
rect 1903 31773 1912 31807
rect 1860 31764 1912 31773
rect 4620 31807 4672 31816
rect 4620 31773 4629 31807
rect 4629 31773 4663 31807
rect 4663 31773 4672 31807
rect 4620 31764 4672 31773
rect 36360 31807 36412 31816
rect 36360 31773 36369 31807
rect 36369 31773 36403 31807
rect 36403 31773 36412 31807
rect 36360 31764 36412 31773
rect 1676 31671 1728 31680
rect 1676 31637 1685 31671
rect 1685 31637 1719 31671
rect 1719 31637 1728 31671
rect 1676 31628 1728 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1860 31424 1912 31476
rect 23388 31424 23440 31476
rect 32312 31424 32364 31476
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 19432 31288 19484 31340
rect 36360 31399 36412 31408
rect 36360 31365 36369 31399
rect 36369 31365 36403 31399
rect 36403 31365 36412 31399
rect 36360 31356 36412 31365
rect 27436 31331 27488 31340
rect 27436 31297 27445 31331
rect 27445 31297 27479 31331
rect 27479 31297 27488 31331
rect 27436 31288 27488 31297
rect 19984 31084 20036 31136
rect 23020 31127 23072 31136
rect 23020 31093 23029 31127
rect 23029 31093 23063 31127
rect 23063 31093 23072 31127
rect 23020 31084 23072 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1768 30923 1820 30932
rect 1768 30889 1777 30923
rect 1777 30889 1811 30923
rect 1811 30889 1820 30923
rect 1768 30880 1820 30889
rect 1860 30676 1912 30728
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 35624 30200 35676 30252
rect 35624 30039 35676 30048
rect 35624 30005 35633 30039
rect 35633 30005 35667 30039
rect 35667 30005 35676 30039
rect 35624 29996 35676 30005
rect 36268 30039 36320 30048
rect 36268 30005 36277 30039
rect 36277 30005 36311 30039
rect 36311 30005 36320 30039
rect 36268 29996 36320 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2688 29792 2740 29844
rect 1952 29588 2004 29640
rect 6092 29631 6144 29640
rect 6092 29597 6101 29631
rect 6101 29597 6135 29631
rect 6135 29597 6144 29631
rect 6092 29588 6144 29597
rect 11060 29588 11112 29640
rect 1676 29495 1728 29504
rect 1676 29461 1685 29495
rect 1685 29461 1719 29495
rect 1719 29461 1728 29495
rect 1676 29452 1728 29461
rect 17224 29452 17276 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 36268 28067 36320 28076
rect 36268 28033 36277 28067
rect 36277 28033 36311 28067
rect 36311 28033 36320 28067
rect 36268 28024 36320 28033
rect 36176 27863 36228 27872
rect 36176 27829 36185 27863
rect 36185 27829 36219 27863
rect 36219 27829 36228 27863
rect 36176 27820 36228 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3700 27412 3752 27464
rect 1676 27319 1728 27328
rect 1676 27285 1685 27319
rect 1685 27285 1719 27319
rect 1719 27285 1728 27319
rect 1676 27276 1728 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 26792 26571 26844 26580
rect 26792 26537 26801 26571
rect 26801 26537 26835 26571
rect 26835 26537 26844 26571
rect 26792 26528 26844 26537
rect 35808 26460 35860 26512
rect 35348 26324 35400 26376
rect 27620 26256 27672 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 4620 24148 4672 24200
rect 30380 24148 30432 24200
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 8944 23808 8996 23860
rect 36360 23851 36412 23860
rect 36360 23817 36369 23851
rect 36369 23817 36403 23851
rect 36403 23817 36412 23851
rect 36360 23808 36412 23817
rect 12716 23672 12768 23724
rect 1952 23536 2004 23588
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 12716 23511 12768 23520
rect 12716 23477 12725 23511
rect 12725 23477 12759 23511
rect 12759 23477 12768 23511
rect 12716 23468 12768 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3700 23264 3752 23316
rect 13268 22924 13320 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 36084 22627 36136 22636
rect 36084 22593 36093 22627
rect 36093 22593 36127 22627
rect 36127 22593 36136 22627
rect 36084 22584 36136 22593
rect 36268 22491 36320 22500
rect 36268 22457 36277 22491
rect 36277 22457 36311 22491
rect 36311 22457 36320 22491
rect 36268 22448 36320 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 24584 21836 24636 21888
rect 27436 21836 27488 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2320 21292 2372 21344
rect 35716 21292 35768 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 35992 21088 36044 21140
rect 4620 20952 4672 21004
rect 1860 20884 1912 20936
rect 35716 20884 35768 20936
rect 17960 20816 18012 20868
rect 33140 20816 33192 20868
rect 9220 20791 9272 20800
rect 9220 20757 9229 20791
rect 9229 20757 9263 20791
rect 9263 20757 9272 20791
rect 9220 20748 9272 20757
rect 36268 20791 36320 20800
rect 36268 20757 36277 20791
rect 36277 20757 36311 20791
rect 36311 20757 36320 20791
rect 36268 20748 36320 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 35716 20247 35768 20256
rect 35716 20213 35725 20247
rect 35725 20213 35759 20247
rect 35759 20213 35768 20247
rect 35716 20204 35768 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 33140 20000 33192 20052
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 21364 19796 21416 19848
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 36084 19456 36136 19508
rect 34612 19320 34664 19372
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 35348 18912 35400 18964
rect 28540 18708 28592 18760
rect 34520 18708 34572 18760
rect 1584 18640 1636 18692
rect 2688 18640 2740 18692
rect 23572 18615 23624 18624
rect 23572 18581 23581 18615
rect 23581 18581 23615 18615
rect 23615 18581 23624 18615
rect 23572 18572 23624 18581
rect 36268 18615 36320 18624
rect 36268 18581 36277 18615
rect 36277 18581 36311 18615
rect 36311 18581 36320 18615
rect 36268 18572 36320 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 24584 18411 24636 18420
rect 24584 18377 24593 18411
rect 24593 18377 24627 18411
rect 24627 18377 24636 18411
rect 24584 18368 24636 18377
rect 30380 18232 30432 18284
rect 23112 18164 23164 18216
rect 25688 18096 25740 18148
rect 5540 18028 5592 18080
rect 22008 18028 22060 18080
rect 22836 18028 22888 18080
rect 23848 18028 23900 18080
rect 24768 18028 24820 18080
rect 26700 18028 26752 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 21364 17867 21416 17876
rect 21364 17833 21373 17867
rect 21373 17833 21407 17867
rect 21407 17833 21416 17867
rect 21364 17824 21416 17833
rect 34520 17824 34572 17876
rect 23204 17756 23256 17808
rect 23112 17731 23164 17740
rect 23112 17697 23121 17731
rect 23121 17697 23155 17731
rect 23155 17697 23164 17731
rect 23112 17688 23164 17697
rect 23848 17663 23900 17672
rect 23848 17629 23857 17663
rect 23857 17629 23891 17663
rect 23891 17629 23900 17663
rect 23848 17620 23900 17629
rect 24584 17620 24636 17672
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 29736 17620 29788 17672
rect 20904 17527 20956 17536
rect 20904 17493 20913 17527
rect 20913 17493 20947 17527
rect 20947 17493 20956 17527
rect 20904 17484 20956 17493
rect 27804 17552 27856 17604
rect 24584 17484 24636 17536
rect 25872 17484 25924 17536
rect 26148 17484 26200 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 24584 17255 24636 17264
rect 24584 17221 24593 17255
rect 24593 17221 24627 17255
rect 24627 17221 24636 17255
rect 24584 17212 24636 17221
rect 21364 17144 21416 17196
rect 22836 17187 22888 17196
rect 22836 17153 22845 17187
rect 22845 17153 22879 17187
rect 22879 17153 22888 17187
rect 22836 17144 22888 17153
rect 27436 17212 27488 17264
rect 25412 17144 25464 17196
rect 26148 17144 26200 17196
rect 36084 17187 36136 17196
rect 36084 17153 36093 17187
rect 36093 17153 36127 17187
rect 36127 17153 36136 17187
rect 36084 17144 36136 17153
rect 20904 17076 20956 17128
rect 21640 17076 21692 17128
rect 25780 17119 25832 17128
rect 23204 17008 23256 17060
rect 25780 17085 25789 17119
rect 25789 17085 25823 17119
rect 25823 17085 25832 17119
rect 25780 17076 25832 17085
rect 26240 17008 26292 17060
rect 20996 16940 21048 16992
rect 21364 16983 21416 16992
rect 21364 16949 21373 16983
rect 21373 16949 21407 16983
rect 21407 16949 21416 16983
rect 21364 16940 21416 16949
rect 35624 17076 35676 17128
rect 26424 17008 26476 17060
rect 35532 17008 35584 17060
rect 36268 17051 36320 17060
rect 36268 17017 36277 17051
rect 36277 17017 36311 17051
rect 36311 17017 36320 17051
rect 36268 17008 36320 17017
rect 26608 16940 26660 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 25412 16736 25464 16788
rect 27620 16736 27672 16788
rect 20720 16643 20772 16652
rect 11704 16532 11756 16584
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 21364 16600 21416 16652
rect 21824 16507 21876 16516
rect 21824 16473 21833 16507
rect 21833 16473 21867 16507
rect 21867 16473 21876 16507
rect 21824 16464 21876 16473
rect 22008 16532 22060 16584
rect 23572 16532 23624 16584
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 27528 16668 27580 16720
rect 26056 16600 26108 16652
rect 26700 16643 26752 16652
rect 26700 16609 26709 16643
rect 26709 16609 26743 16643
rect 26743 16609 26752 16643
rect 26700 16600 26752 16609
rect 29000 16600 29052 16652
rect 27436 16575 27488 16584
rect 27436 16541 27445 16575
rect 27445 16541 27479 16575
rect 27479 16541 27488 16575
rect 27436 16532 27488 16541
rect 22100 16464 22152 16516
rect 22652 16464 22704 16516
rect 26332 16464 26384 16516
rect 26608 16507 26660 16516
rect 26608 16473 26617 16507
rect 26617 16473 26651 16507
rect 26651 16473 26660 16507
rect 26608 16464 26660 16473
rect 27160 16464 27212 16516
rect 27804 16464 27856 16516
rect 28172 16464 28224 16516
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 20168 16439 20220 16448
rect 20168 16405 20177 16439
rect 20177 16405 20211 16439
rect 20211 16405 20220 16439
rect 20168 16396 20220 16405
rect 21916 16439 21968 16448
rect 21916 16405 21925 16439
rect 21925 16405 21959 16439
rect 21959 16405 21968 16439
rect 21916 16396 21968 16405
rect 23480 16396 23532 16448
rect 23848 16439 23900 16448
rect 23848 16405 23857 16439
rect 23857 16405 23891 16439
rect 23891 16405 23900 16439
rect 23848 16396 23900 16405
rect 24860 16396 24912 16448
rect 26148 16396 26200 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11704 16235 11756 16244
rect 11704 16201 11713 16235
rect 11713 16201 11747 16235
rect 11747 16201 11756 16235
rect 11704 16192 11756 16201
rect 17224 16192 17276 16244
rect 19340 16192 19392 16244
rect 22100 16192 22152 16244
rect 9220 16124 9272 16176
rect 22560 16167 22612 16176
rect 22560 16133 22569 16167
rect 22569 16133 22603 16167
rect 22603 16133 22612 16167
rect 22560 16124 22612 16133
rect 27344 16192 27396 16244
rect 25780 16124 25832 16176
rect 26792 16124 26844 16176
rect 20076 15988 20128 16040
rect 26148 16056 26200 16108
rect 26332 16056 26384 16108
rect 26608 16056 26660 16108
rect 20536 15988 20588 16040
rect 23848 15988 23900 16040
rect 24400 16031 24452 16040
rect 24400 15997 24409 16031
rect 24409 15997 24443 16031
rect 24443 15997 24452 16031
rect 24400 15988 24452 15997
rect 27620 16056 27672 16108
rect 22008 15920 22060 15972
rect 23296 15920 23348 15972
rect 23480 15920 23532 15972
rect 20812 15852 20864 15904
rect 21088 15852 21140 15904
rect 23664 15895 23716 15904
rect 23664 15861 23673 15895
rect 23673 15861 23707 15895
rect 23707 15861 23716 15895
rect 23664 15852 23716 15861
rect 26516 15852 26568 15904
rect 27252 15895 27304 15904
rect 27252 15861 27261 15895
rect 27261 15861 27295 15895
rect 27295 15861 27304 15895
rect 27252 15852 27304 15861
rect 27436 15852 27488 15904
rect 36360 15895 36412 15904
rect 36360 15861 36369 15895
rect 36369 15861 36403 15895
rect 36403 15861 36412 15895
rect 36360 15852 36412 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19340 15648 19392 15700
rect 21640 15648 21692 15700
rect 27988 15648 28040 15700
rect 33600 15691 33652 15700
rect 33600 15657 33609 15691
rect 33609 15657 33643 15691
rect 33643 15657 33652 15691
rect 33600 15648 33652 15657
rect 28080 15580 28132 15632
rect 19340 15512 19392 15564
rect 22100 15512 22152 15564
rect 23296 15512 23348 15564
rect 25228 15512 25280 15564
rect 27712 15555 27764 15564
rect 27712 15521 27721 15555
rect 27721 15521 27755 15555
rect 27755 15521 27764 15555
rect 27712 15512 27764 15521
rect 19064 15444 19116 15496
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 27612 15487 27664 15496
rect 27612 15453 27621 15487
rect 27621 15453 27655 15487
rect 27655 15453 27664 15487
rect 27612 15444 27664 15453
rect 33416 15487 33468 15496
rect 4712 15308 4764 15360
rect 20904 15419 20956 15428
rect 20904 15385 20913 15419
rect 20913 15385 20947 15419
rect 20947 15385 20956 15419
rect 20904 15376 20956 15385
rect 21732 15376 21784 15428
rect 22468 15419 22520 15428
rect 22468 15385 22477 15419
rect 22477 15385 22511 15419
rect 22511 15385 22520 15419
rect 22468 15376 22520 15385
rect 23572 15376 23624 15428
rect 24308 15376 24360 15428
rect 22192 15308 22244 15360
rect 26332 15376 26384 15428
rect 26516 15419 26568 15428
rect 26516 15385 26525 15419
rect 26525 15385 26559 15419
rect 26559 15385 26568 15419
rect 26516 15376 26568 15385
rect 26976 15376 27028 15428
rect 27896 15376 27948 15428
rect 27528 15308 27580 15360
rect 28264 15351 28316 15360
rect 28264 15317 28273 15351
rect 28273 15317 28307 15351
rect 28307 15317 28316 15351
rect 28264 15308 28316 15317
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 36360 15487 36412 15496
rect 36360 15453 36369 15487
rect 36369 15453 36403 15487
rect 36403 15453 36412 15487
rect 36360 15444 36412 15453
rect 35532 15308 35584 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 20536 15104 20588 15156
rect 22836 15104 22888 15156
rect 24952 15104 25004 15156
rect 26332 15104 26384 15156
rect 27528 15104 27580 15156
rect 36084 15147 36136 15156
rect 36084 15113 36093 15147
rect 36093 15113 36127 15147
rect 36127 15113 36136 15147
rect 36084 15104 36136 15113
rect 21088 15036 21140 15088
rect 23664 15036 23716 15088
rect 17868 15011 17920 15020
rect 17868 14977 17877 15011
rect 17877 14977 17911 15011
rect 17911 14977 17920 15011
rect 17868 14968 17920 14977
rect 19064 14968 19116 15020
rect 19340 14968 19392 15020
rect 20168 14968 20220 15020
rect 20720 15011 20772 15020
rect 20720 14977 20729 15011
rect 20729 14977 20763 15011
rect 20763 14977 20772 15011
rect 20720 14968 20772 14977
rect 20996 14968 21048 15020
rect 23020 14968 23072 15020
rect 25872 15011 25924 15020
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 27252 14968 27304 15020
rect 27988 15011 28040 15020
rect 27988 14977 27997 15011
rect 27997 14977 28031 15011
rect 28031 14977 28040 15011
rect 27988 14968 28040 14977
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 19984 14900 20036 14952
rect 22836 14900 22888 14952
rect 24860 14900 24912 14952
rect 25320 14943 25372 14952
rect 25320 14909 25329 14943
rect 25329 14909 25363 14943
rect 25363 14909 25372 14943
rect 25320 14900 25372 14909
rect 27344 14900 27396 14952
rect 28724 14968 28776 15020
rect 35992 14968 36044 15020
rect 29092 14900 29144 14952
rect 17408 14764 17460 14816
rect 23480 14832 23532 14884
rect 25136 14832 25188 14884
rect 26056 14832 26108 14884
rect 26148 14832 26200 14884
rect 26884 14832 26936 14884
rect 30840 14832 30892 14884
rect 24400 14764 24452 14816
rect 26240 14807 26292 14816
rect 26240 14773 26249 14807
rect 26249 14773 26283 14807
rect 26283 14773 26292 14807
rect 26240 14764 26292 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 17868 14560 17920 14612
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 22560 14560 22612 14612
rect 22836 14603 22888 14612
rect 22836 14569 22845 14603
rect 22845 14569 22879 14603
rect 22879 14569 22888 14603
rect 22836 14560 22888 14569
rect 23572 14560 23624 14612
rect 26608 14560 26660 14612
rect 27896 14560 27948 14612
rect 18512 14424 18564 14476
rect 20812 14467 20864 14476
rect 20812 14433 20821 14467
rect 20821 14433 20855 14467
rect 20855 14433 20864 14467
rect 20812 14424 20864 14433
rect 21088 14424 21140 14476
rect 27712 14492 27764 14544
rect 27988 14492 28040 14544
rect 30012 14492 30064 14544
rect 20720 14356 20772 14408
rect 21824 14356 21876 14408
rect 23388 14399 23440 14408
rect 2044 14288 2096 14340
rect 20812 14288 20864 14340
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 26148 14399 26200 14408
rect 26148 14365 26157 14399
rect 26157 14365 26191 14399
rect 26191 14365 26200 14399
rect 26148 14356 26200 14365
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 29000 14399 29052 14408
rect 29000 14365 29009 14399
rect 29009 14365 29043 14399
rect 29043 14365 29052 14399
rect 29000 14356 29052 14365
rect 29552 14356 29604 14408
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 19340 14220 19392 14272
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 24400 14288 24452 14340
rect 26608 14331 26660 14340
rect 26608 14297 26617 14331
rect 26617 14297 26651 14331
rect 26651 14297 26660 14331
rect 26608 14288 26660 14297
rect 19432 14220 19484 14229
rect 22284 14220 22336 14272
rect 26240 14220 26292 14272
rect 27712 14288 27764 14340
rect 27896 14331 27948 14340
rect 27896 14297 27905 14331
rect 27905 14297 27939 14331
rect 27939 14297 27948 14331
rect 27896 14288 27948 14297
rect 27988 14331 28040 14340
rect 27988 14297 27997 14331
rect 27997 14297 28031 14331
rect 28031 14297 28040 14331
rect 27988 14288 28040 14297
rect 28632 14288 28684 14340
rect 29736 14220 29788 14272
rect 34612 14220 34664 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 17040 14059 17092 14068
rect 17040 14025 17049 14059
rect 17049 14025 17083 14059
rect 17083 14025 17092 14059
rect 17040 14016 17092 14025
rect 17960 14016 18012 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 22100 14059 22152 14068
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 22744 14059 22796 14068
rect 22100 14016 22152 14025
rect 22744 14025 22753 14059
rect 22753 14025 22787 14059
rect 22787 14025 22796 14059
rect 22744 14016 22796 14025
rect 23388 14016 23440 14068
rect 19340 13948 19392 14000
rect 21824 13880 21876 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 23756 13991 23808 14000
rect 23756 13957 23765 13991
rect 23765 13957 23799 13991
rect 23799 13957 23808 13991
rect 23756 13948 23808 13957
rect 27804 14016 27856 14068
rect 28816 14059 28868 14068
rect 28816 14025 28825 14059
rect 28825 14025 28859 14059
rect 28859 14025 28868 14059
rect 28816 14016 28868 14025
rect 29000 14016 29052 14068
rect 29736 14016 29788 14068
rect 30840 14059 30892 14068
rect 30840 14025 30849 14059
rect 30849 14025 30883 14059
rect 30883 14025 30892 14059
rect 30840 14016 30892 14025
rect 25780 13991 25832 14000
rect 25780 13957 25789 13991
rect 25789 13957 25823 13991
rect 25823 13957 25832 13991
rect 25780 13948 25832 13957
rect 26240 13948 26292 14000
rect 22008 13880 22060 13889
rect 24860 13880 24912 13932
rect 25964 13880 26016 13932
rect 17960 13812 18012 13864
rect 18788 13855 18840 13864
rect 18788 13821 18797 13855
rect 18797 13821 18831 13855
rect 18831 13821 18840 13855
rect 18788 13812 18840 13821
rect 18972 13855 19024 13864
rect 18972 13821 18981 13855
rect 18981 13821 19015 13855
rect 19015 13821 19024 13855
rect 18972 13812 19024 13821
rect 22928 13812 22980 13864
rect 21180 13744 21232 13796
rect 23480 13812 23532 13864
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 18328 13676 18380 13728
rect 22376 13676 22428 13728
rect 23664 13744 23716 13796
rect 25504 13855 25556 13864
rect 25504 13821 25513 13855
rect 25513 13821 25547 13855
rect 25547 13821 25556 13855
rect 25504 13812 25556 13821
rect 26608 13812 26660 13864
rect 29368 13880 29420 13932
rect 27712 13812 27764 13864
rect 27528 13744 27580 13796
rect 28172 13787 28224 13796
rect 28172 13753 28181 13787
rect 28181 13753 28215 13787
rect 28215 13753 28224 13787
rect 28172 13744 28224 13753
rect 28816 13744 28868 13796
rect 33416 13880 33468 13932
rect 28448 13676 28500 13728
rect 28908 13676 28960 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 17960 13472 18012 13524
rect 18972 13472 19024 13524
rect 22192 13472 22244 13524
rect 22468 13472 22520 13524
rect 25044 13472 25096 13524
rect 25964 13472 26016 13524
rect 26056 13472 26108 13524
rect 28632 13472 28684 13524
rect 23664 13404 23716 13456
rect 19340 13336 19392 13388
rect 23388 13336 23440 13388
rect 18328 13268 18380 13320
rect 22192 13311 22244 13320
rect 19156 13132 19208 13184
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 19340 13200 19392 13252
rect 20168 13243 20220 13252
rect 20168 13209 20177 13243
rect 20177 13209 20211 13243
rect 20211 13209 20220 13243
rect 20168 13200 20220 13209
rect 20628 13200 20680 13252
rect 22928 13243 22980 13252
rect 22928 13209 22937 13243
rect 22937 13209 22971 13243
rect 22971 13209 22980 13243
rect 22928 13200 22980 13209
rect 20444 13132 20496 13184
rect 23572 13243 23624 13252
rect 23572 13209 23581 13243
rect 23581 13209 23615 13243
rect 23615 13209 23624 13243
rect 23572 13200 23624 13209
rect 25780 13336 25832 13388
rect 26056 13379 26108 13388
rect 26056 13345 26065 13379
rect 26065 13345 26099 13379
rect 26099 13345 26108 13379
rect 26056 13336 26108 13345
rect 26608 13379 26660 13388
rect 26608 13345 26617 13379
rect 26617 13345 26651 13379
rect 26651 13345 26660 13379
rect 26608 13336 26660 13345
rect 28448 13336 28500 13388
rect 25044 13268 25096 13320
rect 29184 13268 29236 13320
rect 35992 13268 36044 13320
rect 24308 13200 24360 13252
rect 25320 13200 25372 13252
rect 25964 13243 26016 13252
rect 25964 13209 25973 13243
rect 25973 13209 26007 13243
rect 26007 13209 26016 13243
rect 25964 13200 26016 13209
rect 24584 13175 24636 13184
rect 24584 13141 24593 13175
rect 24593 13141 24627 13175
rect 24627 13141 24636 13175
rect 24584 13132 24636 13141
rect 27436 13200 27488 13252
rect 27528 13200 27580 13252
rect 28172 13200 28224 13252
rect 27988 13132 28040 13184
rect 36268 13175 36320 13184
rect 36268 13141 36277 13175
rect 36277 13141 36311 13175
rect 36311 13141 36320 13175
rect 36268 13132 36320 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1860 12928 1912 12980
rect 2688 12928 2740 12980
rect 5632 12860 5684 12912
rect 18328 12860 18380 12912
rect 19432 12928 19484 12980
rect 20720 12928 20772 12980
rect 21824 12928 21876 12980
rect 24584 12928 24636 12980
rect 17684 12792 17736 12844
rect 18788 12792 18840 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20168 12860 20220 12912
rect 21180 12792 21232 12844
rect 18236 12724 18288 12776
rect 20352 12656 20404 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 19340 12588 19392 12640
rect 19984 12588 20036 12640
rect 20536 12631 20588 12640
rect 20536 12597 20545 12631
rect 20545 12597 20579 12631
rect 20579 12597 20588 12631
rect 20536 12588 20588 12597
rect 22192 12860 22244 12912
rect 23480 12860 23532 12912
rect 27160 12860 27212 12912
rect 28264 12860 28316 12912
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 25780 12724 25832 12776
rect 24308 12699 24360 12708
rect 24308 12665 24317 12699
rect 24317 12665 24351 12699
rect 24351 12665 24360 12699
rect 24308 12656 24360 12665
rect 23848 12588 23900 12640
rect 26148 12835 26200 12844
rect 26148 12801 26157 12835
rect 26157 12801 26191 12835
rect 26191 12801 26200 12835
rect 26148 12792 26200 12801
rect 28080 12792 28132 12844
rect 26608 12724 26660 12776
rect 27436 12724 27488 12776
rect 29184 12724 29236 12776
rect 27712 12656 27764 12708
rect 29092 12656 29144 12708
rect 26148 12588 26200 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 17684 12427 17736 12436
rect 17684 12393 17693 12427
rect 17693 12393 17727 12427
rect 17727 12393 17736 12427
rect 17684 12384 17736 12393
rect 20628 12427 20680 12436
rect 14464 12316 14516 12368
rect 18236 12316 18288 12368
rect 19984 12316 20036 12368
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 21180 12427 21232 12436
rect 21180 12393 21189 12427
rect 21189 12393 21223 12427
rect 21223 12393 21232 12427
rect 21180 12384 21232 12393
rect 23204 12384 23256 12436
rect 24492 12384 24544 12436
rect 22928 12316 22980 12368
rect 27988 12384 28040 12436
rect 28356 12384 28408 12436
rect 29092 12427 29144 12436
rect 29092 12393 29101 12427
rect 29101 12393 29135 12427
rect 29135 12393 29144 12427
rect 29092 12384 29144 12393
rect 18052 12248 18104 12300
rect 22008 12248 22060 12300
rect 23572 12291 23624 12300
rect 23572 12257 23581 12291
rect 23581 12257 23615 12291
rect 23615 12257 23624 12291
rect 36176 12384 36228 12436
rect 23572 12248 23624 12257
rect 27712 12248 27764 12300
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 13268 12180 13320 12232
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 18144 12180 18196 12232
rect 17592 12112 17644 12164
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 20444 12180 20496 12232
rect 21180 12180 21232 12232
rect 24492 12180 24544 12232
rect 27344 12223 27396 12232
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 27896 12180 27948 12232
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 18512 12112 18564 12164
rect 19064 12112 19116 12164
rect 21456 12112 21508 12164
rect 22928 12155 22980 12164
rect 1860 12044 1912 12096
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 17500 12044 17552 12096
rect 19616 12044 19668 12096
rect 22928 12121 22937 12155
rect 22937 12121 22971 12155
rect 22971 12121 22980 12155
rect 22928 12112 22980 12121
rect 23480 12155 23532 12164
rect 23480 12121 23489 12155
rect 23489 12121 23523 12155
rect 23523 12121 23532 12155
rect 23480 12112 23532 12121
rect 29828 12112 29880 12164
rect 27344 12044 27396 12096
rect 28816 12044 28868 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 18144 11883 18196 11892
rect 18144 11849 18153 11883
rect 18153 11849 18187 11883
rect 18187 11849 18196 11883
rect 18144 11840 18196 11849
rect 8116 11772 8168 11824
rect 17040 11772 17092 11824
rect 18788 11772 18840 11824
rect 20352 11772 20404 11824
rect 20628 11772 20680 11824
rect 22192 11840 22244 11892
rect 23756 11840 23808 11892
rect 24676 11772 24728 11824
rect 26148 11840 26200 11892
rect 27160 11840 27212 11892
rect 27804 11840 27856 11892
rect 29828 11883 29880 11892
rect 29828 11849 29837 11883
rect 29837 11849 29871 11883
rect 29871 11849 29880 11883
rect 29828 11840 29880 11849
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 26056 11772 26108 11824
rect 27712 11772 27764 11824
rect 18052 11704 18104 11756
rect 18144 11636 18196 11688
rect 20996 11704 21048 11756
rect 23204 11704 23256 11756
rect 23664 11704 23716 11756
rect 5540 11500 5592 11552
rect 18880 11568 18932 11620
rect 20260 11568 20312 11620
rect 19984 11500 20036 11552
rect 20352 11500 20404 11552
rect 21088 11500 21140 11552
rect 21824 11500 21876 11552
rect 23756 11636 23808 11688
rect 26884 11704 26936 11756
rect 27528 11704 27580 11756
rect 27804 11747 27856 11756
rect 27804 11713 27813 11747
rect 27813 11713 27847 11747
rect 27847 11713 27856 11747
rect 27804 11704 27856 11713
rect 28540 11704 28592 11756
rect 29184 11704 29236 11756
rect 29736 11747 29788 11756
rect 29736 11713 29745 11747
rect 29745 11713 29779 11747
rect 29779 11713 29788 11747
rect 29736 11704 29788 11713
rect 22744 11568 22796 11620
rect 27620 11636 27672 11688
rect 25780 11568 25832 11620
rect 35440 11636 35492 11688
rect 24124 11500 24176 11552
rect 24308 11500 24360 11552
rect 27804 11500 27856 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 17500 11339 17552 11348
rect 17500 11305 17509 11339
rect 17509 11305 17543 11339
rect 17543 11305 17552 11339
rect 17500 11296 17552 11305
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 18880 11296 18932 11348
rect 24492 11296 24544 11348
rect 24676 11339 24728 11348
rect 24676 11305 24685 11339
rect 24685 11305 24719 11339
rect 24719 11305 24728 11339
rect 24676 11296 24728 11305
rect 24768 11296 24820 11348
rect 28908 11296 28960 11348
rect 29000 11296 29052 11348
rect 18972 11228 19024 11280
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 19064 11160 19116 11212
rect 20168 11160 20220 11212
rect 21364 11228 21416 11280
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18512 11092 18564 11144
rect 19340 11092 19392 11144
rect 19248 11024 19300 11076
rect 20536 11067 20588 11076
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 19340 10956 19392 11008
rect 20536 11033 20545 11067
rect 20545 11033 20579 11067
rect 20579 11033 20588 11067
rect 20536 11024 20588 11033
rect 22008 11228 22060 11280
rect 25320 11228 25372 11280
rect 22928 11203 22980 11212
rect 22928 11169 22937 11203
rect 22937 11169 22971 11203
rect 22971 11169 22980 11203
rect 22928 11160 22980 11169
rect 25228 11160 25280 11212
rect 26148 11160 26200 11212
rect 27712 11203 27764 11212
rect 27712 11169 27721 11203
rect 27721 11169 27755 11203
rect 27755 11169 27764 11203
rect 27712 11160 27764 11169
rect 23204 11092 23256 11144
rect 23756 11092 23808 11144
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 22100 10956 22152 11008
rect 23940 11024 23992 11076
rect 24032 11024 24084 11076
rect 25504 11067 25556 11076
rect 25504 11033 25513 11067
rect 25513 11033 25547 11067
rect 25547 11033 25556 11067
rect 25504 11024 25556 11033
rect 25780 11024 25832 11076
rect 28540 11135 28592 11144
rect 28540 11101 28549 11135
rect 28549 11101 28583 11135
rect 28583 11101 28592 11135
rect 28540 11092 28592 11101
rect 30104 11092 30156 11144
rect 36084 11135 36136 11144
rect 36084 11101 36093 11135
rect 36093 11101 36127 11135
rect 36127 11101 36136 11135
rect 36084 11092 36136 11101
rect 31484 11024 31536 11076
rect 36268 11067 36320 11076
rect 36268 11033 36277 11067
rect 36277 11033 36311 11067
rect 36311 11033 36320 11067
rect 36268 11024 36320 11033
rect 27620 10956 27672 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 18052 10752 18104 10804
rect 19524 10752 19576 10804
rect 18144 10684 18196 10736
rect 19248 10684 19300 10736
rect 21732 10752 21784 10804
rect 23296 10684 23348 10736
rect 24492 10727 24544 10736
rect 24492 10693 24501 10727
rect 24501 10693 24535 10727
rect 24535 10693 24544 10727
rect 24492 10684 24544 10693
rect 30012 10752 30064 10804
rect 26148 10684 26200 10736
rect 27896 10684 27948 10736
rect 28080 10684 28132 10736
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 28632 10616 28684 10668
rect 29000 10616 29052 10668
rect 19432 10548 19484 10600
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 19984 10548 20036 10600
rect 20812 10548 20864 10600
rect 22744 10548 22796 10600
rect 23020 10591 23072 10600
rect 23020 10557 23029 10591
rect 23029 10557 23063 10591
rect 23063 10557 23072 10591
rect 23020 10548 23072 10557
rect 23296 10548 23348 10600
rect 23664 10548 23716 10600
rect 24768 10548 24820 10600
rect 26976 10548 27028 10600
rect 27712 10591 27764 10600
rect 27712 10557 27721 10591
rect 27721 10557 27755 10591
rect 27755 10557 27764 10591
rect 27712 10548 27764 10557
rect 29276 10548 29328 10600
rect 6092 10480 6144 10532
rect 18972 10412 19024 10464
rect 19248 10412 19300 10464
rect 22836 10412 22888 10464
rect 23296 10412 23348 10464
rect 25044 10412 25096 10464
rect 26424 10480 26476 10532
rect 28448 10480 28500 10532
rect 27620 10412 27672 10464
rect 36544 10412 36596 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5632 10208 5684 10260
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 19340 10208 19392 10260
rect 19616 10208 19668 10260
rect 21640 10208 21692 10260
rect 23112 10208 23164 10260
rect 24768 10208 24820 10260
rect 25504 10208 25556 10260
rect 26240 10208 26292 10260
rect 28264 10208 28316 10260
rect 22192 10183 22244 10192
rect 22192 10149 22201 10183
rect 22201 10149 22235 10183
rect 22235 10149 22244 10183
rect 22192 10140 22244 10149
rect 22928 10140 22980 10192
rect 26424 10183 26476 10192
rect 26424 10149 26433 10183
rect 26433 10149 26467 10183
rect 26467 10149 26476 10183
rect 26424 10140 26476 10149
rect 26976 10183 27028 10192
rect 26976 10149 26985 10183
rect 26985 10149 27019 10183
rect 27019 10149 27028 10183
rect 26976 10140 27028 10149
rect 19340 10072 19392 10124
rect 22468 10072 22520 10124
rect 22836 10115 22888 10124
rect 22836 10081 22845 10115
rect 22845 10081 22879 10115
rect 22879 10081 22888 10115
rect 22836 10072 22888 10081
rect 23020 10072 23072 10124
rect 23204 10072 23256 10124
rect 27620 10047 27672 10056
rect 27620 10013 27629 10047
rect 27629 10013 27663 10047
rect 27663 10013 27672 10047
rect 27620 10004 27672 10013
rect 28356 10004 28408 10056
rect 29460 10004 29512 10056
rect 36360 10047 36412 10056
rect 36360 10013 36369 10047
rect 36369 10013 36403 10047
rect 36403 10013 36412 10047
rect 36360 10004 36412 10013
rect 19340 9936 19392 9988
rect 17868 9868 17920 9920
rect 19616 9868 19668 9920
rect 19984 9936 20036 9988
rect 20536 9936 20588 9988
rect 20168 9868 20220 9920
rect 20260 9868 20312 9920
rect 21732 9979 21784 9988
rect 21732 9945 21741 9979
rect 21741 9945 21775 9979
rect 21775 9945 21784 9979
rect 21732 9936 21784 9945
rect 24124 9936 24176 9988
rect 24676 9868 24728 9920
rect 35624 9868 35676 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 20076 9664 20128 9716
rect 20720 9664 20772 9716
rect 21732 9664 21784 9716
rect 23296 9664 23348 9716
rect 23572 9664 23624 9716
rect 12808 9596 12860 9648
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 19156 9596 19208 9648
rect 22560 9596 22612 9648
rect 24768 9596 24820 9648
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 18788 9460 18840 9469
rect 21548 9460 21600 9512
rect 22008 9503 22060 9512
rect 22008 9469 22017 9503
rect 22017 9469 22051 9503
rect 22051 9469 22060 9503
rect 22008 9460 22060 9469
rect 21916 9392 21968 9444
rect 18420 9324 18472 9376
rect 19064 9324 19116 9376
rect 22652 9460 22704 9512
rect 24216 9503 24268 9512
rect 24216 9469 24225 9503
rect 24225 9469 24259 9503
rect 24259 9469 24268 9503
rect 24216 9460 24268 9469
rect 23572 9392 23624 9444
rect 26792 9596 26844 9648
rect 27896 9639 27948 9648
rect 27896 9605 27905 9639
rect 27905 9605 27939 9639
rect 27939 9605 27948 9639
rect 27896 9596 27948 9605
rect 31024 9596 31076 9648
rect 36360 9639 36412 9648
rect 36360 9605 36369 9639
rect 36369 9605 36403 9639
rect 36403 9605 36412 9639
rect 36360 9596 36412 9605
rect 27068 9528 27120 9580
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 27436 9528 27488 9580
rect 32772 9460 32824 9512
rect 23756 9367 23808 9376
rect 23756 9333 23765 9367
rect 23765 9333 23799 9367
rect 23799 9333 23808 9367
rect 23756 9324 23808 9333
rect 24308 9324 24360 9376
rect 24676 9324 24728 9376
rect 29184 9392 29236 9444
rect 32312 9392 32364 9444
rect 25964 9367 26016 9376
rect 25964 9333 25973 9367
rect 25973 9333 26007 9367
rect 26007 9333 26016 9367
rect 25964 9324 26016 9333
rect 27160 9324 27212 9376
rect 28448 9324 28500 9376
rect 32864 9324 32916 9376
rect 34796 9324 34848 9376
rect 36176 9324 36228 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6552 9120 6604 9172
rect 19432 9120 19484 9172
rect 20260 9120 20312 9172
rect 20444 9120 20496 9172
rect 17592 9052 17644 9104
rect 21456 9052 21508 9104
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 19340 8984 19392 9036
rect 20076 8984 20128 9036
rect 22192 9120 22244 9172
rect 24032 9120 24084 9172
rect 25964 9120 26016 9172
rect 27620 9120 27672 9172
rect 28172 9120 28224 9172
rect 29368 9120 29420 9172
rect 32312 9163 32364 9172
rect 22928 9052 22980 9104
rect 23388 9052 23440 9104
rect 23756 9052 23808 9104
rect 22008 8984 22060 9036
rect 24216 8984 24268 9036
rect 28264 9052 28316 9104
rect 31392 9052 31444 9104
rect 32312 9129 32321 9163
rect 32321 9129 32355 9163
rect 32355 9129 32364 9163
rect 32312 9120 32364 9129
rect 32864 9163 32916 9172
rect 32864 9129 32873 9163
rect 32873 9129 32907 9163
rect 32907 9129 32916 9163
rect 32864 9120 32916 9129
rect 33140 9052 33192 9104
rect 25228 8984 25280 9036
rect 17224 8916 17276 8968
rect 17960 8916 18012 8968
rect 19248 8916 19300 8968
rect 25964 8916 26016 8968
rect 29184 8984 29236 9036
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 21824 8848 21876 8900
rect 22468 8848 22520 8900
rect 23848 8891 23900 8900
rect 20812 8780 20864 8832
rect 20996 8780 21048 8832
rect 21732 8780 21784 8832
rect 23848 8857 23857 8891
rect 23857 8857 23891 8891
rect 23891 8857 23900 8891
rect 23848 8848 23900 8857
rect 24124 8848 24176 8900
rect 23388 8780 23440 8832
rect 25136 8848 25188 8900
rect 34520 8916 34572 8968
rect 30472 8848 30524 8900
rect 35900 8891 35952 8900
rect 35900 8857 35909 8891
rect 35909 8857 35943 8891
rect 35943 8857 35952 8891
rect 35900 8848 35952 8857
rect 28448 8780 28500 8832
rect 28632 8780 28684 8832
rect 29184 8780 29236 8832
rect 34244 8780 34296 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 17776 8576 17828 8628
rect 19524 8576 19576 8628
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 20904 8576 20956 8628
rect 19892 8551 19944 8560
rect 19892 8517 19901 8551
rect 19901 8517 19935 8551
rect 19935 8517 19944 8551
rect 19892 8508 19944 8517
rect 20996 8440 21048 8492
rect 21548 8576 21600 8628
rect 36084 8576 36136 8628
rect 23296 8508 23348 8560
rect 28264 8508 28316 8560
rect 31576 8508 31628 8560
rect 31852 8508 31904 8560
rect 32312 8508 32364 8560
rect 22100 8440 22152 8492
rect 24216 8440 24268 8492
rect 28172 8440 28224 8492
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 19340 8372 19392 8424
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 24676 8372 24728 8424
rect 19432 8236 19484 8288
rect 21732 8304 21784 8356
rect 22100 8347 22152 8356
rect 22100 8313 22109 8347
rect 22109 8313 22143 8347
rect 22143 8313 22152 8347
rect 27528 8372 27580 8424
rect 22100 8304 22152 8313
rect 21180 8236 21232 8288
rect 21456 8236 21508 8288
rect 27436 8304 27488 8356
rect 30288 8304 30340 8356
rect 31760 8304 31812 8356
rect 34520 8304 34572 8356
rect 35348 8304 35400 8356
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 26056 8279 26108 8288
rect 26056 8245 26065 8279
rect 26065 8245 26099 8279
rect 26099 8245 26108 8279
rect 26056 8236 26108 8245
rect 34152 8236 34204 8288
rect 35440 8279 35492 8288
rect 35440 8245 35449 8279
rect 35449 8245 35483 8279
rect 35483 8245 35492 8279
rect 35440 8236 35492 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 22192 8032 22244 8084
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 24492 8032 24544 8084
rect 26056 8032 26108 8084
rect 29092 8032 29144 8084
rect 31208 8032 31260 8084
rect 31852 8032 31904 8084
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 23020 7964 23072 8016
rect 28724 7964 28776 8016
rect 33416 7964 33468 8016
rect 24124 7896 24176 7948
rect 24676 7896 24728 7948
rect 26148 7896 26200 7948
rect 29184 7896 29236 7948
rect 32864 7896 32916 7948
rect 20812 7828 20864 7880
rect 23664 7828 23716 7880
rect 24032 7871 24084 7880
rect 24032 7837 24041 7871
rect 24041 7837 24075 7871
rect 24075 7837 24084 7871
rect 24032 7828 24084 7837
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 29644 7828 29696 7880
rect 29920 7828 29972 7880
rect 34520 7896 34572 7948
rect 35440 7896 35492 7948
rect 36360 7871 36412 7880
rect 36360 7837 36369 7871
rect 36369 7837 36403 7871
rect 36403 7837 36412 7871
rect 36360 7828 36412 7837
rect 21180 7803 21232 7812
rect 19064 7692 19116 7744
rect 19248 7692 19300 7744
rect 21180 7769 21189 7803
rect 21189 7769 21223 7803
rect 21223 7769 21232 7803
rect 21180 7760 21232 7769
rect 22744 7692 22796 7744
rect 22836 7692 22888 7744
rect 24032 7692 24084 7744
rect 29184 7692 29236 7744
rect 30288 7692 30340 7744
rect 32128 7760 32180 7812
rect 32036 7692 32088 7744
rect 32312 7735 32364 7744
rect 32312 7701 32321 7735
rect 32321 7701 32355 7735
rect 32355 7701 32364 7735
rect 32312 7692 32364 7701
rect 34152 7735 34204 7744
rect 34152 7701 34161 7735
rect 34161 7701 34195 7735
rect 34195 7701 34204 7735
rect 34152 7692 34204 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 20536 7488 20588 7540
rect 22192 7488 22244 7540
rect 23848 7488 23900 7540
rect 18236 7463 18288 7472
rect 18236 7429 18245 7463
rect 18245 7429 18279 7463
rect 18279 7429 18288 7463
rect 18236 7420 18288 7429
rect 19064 7463 19116 7472
rect 19064 7429 19073 7463
rect 19073 7429 19107 7463
rect 19107 7429 19116 7463
rect 19064 7420 19116 7429
rect 19340 7420 19392 7472
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 23756 7420 23808 7472
rect 23020 7352 23072 7404
rect 24308 7420 24360 7472
rect 26148 7488 26200 7540
rect 28908 7488 28960 7540
rect 36360 7531 36412 7540
rect 26516 7420 26568 7472
rect 27252 7420 27304 7472
rect 31760 7420 31812 7472
rect 25412 7352 25464 7404
rect 25964 7352 26016 7404
rect 27344 7352 27396 7404
rect 31208 7395 31260 7404
rect 31208 7361 31217 7395
rect 31217 7361 31251 7395
rect 31251 7361 31260 7395
rect 31208 7352 31260 7361
rect 34704 7420 34756 7472
rect 35348 7420 35400 7472
rect 36360 7497 36369 7531
rect 36369 7497 36403 7531
rect 36403 7497 36412 7531
rect 36360 7488 36412 7497
rect 36452 7420 36504 7472
rect 19432 7284 19484 7336
rect 20260 7284 20312 7336
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 20720 7284 20772 7336
rect 24032 7327 24084 7336
rect 24032 7293 24041 7327
rect 24041 7293 24075 7327
rect 24075 7293 24084 7327
rect 24308 7327 24360 7336
rect 24032 7284 24084 7293
rect 24308 7293 24317 7327
rect 24317 7293 24351 7327
rect 24351 7293 24360 7327
rect 24308 7284 24360 7293
rect 27896 7284 27948 7336
rect 28908 7327 28960 7336
rect 28908 7293 28917 7327
rect 28917 7293 28951 7327
rect 28951 7293 28960 7327
rect 28908 7284 28960 7293
rect 29184 7327 29236 7336
rect 29184 7293 29193 7327
rect 29193 7293 29227 7327
rect 29227 7293 29236 7327
rect 29184 7284 29236 7293
rect 32312 7352 32364 7404
rect 18604 7216 18656 7268
rect 19248 7216 19300 7268
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 19340 7148 19392 7200
rect 21180 7148 21232 7200
rect 22744 7148 22796 7200
rect 25504 7148 25556 7200
rect 28448 7148 28500 7200
rect 30932 7216 30984 7268
rect 32772 7352 32824 7404
rect 34152 7352 34204 7404
rect 35532 7352 35584 7404
rect 34704 7216 34756 7268
rect 31852 7148 31904 7200
rect 31944 7148 31996 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19432 6944 19484 6996
rect 25412 6944 25464 6996
rect 32956 6944 33008 6996
rect 35532 6987 35584 6996
rect 35532 6953 35541 6987
rect 35541 6953 35575 6987
rect 35575 6953 35584 6987
rect 35532 6944 35584 6953
rect 18236 6808 18288 6860
rect 1952 6740 2004 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 17592 6740 17644 6792
rect 20628 6808 20680 6860
rect 20812 6851 20864 6860
rect 20812 6817 20821 6851
rect 20821 6817 20855 6851
rect 20855 6817 20864 6851
rect 20812 6808 20864 6817
rect 21640 6808 21692 6860
rect 23204 6808 23256 6860
rect 24032 6808 24084 6860
rect 26056 6808 26108 6860
rect 26332 6808 26384 6860
rect 29368 6876 29420 6928
rect 29552 6876 29604 6928
rect 27344 6808 27396 6860
rect 32588 6808 32640 6860
rect 32864 6851 32916 6860
rect 32864 6817 32873 6851
rect 32873 6817 32907 6851
rect 32907 6817 32916 6851
rect 32864 6808 32916 6817
rect 33048 6808 33100 6860
rect 34520 6808 34572 6860
rect 19340 6740 19392 6792
rect 18972 6672 19024 6724
rect 18512 6604 18564 6656
rect 21180 6672 21232 6724
rect 21364 6672 21416 6724
rect 25688 6672 25740 6724
rect 26240 6672 26292 6724
rect 31852 6740 31904 6792
rect 32772 6740 32824 6792
rect 33232 6740 33284 6792
rect 33692 6740 33744 6792
rect 34704 6740 34756 6792
rect 35072 6783 35124 6792
rect 35072 6749 35081 6783
rect 35081 6749 35115 6783
rect 35115 6749 35124 6783
rect 35072 6740 35124 6749
rect 34520 6672 34572 6724
rect 20260 6604 20312 6656
rect 23020 6604 23072 6656
rect 24400 6604 24452 6656
rect 24768 6604 24820 6656
rect 24952 6604 25004 6656
rect 25780 6604 25832 6656
rect 27988 6604 28040 6656
rect 28080 6647 28132 6656
rect 28080 6613 28089 6647
rect 28089 6613 28123 6647
rect 28123 6613 28132 6647
rect 28080 6604 28132 6613
rect 29184 6647 29236 6656
rect 29184 6613 29193 6647
rect 29193 6613 29227 6647
rect 29227 6613 29236 6647
rect 29184 6604 29236 6613
rect 29552 6604 29604 6656
rect 30748 6647 30800 6656
rect 30748 6613 30757 6647
rect 30757 6613 30791 6647
rect 30791 6613 30800 6647
rect 30748 6604 30800 6613
rect 31116 6604 31168 6656
rect 32404 6604 32456 6656
rect 33232 6604 33284 6656
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 33600 6604 33652 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1860 6400 1912 6452
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 17500 6332 17552 6384
rect 20812 6400 20864 6452
rect 22192 6400 22244 6452
rect 24400 6400 24452 6452
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 18696 6264 18748 6316
rect 18972 6264 19024 6316
rect 18604 6196 18656 6248
rect 20260 6332 20312 6384
rect 30380 6400 30432 6452
rect 31392 6400 31444 6452
rect 32588 6443 32640 6452
rect 32588 6409 32597 6443
rect 32597 6409 32631 6443
rect 32631 6409 32640 6443
rect 32588 6400 32640 6409
rect 32772 6400 32824 6452
rect 33600 6400 33652 6452
rect 34520 6443 34572 6452
rect 34520 6409 34529 6443
rect 34529 6409 34563 6443
rect 34563 6409 34572 6443
rect 34520 6400 34572 6409
rect 35532 6400 35584 6452
rect 22008 6264 22060 6316
rect 19616 6128 19668 6180
rect 20444 6060 20496 6112
rect 22192 6060 22244 6112
rect 24952 6332 25004 6384
rect 27528 6332 27580 6384
rect 33508 6332 33560 6384
rect 24032 6264 24084 6316
rect 26608 6239 26660 6248
rect 26608 6205 26617 6239
rect 26617 6205 26651 6239
rect 26651 6205 26660 6239
rect 26608 6196 26660 6205
rect 30564 6264 30616 6316
rect 31852 6264 31904 6316
rect 32680 6307 32732 6316
rect 32680 6273 32689 6307
rect 32689 6273 32723 6307
rect 32723 6273 32732 6307
rect 32680 6264 32732 6273
rect 32864 6264 32916 6316
rect 33692 6264 33744 6316
rect 35072 6332 35124 6384
rect 35440 6332 35492 6384
rect 29276 6239 29328 6248
rect 29276 6205 29285 6239
rect 29285 6205 29319 6239
rect 29319 6205 29328 6239
rect 29276 6196 29328 6205
rect 23848 6128 23900 6180
rect 24584 6128 24636 6180
rect 27160 6103 27212 6112
rect 27160 6069 27169 6103
rect 27169 6069 27203 6103
rect 27203 6069 27212 6103
rect 27160 6060 27212 6069
rect 30472 6196 30524 6248
rect 29644 6128 29696 6180
rect 29184 6060 29236 6112
rect 29552 6060 29604 6112
rect 30472 6060 30524 6112
rect 31576 6060 31628 6112
rect 32588 6060 32640 6112
rect 32680 6060 32732 6112
rect 34520 6196 34572 6248
rect 34704 6196 34756 6248
rect 34704 6060 34756 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 17960 5856 18012 5908
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 22100 5856 22152 5908
rect 2320 5652 2372 5704
rect 17776 5652 17828 5704
rect 18696 5720 18748 5772
rect 20812 5763 20864 5772
rect 20812 5729 20821 5763
rect 20821 5729 20855 5763
rect 20855 5729 20864 5763
rect 20812 5720 20864 5729
rect 22928 5720 22980 5772
rect 20352 5652 20404 5704
rect 19616 5627 19668 5636
rect 19616 5593 19625 5627
rect 19625 5593 19659 5627
rect 19659 5593 19668 5627
rect 19616 5584 19668 5593
rect 20444 5584 20496 5636
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 17868 5516 17920 5568
rect 18788 5516 18840 5568
rect 21180 5516 21232 5568
rect 26608 5788 26660 5840
rect 23848 5720 23900 5772
rect 27252 5788 27304 5840
rect 27160 5720 27212 5772
rect 28080 5720 28132 5772
rect 29092 5899 29144 5908
rect 29092 5865 29101 5899
rect 29101 5865 29135 5899
rect 29135 5865 29144 5899
rect 29092 5856 29144 5865
rect 28724 5788 28776 5840
rect 31484 5899 31536 5908
rect 31484 5865 31493 5899
rect 31493 5865 31527 5899
rect 31527 5865 31536 5899
rect 31484 5856 31536 5865
rect 32036 5899 32088 5908
rect 32036 5865 32045 5899
rect 32045 5865 32079 5899
rect 32079 5865 32088 5899
rect 32036 5856 32088 5865
rect 32588 5856 32640 5908
rect 31024 5788 31076 5840
rect 32956 5856 33008 5908
rect 32312 5720 32364 5772
rect 25688 5652 25740 5704
rect 26148 5584 26200 5636
rect 25504 5559 25556 5568
rect 25504 5525 25513 5559
rect 25513 5525 25547 5559
rect 25547 5525 25556 5559
rect 25504 5516 25556 5525
rect 26056 5559 26108 5568
rect 26056 5525 26065 5559
rect 26065 5525 26099 5559
rect 26099 5525 26108 5559
rect 26056 5516 26108 5525
rect 29644 5652 29696 5704
rect 31116 5652 31168 5704
rect 31668 5652 31720 5704
rect 33140 5720 33192 5772
rect 27620 5627 27672 5636
rect 27620 5593 27629 5627
rect 27629 5593 27663 5627
rect 27663 5593 27672 5627
rect 27620 5584 27672 5593
rect 29828 5516 29880 5568
rect 32680 5584 32732 5636
rect 33784 5652 33836 5704
rect 34060 5695 34112 5704
rect 34060 5661 34069 5695
rect 34069 5661 34103 5695
rect 34103 5661 34112 5695
rect 34060 5652 34112 5661
rect 35440 5652 35492 5704
rect 36360 5695 36412 5704
rect 36360 5661 36369 5695
rect 36369 5661 36403 5695
rect 36403 5661 36412 5695
rect 36360 5652 36412 5661
rect 31760 5516 31812 5568
rect 33140 5516 33192 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 19156 5312 19208 5364
rect 19984 5312 20036 5364
rect 22008 5312 22060 5364
rect 16764 5244 16816 5296
rect 20076 5244 20128 5296
rect 13544 5176 13596 5228
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 17960 5108 18012 5160
rect 15292 5040 15344 5092
rect 17592 5040 17644 5092
rect 22928 5108 22980 5160
rect 20812 5040 20864 5092
rect 22008 5083 22060 5092
rect 22008 5049 22017 5083
rect 22017 5049 22051 5083
rect 22051 5049 22060 5083
rect 22008 5040 22060 5049
rect 29000 5312 29052 5364
rect 33048 5312 33100 5364
rect 33784 5312 33836 5364
rect 34428 5312 34480 5364
rect 35440 5355 35492 5364
rect 35440 5321 35449 5355
rect 35449 5321 35483 5355
rect 35483 5321 35492 5355
rect 35440 5312 35492 5321
rect 27160 5219 27212 5228
rect 27160 5185 27169 5219
rect 27169 5185 27203 5219
rect 27203 5185 27212 5219
rect 27160 5176 27212 5185
rect 30380 5287 30432 5296
rect 30380 5253 30389 5287
rect 30389 5253 30423 5287
rect 30423 5253 30432 5287
rect 30380 5244 30432 5253
rect 30564 5244 30616 5296
rect 30748 5244 30800 5296
rect 29092 5176 29144 5228
rect 30104 5176 30156 5228
rect 30472 5219 30524 5228
rect 30472 5185 30481 5219
rect 30481 5185 30515 5219
rect 30515 5185 30524 5219
rect 30472 5176 30524 5185
rect 31668 5244 31720 5296
rect 27528 5108 27580 5160
rect 26424 5040 26476 5092
rect 29184 5108 29236 5160
rect 31760 5219 31812 5228
rect 31760 5185 31769 5219
rect 31769 5185 31803 5219
rect 31803 5185 31812 5219
rect 31760 5176 31812 5185
rect 32404 5219 32456 5228
rect 32404 5185 32413 5219
rect 32413 5185 32447 5219
rect 32447 5185 32456 5219
rect 32404 5176 32456 5185
rect 32864 5244 32916 5296
rect 33232 5176 33284 5228
rect 33508 5176 33560 5228
rect 34060 5176 34112 5228
rect 30748 5108 30800 5160
rect 32588 5040 32640 5092
rect 33048 5083 33100 5092
rect 33048 5049 33057 5083
rect 33057 5049 33091 5083
rect 33091 5049 33100 5083
rect 33048 5040 33100 5049
rect 33508 5040 33560 5092
rect 34060 5040 34112 5092
rect 23664 5015 23716 5024
rect 23664 4981 23673 5015
rect 23673 4981 23707 5015
rect 23707 4981 23716 5015
rect 23664 4972 23716 4981
rect 24124 5015 24176 5024
rect 24124 4981 24133 5015
rect 24133 4981 24167 5015
rect 24167 4981 24176 5015
rect 24124 4972 24176 4981
rect 26056 5015 26108 5024
rect 26056 4981 26065 5015
rect 26065 4981 26099 5015
rect 26099 4981 26108 5015
rect 26056 4972 26108 4981
rect 29092 4972 29144 5024
rect 29644 5015 29696 5024
rect 29644 4981 29653 5015
rect 29653 4981 29687 5015
rect 29687 4981 29696 5015
rect 29644 4972 29696 4981
rect 29828 4972 29880 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 16764 4811 16816 4820
rect 16764 4777 16773 4811
rect 16773 4777 16807 4811
rect 16807 4777 16816 4811
rect 16764 4768 16816 4777
rect 22652 4811 22704 4820
rect 17776 4700 17828 4752
rect 22652 4777 22661 4811
rect 22661 4777 22695 4811
rect 22695 4777 22704 4811
rect 22652 4768 22704 4777
rect 25228 4768 25280 4820
rect 33048 4768 33100 4820
rect 35440 4811 35492 4820
rect 35440 4777 35449 4811
rect 35449 4777 35483 4811
rect 35483 4777 35492 4811
rect 35440 4768 35492 4777
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 20812 4632 20864 4684
rect 21640 4632 21692 4684
rect 23664 4632 23716 4684
rect 26056 4632 26108 4684
rect 27160 4632 27212 4684
rect 29092 4700 29144 4752
rect 29736 4743 29788 4752
rect 29736 4709 29745 4743
rect 29745 4709 29779 4743
rect 29779 4709 29788 4743
rect 29736 4700 29788 4709
rect 31484 4700 31536 4752
rect 30472 4632 30524 4684
rect 32588 4675 32640 4684
rect 32588 4641 32597 4675
rect 32597 4641 32631 4675
rect 32631 4641 32640 4675
rect 32588 4632 32640 4641
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 19248 4564 19300 4616
rect 29920 4564 29972 4616
rect 25228 4496 25280 4548
rect 26332 4496 26384 4548
rect 27620 4539 27672 4548
rect 27620 4505 27629 4539
rect 27629 4505 27663 4539
rect 27663 4505 27672 4539
rect 27620 4496 27672 4505
rect 21456 4428 21508 4480
rect 25320 4428 25372 4480
rect 29368 4428 29420 4480
rect 30748 4496 30800 4548
rect 31760 4564 31812 4616
rect 32680 4607 32732 4616
rect 32680 4573 32689 4607
rect 32689 4573 32723 4607
rect 32723 4573 32732 4607
rect 32680 4564 32732 4573
rect 33508 4564 33560 4616
rect 33784 4564 33836 4616
rect 35900 4564 35952 4616
rect 31484 4428 31536 4480
rect 32036 4471 32088 4480
rect 32036 4437 32045 4471
rect 32045 4437 32079 4471
rect 32079 4437 32088 4471
rect 32036 4428 32088 4437
rect 33232 4539 33284 4548
rect 33232 4505 33241 4539
rect 33241 4505 33275 4539
rect 33275 4505 33284 4539
rect 33232 4496 33284 4505
rect 33324 4428 33376 4480
rect 33876 4471 33928 4480
rect 33876 4437 33885 4471
rect 33885 4437 33919 4471
rect 33919 4437 33928 4471
rect 33876 4428 33928 4437
rect 36268 4471 36320 4480
rect 36268 4437 36277 4471
rect 36277 4437 36311 4471
rect 36311 4437 36320 4471
rect 36268 4428 36320 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 13544 4224 13596 4276
rect 20812 4224 20864 4276
rect 17684 4088 17736 4140
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 18972 4131 19024 4140
rect 17868 4088 17920 4097
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 21456 4156 21508 4208
rect 22376 4156 22428 4208
rect 32680 4224 32732 4276
rect 32864 4224 32916 4276
rect 25320 4156 25372 4208
rect 28448 4156 28500 4208
rect 29000 4156 29052 4208
rect 34704 4156 34756 4208
rect 19064 4088 19116 4097
rect 26056 4131 26108 4140
rect 26056 4097 26065 4131
rect 26065 4097 26099 4131
rect 26099 4097 26108 4131
rect 26056 4088 26108 4097
rect 26608 4088 26660 4140
rect 14188 4063 14240 4072
rect 14188 4029 14197 4063
rect 14197 4029 14231 4063
rect 14231 4029 14240 4063
rect 14188 4020 14240 4029
rect 17960 3884 18012 3936
rect 21640 3884 21692 3936
rect 22836 4020 22888 4072
rect 22928 4020 22980 4072
rect 23480 3952 23532 4004
rect 26240 4020 26292 4072
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 31208 4088 31260 4140
rect 28448 4020 28500 4072
rect 28908 4063 28960 4072
rect 28908 4029 28917 4063
rect 28917 4029 28951 4063
rect 28951 4029 28960 4063
rect 28908 4020 28960 4029
rect 29184 4063 29236 4072
rect 29184 4029 29193 4063
rect 29193 4029 29227 4063
rect 29227 4029 29236 4063
rect 29644 4063 29696 4072
rect 29184 4020 29236 4029
rect 29644 4029 29653 4063
rect 29653 4029 29687 4063
rect 29687 4029 29696 4063
rect 29644 4020 29696 4029
rect 31576 4020 31628 4072
rect 32312 4088 32364 4140
rect 32864 4088 32916 4140
rect 33048 4131 33100 4140
rect 33048 4097 33057 4131
rect 33057 4097 33091 4131
rect 33091 4097 33100 4131
rect 33048 4088 33100 4097
rect 33324 4088 33376 4140
rect 33784 4131 33836 4140
rect 33784 4097 33793 4131
rect 33793 4097 33827 4131
rect 33827 4097 33836 4131
rect 33784 4088 33836 4097
rect 34704 4020 34756 4072
rect 23756 3884 23808 3936
rect 24308 3884 24360 3936
rect 24400 3884 24452 3936
rect 29644 3884 29696 3936
rect 32036 3952 32088 4004
rect 35992 3952 36044 4004
rect 31208 3884 31260 3936
rect 33692 3927 33744 3936
rect 33692 3893 33701 3927
rect 33701 3893 33735 3927
rect 33735 3893 33744 3927
rect 33692 3884 33744 3893
rect 33784 3884 33836 3936
rect 35440 3927 35492 3936
rect 35440 3893 35449 3927
rect 35449 3893 35483 3927
rect 35483 3893 35492 3927
rect 35440 3884 35492 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 13544 3680 13596 3732
rect 20812 3680 20864 3732
rect 22560 3612 22612 3664
rect 29184 3680 29236 3732
rect 31392 3680 31444 3732
rect 15200 3544 15252 3596
rect 17684 3544 17736 3596
rect 20536 3544 20588 3596
rect 20812 3544 20864 3596
rect 21640 3544 21692 3596
rect 23848 3544 23900 3596
rect 24124 3544 24176 3596
rect 24400 3476 24452 3528
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 14188 3408 14240 3460
rect 17960 3340 18012 3392
rect 20720 3408 20772 3460
rect 24860 3544 24912 3596
rect 26056 3544 26108 3596
rect 26792 3587 26844 3596
rect 26792 3553 26801 3587
rect 26801 3553 26835 3587
rect 26835 3553 26844 3587
rect 26792 3544 26844 3553
rect 30104 3612 30156 3664
rect 32496 3680 32548 3732
rect 32680 3723 32732 3732
rect 32680 3689 32689 3723
rect 32689 3689 32723 3723
rect 32723 3689 32732 3723
rect 32680 3680 32732 3689
rect 34704 3680 34756 3732
rect 31576 3612 31628 3664
rect 35348 3612 35400 3664
rect 32036 3544 32088 3596
rect 33508 3544 33560 3596
rect 28448 3476 28500 3528
rect 29920 3476 29972 3528
rect 31760 3476 31812 3528
rect 33232 3476 33284 3528
rect 33324 3476 33376 3528
rect 35440 3544 35492 3596
rect 36176 3476 36228 3528
rect 27068 3451 27120 3460
rect 27068 3417 27077 3451
rect 27077 3417 27111 3451
rect 27111 3417 27120 3451
rect 27068 3408 27120 3417
rect 26148 3340 26200 3392
rect 26240 3340 26292 3392
rect 26424 3340 26476 3392
rect 27712 3340 27764 3392
rect 28540 3383 28592 3392
rect 28540 3349 28549 3383
rect 28549 3349 28583 3383
rect 28583 3349 28592 3383
rect 28540 3340 28592 3349
rect 28908 3340 28960 3392
rect 30932 3408 30984 3460
rect 31116 3408 31168 3460
rect 32036 3383 32088 3392
rect 32036 3349 32045 3383
rect 32045 3349 32079 3383
rect 32079 3349 32088 3383
rect 32036 3340 32088 3349
rect 35992 3340 36044 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 15200 3136 15252 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 17776 3136 17828 3188
rect 23572 3136 23624 3188
rect 15292 3068 15344 3120
rect 20904 3068 20956 3120
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 16948 3000 17000 3052
rect 24860 3136 24912 3188
rect 26148 3136 26200 3188
rect 31576 3136 31628 3188
rect 31668 3136 31720 3188
rect 32036 3136 32088 3188
rect 32496 3136 32548 3188
rect 25872 3111 25924 3120
rect 23112 3000 23164 3052
rect 23756 3000 23808 3052
rect 25872 3077 25881 3111
rect 25881 3077 25915 3111
rect 25915 3077 25924 3111
rect 25872 3068 25924 3077
rect 26424 3111 26476 3120
rect 26424 3077 26433 3111
rect 26433 3077 26467 3111
rect 26467 3077 26476 3111
rect 26424 3068 26476 3077
rect 26700 3068 26752 3120
rect 29736 3068 29788 3120
rect 33692 3068 33744 3120
rect 34796 3068 34848 3120
rect 35348 3068 35400 3120
rect 19064 2932 19116 2984
rect 21180 2975 21232 2984
rect 21180 2941 21189 2975
rect 21189 2941 21223 2975
rect 21223 2941 21232 2975
rect 21180 2932 21232 2941
rect 12440 2864 12492 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 4620 2796 4672 2848
rect 14096 2839 14148 2848
rect 14096 2805 14105 2839
rect 14105 2805 14139 2839
rect 14139 2805 14148 2839
rect 14096 2796 14148 2805
rect 19248 2796 19300 2848
rect 29184 3000 29236 3052
rect 29368 3043 29420 3052
rect 29368 3009 29377 3043
rect 29377 3009 29411 3043
rect 29411 3009 29420 3043
rect 29368 3000 29420 3009
rect 31484 3000 31536 3052
rect 31760 3043 31812 3052
rect 31760 3009 31769 3043
rect 31769 3009 31803 3043
rect 31803 3009 31812 3043
rect 32312 3043 32364 3052
rect 31760 3000 31812 3009
rect 32312 3009 32321 3043
rect 32321 3009 32355 3043
rect 32355 3009 32364 3043
rect 32312 3000 32364 3009
rect 33232 3043 33284 3052
rect 33232 3009 33241 3043
rect 33241 3009 33275 3043
rect 33275 3009 33284 3043
rect 33232 3000 33284 3009
rect 36084 3043 36136 3052
rect 36084 3009 36093 3043
rect 36093 3009 36127 3043
rect 36127 3009 36136 3043
rect 36084 3000 36136 3009
rect 22560 2796 22612 2848
rect 29000 2932 29052 2984
rect 29736 2932 29788 2984
rect 36360 2975 36412 2984
rect 36360 2941 36369 2975
rect 36369 2941 36403 2975
rect 36403 2941 36412 2975
rect 36360 2932 36412 2941
rect 28908 2864 28960 2916
rect 29092 2796 29144 2848
rect 29644 2796 29696 2848
rect 34796 2907 34848 2916
rect 34796 2873 34805 2907
rect 34805 2873 34839 2907
rect 34839 2873 34848 2907
rect 34796 2864 34848 2873
rect 31116 2839 31168 2848
rect 31116 2805 31125 2839
rect 31125 2805 31159 2839
rect 31159 2805 31168 2839
rect 31116 2796 31168 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1952 2592 2004 2644
rect 4712 2635 4764 2644
rect 4712 2601 4721 2635
rect 4721 2601 4755 2635
rect 4755 2601 4764 2635
rect 4712 2592 4764 2601
rect 19064 2592 19116 2644
rect 21272 2592 21324 2644
rect 25964 2592 26016 2644
rect 26792 2592 26844 2644
rect 13268 2524 13320 2576
rect 16948 2524 17000 2576
rect 28356 2592 28408 2644
rect 29276 2592 29328 2644
rect 29552 2592 29604 2644
rect 34612 2592 34664 2644
rect 35992 2592 36044 2644
rect 4620 2456 4672 2508
rect 20 2320 72 2372
rect 4712 2388 4764 2440
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 14096 2456 14148 2508
rect 12440 2388 12492 2440
rect 17684 2456 17736 2508
rect 17408 2388 17460 2440
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 5172 2252 5224 2304
rect 6460 2252 6512 2304
rect 8392 2252 8444 2304
rect 10324 2320 10376 2372
rect 18696 2388 18748 2440
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10600 2252 10652 2261
rect 11612 2252 11664 2304
rect 13544 2252 13596 2304
rect 15476 2252 15528 2304
rect 17408 2252 17460 2304
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 20628 2252 20680 2304
rect 22284 2456 22336 2508
rect 23756 2499 23808 2508
rect 23756 2465 23765 2499
rect 23765 2465 23799 2499
rect 23799 2465 23808 2499
rect 23756 2456 23808 2465
rect 24860 2499 24912 2508
rect 24860 2465 24869 2499
rect 24869 2465 24903 2499
rect 24903 2465 24912 2499
rect 24860 2456 24912 2465
rect 24952 2456 25004 2508
rect 28632 2524 28684 2576
rect 26332 2499 26384 2508
rect 26332 2465 26341 2499
rect 26341 2465 26375 2499
rect 26375 2465 26384 2499
rect 26332 2456 26384 2465
rect 26792 2456 26844 2508
rect 29460 2456 29512 2508
rect 29552 2388 29604 2440
rect 32772 2524 32824 2576
rect 24952 2320 25004 2372
rect 25872 2320 25924 2372
rect 29920 2320 29972 2372
rect 31392 2388 31444 2440
rect 32128 2388 32180 2440
rect 31484 2320 31536 2372
rect 32864 2388 32916 2440
rect 34244 2388 34296 2440
rect 34796 2388 34848 2440
rect 35624 2388 35676 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 18328 2048 18380 2100
rect 25596 2048 25648 2100
rect 20536 1980 20588 2032
rect 31484 2048 31536 2100
rect 29920 1980 29972 2032
rect 33140 1980 33192 2032
rect 10600 1912 10652 1964
rect 25044 1912 25096 1964
rect 25872 1912 25924 1964
rect 33876 1912 33928 1964
rect 28356 1844 28408 1896
rect 31208 1844 31260 1896
<< metal2 >>
rect 18 39200 74 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 14186 39200 14242 39800
rect 16118 39200 16174 39800
rect 17406 39200 17462 39800
rect 19338 39200 19394 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 26422 39200 26478 39800
rect 28354 39200 28410 39800
rect 29642 39200 29698 39800
rect 31574 39200 31630 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 32 37466 60 39200
rect 20 37460 72 37466
rect 20 37402 72 37408
rect 1964 37262 1992 39200
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 1964 36922 1992 37198
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 1952 36916 2004 36922
rect 1952 36858 2004 36864
rect 1688 36825 1716 36858
rect 1674 36816 1730 36825
rect 1674 36751 1730 36760
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1676 34944 1728 34950
rect 1676 34886 1728 34892
rect 1688 34785 1716 34886
rect 1674 34776 1730 34785
rect 1674 34711 1730 34720
rect 1676 32836 1728 32842
rect 1676 32778 1728 32784
rect 1688 32745 1716 32778
rect 1674 32736 1730 32745
rect 1674 32671 1730 32680
rect 1688 32570 1716 32671
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1676 31680 1728 31686
rect 1676 31622 1728 31628
rect 1688 31385 1716 31622
rect 1674 31376 1730 31385
rect 1674 31311 1730 31320
rect 1780 30938 1808 36722
rect 2792 36378 2820 38111
rect 3056 37256 3108 37262
rect 3056 37198 3108 37204
rect 3068 36922 3096 37198
rect 3896 37126 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5184 37262 5212 39200
rect 7116 37330 7144 39200
rect 5540 37324 5592 37330
rect 5540 37266 5592 37272
rect 7104 37324 7156 37330
rect 7104 37266 7156 37272
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3056 36916 3108 36922
rect 3056 36858 3108 36864
rect 2780 36372 2832 36378
rect 2780 36314 2832 36320
rect 2688 35080 2740 35086
rect 2688 35022 2740 35028
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1872 31482 1900 31758
rect 1860 31476 1912 31482
rect 1860 31418 1912 31424
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1768 30932 1820 30938
rect 1768 30874 1820 30880
rect 1860 30728 1912 30734
rect 1860 30670 1912 30676
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29345 1716 29446
rect 1674 29336 1730 29345
rect 1674 29271 1730 29280
rect 1676 27328 1728 27334
rect 1674 27296 1676 27305
rect 1728 27296 1730 27305
rect 1674 27231 1730 27240
rect 1872 25294 1900 30670
rect 1952 29640 2004 29646
rect 1952 29582 2004 29588
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1860 25288 1912 25294
rect 1636 25256 1638 25265
rect 1860 25230 1912 25236
rect 1582 25191 1638 25200
rect 1596 24954 1624 25191
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 1596 23905 1624 24142
rect 1582 23896 1638 23905
rect 1582 23831 1584 23840
rect 1636 23831 1638 23840
rect 1584 23802 1636 23808
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21865 1624 21966
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 1596 21690 1624 21791
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1872 20942 1900 25230
rect 1964 23594 1992 29582
rect 1952 23588 2004 23594
rect 1952 23530 2004 23536
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1584 19848 1636 19854
rect 1582 19816 1584 19825
rect 1636 19816 1638 19825
rect 1582 19751 1638 19760
rect 1596 19514 1624 19751
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1584 18692 1636 18698
rect 1584 18634 1636 18640
rect 1596 18465 1624 18634
rect 1582 18456 1638 18465
rect 1582 18391 1584 18400
rect 1636 18391 1638 18400
rect 1584 18362 1636 18368
rect 1676 16448 1728 16454
rect 1674 16416 1676 16425
rect 1728 16416 1730 16425
rect 1674 16351 1730 16360
rect 1860 14408 1912 14414
rect 1674 14376 1730 14385
rect 1860 14350 1912 14356
rect 1674 14311 1730 14320
rect 1688 14278 1716 14311
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1872 12986 1900 14350
rect 2056 14346 2084 31282
rect 2700 29850 2728 35022
rect 3988 32026 4016 37198
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3976 32020 4028 32026
rect 3976 31962 4028 31968
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 3712 23322 3740 27406
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24206 4660 31758
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3700 23316 3752 23322
rect 3700 23258 3752 23264
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2044 14340 2096 14346
rect 2044 14282 2096 14288
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 11150 1900 12038
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1676 11008 1728 11014
rect 1674 10976 1676 10985
rect 1728 10976 1730 10985
rect 1674 10911 1730 10920
rect 1674 8936 1730 8945
rect 1674 8871 1730 8880
rect 1688 8838 1716 8871
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6905 1716 7142
rect 1674 6896 1730 6905
rect 1674 6831 1730 6840
rect 1872 6458 1900 7346
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1964 6322 1992 6734
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1676 5568 1728 5574
rect 1674 5536 1676 5545
rect 1728 5536 1730 5545
rect 1674 5471 1730 5480
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 1964 2650 1992 6258
rect 2332 5914 2360 21286
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21010 4660 24142
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2700 12986 2728 18634
rect 5552 18086 5580 37266
rect 9048 37262 9076 39200
rect 10336 37330 10364 39200
rect 12268 37346 12296 39200
rect 13544 37460 13596 37466
rect 13544 37402 13596 37408
rect 10324 37324 10376 37330
rect 12268 37318 12480 37346
rect 10324 37266 10376 37272
rect 12452 37262 12480 37318
rect 7472 37256 7524 37262
rect 7472 37198 7524 37204
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 10876 37256 10928 37262
rect 10876 37198 10928 37204
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 7484 36786 7512 37198
rect 8944 37188 8996 37194
rect 8944 37130 8996 37136
rect 7472 36780 7524 36786
rect 7472 36722 7524 36728
rect 6092 29640 6144 29646
rect 6092 29582 6144 29588
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2332 5710 2360 5850
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 4632 2514 4660 2790
rect 4724 2650 4752 15302
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4724 2446 4752 2586
rect 5552 2446 5580 11494
rect 5644 10266 5672 12854
rect 6104 10538 6132 29582
rect 8956 23866 8984 37130
rect 10888 36854 10916 37198
rect 10876 36848 10928 36854
rect 10876 36790 10928 36796
rect 11060 36780 11112 36786
rect 11060 36722 11112 36728
rect 11072 29646 11100 36722
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12728 23526 12756 23666
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 6564 9178 6592 23462
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9232 16182 9260 20742
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16250 11744 16526
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 12728 12434 12756 23462
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 12728 12406 12848 12434
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11830 8156 12174
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 12820 9654 12848 12406
rect 13280 12238 13308 22918
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 12102 13308 12174
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12452 2446 12480 2858
rect 13280 2582 13308 12038
rect 13556 5234 13584 37402
rect 14200 37262 14228 39200
rect 16132 37466 16160 39200
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 16132 37330 16160 37402
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 17040 37324 17092 37330
rect 17040 37266 17092 37272
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 14464 37120 14516 37126
rect 14464 37062 14516 37068
rect 14476 12374 14504 37062
rect 17052 14074 17080 37266
rect 17420 37262 17448 39200
rect 17408 37256 17460 37262
rect 17408 37198 17460 37204
rect 18880 37256 18932 37262
rect 18880 37198 18932 37204
rect 18892 36922 18920 37198
rect 19352 37126 19380 39200
rect 21284 37466 21312 39200
rect 21272 37460 21324 37466
rect 21272 37402 21324 37408
rect 22572 37262 22600 39200
rect 22652 37324 22704 37330
rect 22652 37266 22704 37272
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 19248 37120 19300 37126
rect 19248 37062 19300 37068
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 18880 36916 18932 36922
rect 18880 36858 18932 36864
rect 19260 36854 19288 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19248 36848 19300 36854
rect 19248 36790 19300 36796
rect 17592 36780 17644 36786
rect 17592 36722 17644 36728
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 17604 36106 17632 36722
rect 17592 36100 17644 36106
rect 17592 36042 17644 36048
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 17236 16250 17264 29446
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17880 15026 17908 32710
rect 19444 31346 19472 36722
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 17052 11830 17080 14010
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13556 4622 13584 5170
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 4282 13584 4558
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13556 3738 13584 4218
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 14200 3466 14228 4014
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 15212 3194 15240 3538
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15304 3126 15332 5034
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14844 2961 14872 2994
rect 16684 2961 16712 5510
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16776 4826 16804 5238
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17236 3505 17264 8910
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17328 4690 17356 5102
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16960 3058 16988 3130
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 14830 2952 14886 2961
rect 14830 2887 14886 2896
rect 16670 2952 16726 2961
rect 16670 2887 16726 2896
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 14108 2514 14136 2790
rect 16960 2582 16988 2994
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 17420 2446 17448 14758
rect 17880 14618 17908 14962
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17972 14074 18000 20810
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19352 15706 19380 16186
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19352 15570 19380 15642
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 15026 19104 15438
rect 19352 15026 19380 15506
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18524 14482 18552 14894
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17972 13870 18000 14010
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 17972 13530 18000 13806
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17696 12442 17724 12786
rect 18248 12782 18276 13670
rect 18340 13326 18368 13670
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18340 12918 18368 13262
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18800 12850 18828 13806
rect 18984 13530 19012 13806
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 18248 12374 18276 12718
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17512 11354 17540 12038
rect 17604 11898 17632 12106
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 9110 17632 11086
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17604 6798 17632 9046
rect 17788 8634 17816 12174
rect 18064 11762 18092 12242
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18156 11898 18184 12174
rect 19076 12170 19104 14962
rect 19996 14958 20024 31078
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21376 17882 21404 19790
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 17134 20944 17478
rect 21376 17202 21404 17818
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19352 14006 19380 14214
rect 19444 14074 19472 14214
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19352 13394 19380 13942
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12850 19196 13126
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19352 12646 19380 13194
rect 19444 12986 19472 14010
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18156 11354 18184 11630
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18524 11150 18552 12106
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 19338 11792 19394 11801
rect 18800 11354 18828 11766
rect 19338 11727 19394 11736
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18892 11354 18920 11562
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18972 11280 19024 11286
rect 18800 11228 18972 11234
rect 18800 11222 19024 11228
rect 18800 11206 19012 11222
rect 19064 11212 19116 11218
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18064 10810 18092 11086
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17880 9926 17908 10610
rect 18156 10266 18184 10678
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 18800 9518 18828 11206
rect 19064 11154 19116 11160
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 9586 19012 10406
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18432 9042 18460 9318
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17788 8498 17816 8570
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17512 6390 17540 6734
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17972 5914 18000 8910
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18248 6866 18276 7414
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18524 6662 18552 8366
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18616 6458 18644 7210
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 5914 18644 6190
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18708 5778 18736 6258
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17604 2774 17632 5034
rect 17788 4758 17816 5646
rect 18800 5574 18828 9454
rect 19076 9382 19104 11154
rect 19352 11150 19380 11727
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19260 10742 19288 11018
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19076 7478 19104 7686
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18984 6322 19012 6666
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 3602 17724 4082
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17788 3194 17816 4694
rect 17880 4146 17908 5510
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17972 3942 18000 5102
rect 18984 4146 19012 6258
rect 19168 5370 19196 9590
rect 19260 8974 19288 10406
rect 19352 10266 19380 10950
rect 19444 10606 19472 12922
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 12374 20024 12582
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19628 12102 19656 12174
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11642 20024 12310
rect 20088 11801 20116 15982
rect 20180 15026 20208 16390
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20548 15162 20576 15982
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20732 15026 20760 16594
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15416 20852 15846
rect 20904 15428 20956 15434
rect 20824 15388 20904 15416
rect 20904 15370 20956 15376
rect 21008 15026 21036 16934
rect 21376 16658 21404 16934
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15094 21128 15846
rect 21652 15706 21680 17070
rect 22020 16590 22048 18022
rect 22008 16584 22060 16590
rect 21836 16532 22008 16538
rect 21836 16526 22060 16532
rect 21836 16522 22048 16526
rect 22664 16522 22692 37266
rect 24504 37262 24532 39200
rect 25504 37392 25556 37398
rect 25504 37334 25556 37340
rect 24860 37324 24912 37330
rect 24860 37266 24912 37272
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 23204 37188 23256 37194
rect 23204 37130 23256 37136
rect 23216 36786 23244 37130
rect 24504 36922 24532 37198
rect 24492 36916 24544 36922
rect 24492 36858 24544 36864
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 23400 31482 23428 36722
rect 24872 35894 24900 37266
rect 24872 35866 24992 35894
rect 23388 31476 23440 31482
rect 23388 31418 23440 31424
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22848 17202 22876 18022
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 21824 16516 22048 16522
rect 21876 16510 22048 16516
rect 22100 16516 22152 16522
rect 21824 16458 21876 16464
rect 22100 16458 22152 16464
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21100 14482 21128 15030
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20180 12918 20208 13194
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20074 11792 20130 11801
rect 20074 11727 20130 11736
rect 19996 11614 20116 11642
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19338 10160 19394 10169
rect 19338 10095 19340 10104
rect 19392 10095 19394 10104
rect 19340 10066 19392 10072
rect 19340 9988 19392 9994
rect 19536 9976 19564 10746
rect 19996 10606 20024 11494
rect 19616 10600 19668 10606
rect 19614 10568 19616 10577
rect 19984 10600 20036 10606
rect 19668 10568 19670 10577
rect 19984 10542 20036 10548
rect 19614 10503 19670 10512
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19392 9948 19564 9976
rect 19340 9930 19392 9936
rect 19352 9042 19380 9930
rect 19628 9926 19656 10202
rect 19996 10146 20024 10542
rect 20088 10282 20116 11614
rect 20180 11218 20208 12854
rect 20352 12708 20404 12714
rect 20352 12650 20404 12656
rect 20364 11830 20392 12650
rect 20456 12238 20484 13126
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20548 11642 20576 12582
rect 20640 12442 20668 13194
rect 20732 12986 20760 14350
rect 20824 14346 20852 14418
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20718 11792 20774 11801
rect 20272 11626 20576 11642
rect 20260 11620 20576 11626
rect 20312 11614 20576 11620
rect 20260 11562 20312 11568
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20088 10254 20208 10282
rect 19996 10118 20116 10146
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19444 9178 19472 9658
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19536 8537 19564 8570
rect 19892 8560 19944 8566
rect 19522 8528 19578 8537
rect 19522 8463 19578 8472
rect 19890 8528 19892 8537
rect 19944 8528 19946 8537
rect 19890 8463 19946 8472
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7274 19288 7686
rect 19352 7478 19380 8366
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19444 7342 19472 8230
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 6798 19380 7142
rect 19444 7002 19472 7278
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 19628 5642 19656 6122
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 5370 20024 9930
rect 20088 9722 20116 10118
rect 20180 9926 20208 10254
rect 20272 9926 20300 11562
rect 20352 11552 20404 11558
rect 20640 11506 20668 11766
rect 20718 11727 20774 11736
rect 20352 11494 20404 11500
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 20088 5302 20116 8978
rect 20272 7342 20300 9114
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6390 20300 6598
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20364 5710 20392 11494
rect 20548 11478 20668 11506
rect 20548 11082 20576 11478
rect 20732 11370 20760 11727
rect 20640 11342 20760 11370
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20442 10568 20498 10577
rect 20442 10503 20498 10512
rect 20456 9178 20484 10503
rect 20548 9994 20576 11018
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20548 7546 20576 9930
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 7426 20668 11342
rect 20824 10606 20852 14282
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21192 12850 21220 13738
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21192 12442 21220 12786
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21454 12200 21510 12209
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20456 7398 20668 7426
rect 20456 6118 20484 7398
rect 20732 7342 20760 9658
rect 21008 8838 21036 11698
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 20824 7886 20852 8774
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20916 7954 20944 8570
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20640 6866 20668 7278
rect 20824 7188 20852 7822
rect 20732 7160 20852 7188
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20456 5642 20484 6054
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17972 3398 18000 3878
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 19076 2990 19104 4082
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 17604 2746 17724 2774
rect 17696 2514 17724 2746
rect 19076 2650 19104 2926
rect 19260 2854 19288 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2246
rect 5184 800 5212 2246
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 10336 800 10364 2314
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 10612 1970 10640 2246
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 11624 800 11652 2246
rect 13556 800 13584 2246
rect 15488 800 15516 2246
rect 17420 800 17448 2246
rect 18340 2106 18368 2246
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18708 800 18736 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20548 2038 20576 3538
rect 20732 3466 20760 7160
rect 20916 6882 20944 7890
rect 20824 6866 20944 6882
rect 20812 6860 20944 6866
rect 20864 6854 20944 6860
rect 20812 6802 20864 6808
rect 20824 6458 20852 6802
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20824 5778 20852 6394
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20824 5098 20852 5714
rect 21008 5273 21036 8434
rect 20994 5264 21050 5273
rect 20994 5199 21050 5208
rect 20812 5092 20864 5098
rect 20812 5034 20864 5040
rect 20824 4690 20852 5034
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4282 20852 4626
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20824 3738 20852 4218
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20824 3602 20852 3674
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20824 3210 20852 3538
rect 20824 3182 20944 3210
rect 20916 3126 20944 3182
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 21100 2774 21128 11494
rect 21192 8294 21220 12174
rect 21454 12135 21456 12144
rect 21508 12135 21510 12144
rect 21456 12106 21508 12112
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21270 10976 21326 10985
rect 21270 10911 21326 10920
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21192 7818 21220 8230
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21192 7206 21220 7754
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21192 5574 21220 6666
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21284 3074 21312 10911
rect 21376 9586 21404 11222
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21468 9466 21496 12106
rect 21652 10266 21680 15642
rect 21732 15428 21784 15434
rect 21732 15370 21784 15376
rect 21744 11218 21772 15370
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21836 13938 21864 14350
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21836 11558 21864 12922
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21744 10810 21772 11154
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 21928 10690 21956 16390
rect 22112 16250 22140 16458
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 22020 13938 22048 15914
rect 22112 15688 22140 16186
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22112 15660 22232 15688
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22112 14074 22140 15506
rect 22204 15366 22232 15660
rect 22468 15428 22520 15434
rect 22468 15370 22520 15376
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22190 13560 22246 13569
rect 22190 13495 22192 13504
rect 22244 13495 22246 13504
rect 22192 13466 22244 13472
rect 22204 13326 22232 13466
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22020 11286 22048 12242
rect 22204 11898 22232 12854
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 21836 10662 21956 10690
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21376 9438 21496 9466
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21376 6730 21404 9438
rect 21456 9104 21508 9110
rect 21456 9046 21508 9052
rect 21468 8294 21496 9046
rect 21560 8634 21588 9454
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21652 6866 21680 10202
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21744 9722 21772 9930
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21836 9081 21864 10662
rect 21914 9616 21970 9625
rect 21914 9551 21970 9560
rect 21928 9450 21956 9551
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 21822 9072 21878 9081
rect 22020 9042 22048 9454
rect 21822 9007 21878 9016
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21744 8362 21772 8774
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21652 4690 21680 6802
rect 21836 5137 21864 8842
rect 22020 8650 22048 8978
rect 22112 8786 22140 10950
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22204 9178 22232 10134
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22112 8758 22232 8786
rect 22020 8622 22140 8650
rect 22112 8498 22140 8622
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22098 8392 22154 8401
rect 22098 8327 22100 8336
rect 22152 8327 22154 8336
rect 22100 8298 22152 8304
rect 22006 6352 22062 6361
rect 22006 6287 22008 6296
rect 22060 6287 22062 6296
rect 22008 6258 22060 6264
rect 22112 5914 22140 8298
rect 22204 8090 22232 8758
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22296 7970 22324 14214
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 8888 22416 13670
rect 22480 13530 22508 15370
rect 22572 14618 22600 16118
rect 22848 15162 22876 17138
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23032 15026 23060 31078
rect 24964 22094 24992 35866
rect 24964 22066 25084 22094
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23124 17746 23152 18158
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 23216 17066 23244 17750
rect 23204 17060 23256 17066
rect 23204 17002 23256 17008
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22848 14618 22876 14894
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22742 14104 22798 14113
rect 22742 14039 22744 14048
rect 22796 14039 22798 14048
rect 22744 14010 22796 14016
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 22742 13560 22798 13569
rect 22468 13524 22520 13530
rect 22742 13495 22798 13504
rect 22468 13466 22520 13472
rect 22650 12744 22706 12753
rect 22650 12679 22706 12688
rect 22664 12434 22692 12679
rect 22572 12406 22692 12434
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22480 9024 22508 10066
rect 22572 9654 22600 12406
rect 22756 12356 22784 13495
rect 22940 13258 22968 13806
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22940 12374 22968 13194
rect 23216 12753 23244 17002
rect 23584 16590 23612 18566
rect 24596 18426 24624 21830
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23860 17678 23888 18022
rect 24596 17678 24624 18362
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 17270 24624 17478
rect 24584 17264 24636 17270
rect 24584 17206 24636 17212
rect 24780 16590 24808 18022
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 23492 15978 23520 16390
rect 23860 16046 23888 16390
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 23296 15972 23348 15978
rect 23296 15914 23348 15920
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23308 15570 23336 15914
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23492 14890 23520 15914
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 23584 14618 23612 15370
rect 23676 15094 23704 15846
rect 24308 15428 24360 15434
rect 24308 15370 24360 15376
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23400 14074 23428 14350
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23400 13394 23428 14010
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23492 12918 23520 13806
rect 23664 13796 23716 13802
rect 23664 13738 23716 13744
rect 23676 13462 23704 13738
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23202 12744 23258 12753
rect 23202 12679 23258 12688
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 22664 12328 22784 12356
rect 22928 12368 22980 12374
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22664 9602 22692 12328
rect 22928 12310 22980 12316
rect 23018 12336 23074 12345
rect 23018 12271 23074 12280
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22756 10606 22784 11562
rect 22940 11218 22968 12106
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 10130 22876 10406
rect 22940 10198 22968 11154
rect 23032 10606 23060 12271
rect 23216 11762 23244 12378
rect 23584 12306 23612 13194
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23492 11801 23520 12106
rect 23478 11792 23534 11801
rect 23204 11756 23256 11762
rect 23676 11762 23704 13398
rect 23768 12889 23796 13942
rect 24320 13258 24348 15370
rect 24412 14822 24440 15982
rect 24872 14958 24900 16390
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24412 14346 24440 14758
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24400 14340 24452 14346
rect 24400 14282 24452 14288
rect 24308 13252 24360 13258
rect 24308 13194 24360 13200
rect 23754 12880 23810 12889
rect 23754 12815 23810 12824
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23768 11898 23796 12718
rect 24320 12714 24348 13194
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24596 12986 24624 13126
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23478 11727 23534 11736
rect 23664 11756 23716 11762
rect 23204 11698 23256 11704
rect 23664 11698 23716 11704
rect 23216 11150 23244 11698
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 23032 10130 23060 10542
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23018 10024 23074 10033
rect 23018 9959 23074 9968
rect 22664 9574 22968 9602
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22480 8996 22600 9024
rect 22468 8900 22520 8906
rect 22388 8860 22468 8888
rect 22388 8401 22416 8860
rect 22468 8842 22520 8848
rect 22374 8392 22430 8401
rect 22374 8327 22430 8336
rect 22204 7942 22324 7970
rect 22204 7546 22232 7942
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22204 6118 22232 6394
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21822 5128 21878 5137
rect 22020 5098 22048 5306
rect 21822 5063 21878 5072
rect 22008 5092 22060 5098
rect 22008 5034 22060 5040
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21468 4214 21496 4422
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21652 3602 21680 3878
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 21192 3046 21312 3074
rect 21192 2990 21220 3046
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21008 2746 21128 2774
rect 21008 2446 21036 2746
rect 21284 2650 21312 3046
rect 22388 2774 22416 4150
rect 22572 3670 22600 8996
rect 22664 4826 22692 9454
rect 22940 9110 22968 9574
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22756 7206 22784 7686
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22848 4078 22876 7686
rect 22940 5778 22968 9046
rect 23032 8022 23060 9959
rect 23020 8016 23072 8022
rect 23020 7958 23072 7964
rect 23032 7410 23060 7958
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23032 6662 23060 7346
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 22940 4078 22968 5102
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 23124 3058 23152 10202
rect 23216 10130 23244 11086
rect 23296 10736 23348 10742
rect 23348 10684 23612 10690
rect 23296 10678 23612 10684
rect 23308 10662 23612 10678
rect 23296 10600 23348 10606
rect 23294 10568 23296 10577
rect 23348 10568 23350 10577
rect 23294 10503 23350 10512
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23216 6866 23244 10066
rect 23308 9722 23336 10406
rect 23584 9722 23612 10662
rect 23676 10606 23704 11698
rect 23768 11694 23796 11834
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23768 9466 23796 11086
rect 23860 10033 23888 12582
rect 24492 12436 24544 12442
rect 24780 12434 24808 14350
rect 24860 13932 24912 13938
rect 24964 13920 24992 15098
rect 24912 13892 24992 13920
rect 24860 13874 24912 13880
rect 24492 12378 24544 12384
rect 24596 12406 24808 12434
rect 24872 12434 24900 13874
rect 25056 13530 25084 22066
rect 25516 17678 25544 37334
rect 26436 37126 26464 39200
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 26804 26586 26832 37198
rect 28368 37126 28396 39200
rect 28816 37256 28868 37262
rect 28816 37198 28868 37204
rect 28632 37188 28684 37194
rect 28632 37130 28684 37136
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 28644 36582 28672 37130
rect 28828 36582 28856 37198
rect 29656 37126 29684 39200
rect 31588 37346 31616 39200
rect 31588 37318 31708 37346
rect 29736 37256 29788 37262
rect 29736 37198 29788 37204
rect 31680 37210 31708 37318
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29748 36650 29776 37198
rect 31680 37182 31800 37210
rect 31772 37126 31800 37182
rect 33520 37126 33548 39200
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 31760 37120 31812 37126
rect 31760 37062 31812 37068
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 29736 36644 29788 36650
rect 29736 36586 29788 36592
rect 33612 36582 33640 37198
rect 34808 36922 34836 39200
rect 35530 38856 35586 38865
rect 35530 38791 35586 38800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35544 37330 35572 38791
rect 35532 37324 35584 37330
rect 35532 37266 35584 37272
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 34796 36916 34848 36922
rect 34796 36858 34848 36864
rect 28632 36576 28684 36582
rect 28632 36518 28684 36524
rect 28816 36576 28868 36582
rect 28816 36518 28868 36524
rect 33600 36576 33652 36582
rect 33600 36518 33652 36524
rect 27436 31340 27488 31346
rect 27436 31282 27488 31288
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 27448 21894 27476 31282
rect 27620 26308 27672 26314
rect 27620 26250 27672 26256
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 25688 18148 25740 18154
rect 25688 18090 25740 18096
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25424 16794 25452 17138
rect 25412 16788 25464 16794
rect 25412 16730 25464 16736
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 25136 14884 25188 14890
rect 25136 14826 25188 14832
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 25056 13326 25084 13466
rect 25044 13320 25096 13326
rect 25148 13297 25176 14826
rect 25044 13262 25096 13268
rect 25134 13288 25190 13297
rect 25134 13223 25190 13232
rect 24872 12406 25084 12434
rect 24504 12238 24532 12378
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24030 11112 24086 11121
rect 23940 11076 23992 11082
rect 24030 11047 24032 11056
rect 23940 11018 23992 11024
rect 24084 11047 24086 11056
rect 24032 11018 24084 11024
rect 23846 10024 23902 10033
rect 23846 9959 23902 9968
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23676 9438 23796 9466
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 23400 8838 23428 9046
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23308 4593 23336 8502
rect 23478 6352 23534 6361
rect 23478 6287 23534 6296
rect 23294 4584 23350 4593
rect 23294 4519 23350 4528
rect 23492 4010 23520 6287
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23584 3194 23612 9386
rect 23676 7886 23704 9438
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 9110 23796 9318
rect 23756 9104 23808 9110
rect 23756 9046 23808 9052
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23676 6202 23704 7822
rect 23768 7478 23796 9046
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23860 7546 23888 8842
rect 23952 8090 23980 11018
rect 24136 9994 24164 11494
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 24044 7886 24072 9114
rect 24228 9042 24256 9454
rect 24320 9382 24348 11494
rect 24504 11354 24532 12174
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24492 10736 24544 10742
rect 24492 10678 24544 10684
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 24136 7954 24164 8842
rect 24228 8498 24256 8978
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24504 8090 24532 10678
rect 24596 8430 24624 12406
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 24688 11354 24716 11766
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24780 11150 24808 11290
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24780 10266 24808 10542
rect 25056 10470 25084 12406
rect 25148 11830 25176 13223
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25240 11218 25268 15506
rect 25318 15056 25374 15065
rect 25318 14991 25374 15000
rect 25332 14958 25360 14991
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25320 13252 25372 13258
rect 25320 13194 25372 13200
rect 25332 11286 25360 13194
rect 25320 11280 25372 11286
rect 25320 11222 25372 11228
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24688 9382 24716 9862
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24780 9654 24808 9687
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24950 9616 25006 9625
rect 24950 9551 25006 9560
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24044 7750 24072 7822
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 24320 7342 24348 7414
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24308 7336 24360 7342
rect 24308 7278 24360 7284
rect 24044 6866 24072 7278
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24044 6322 24072 6802
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24412 6458 24440 6598
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23676 6186 23888 6202
rect 24596 6186 24624 8366
rect 24688 7954 24716 8366
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24780 6662 24808 7822
rect 24964 6662 24992 9551
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 23676 6180 23900 6186
rect 23676 6174 23848 6180
rect 23848 6122 23900 6128
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 23860 5778 23888 6122
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 24124 5024 24176 5030
rect 24124 4966 24176 4972
rect 23676 4690 23704 4966
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23754 4040 23810 4049
rect 23754 3975 23810 3984
rect 23768 3942 23796 3975
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 24136 3602 24164 4966
rect 24308 3936 24360 3942
rect 24306 3904 24308 3913
rect 24400 3936 24452 3942
rect 24360 3904 24362 3913
rect 24400 3878 24452 3884
rect 24306 3839 24362 3848
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22296 2746 22416 2774
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 22296 2514 22324 2746
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20536 2032 20588 2038
rect 20536 1974 20588 1980
rect 20640 800 20668 2246
rect 22572 800 22600 2790
rect 23768 2514 23796 2994
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23860 800 23888 3538
rect 24412 3534 24440 3878
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24780 3097 24808 6598
rect 24964 6390 24992 6598
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24872 3194 24900 3538
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24766 3088 24822 3097
rect 24766 3023 24822 3032
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 24872 2514 24900 2751
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 24964 2378 24992 2450
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 25056 1970 25084 10406
rect 25424 9625 25452 16730
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25516 12345 25544 13806
rect 25700 12434 25728 18090
rect 26700 18080 26752 18086
rect 26700 18022 26752 18028
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 25792 16182 25820 17070
rect 25780 16176 25832 16182
rect 25780 16118 25832 16124
rect 25884 15026 25912 17478
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26252 17066 26464 17082
rect 26240 17060 26476 17066
rect 26292 17054 26424 17060
rect 26240 17002 26292 17008
rect 26424 17002 26476 17008
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 25884 14906 25912 14962
rect 25792 14878 25912 14906
rect 26068 14890 26096 16594
rect 26620 16522 26648 16934
rect 26712 16658 26740 18022
rect 27436 17264 27488 17270
rect 27436 17206 27488 17212
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 27448 16590 27476 17206
rect 27632 16794 27660 26250
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27528 16720 27580 16726
rect 27528 16662 27580 16668
rect 27436 16584 27488 16590
rect 27436 16526 27488 16532
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26608 16516 26660 16522
rect 26608 16458 26660 16464
rect 27160 16516 27212 16522
rect 27160 16458 27212 16464
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26160 16114 26188 16390
rect 26344 16114 26372 16458
rect 26792 16176 26844 16182
rect 26792 16118 26844 16124
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26516 15904 26568 15910
rect 26516 15846 26568 15852
rect 26528 15434 26556 15846
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26344 15162 26372 15370
rect 26620 15314 26648 16050
rect 26528 15286 26648 15314
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 26056 14884 26108 14890
rect 25792 14006 25820 14878
rect 26056 14826 26108 14832
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26160 14414 26188 14826
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26252 14278 26280 14758
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26252 14006 26280 14214
rect 25780 14000 25832 14006
rect 25780 13942 25832 13948
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 25976 13530 26004 13874
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25962 13424 26018 13433
rect 25780 13388 25832 13394
rect 26068 13394 26096 13466
rect 25962 13359 26018 13368
rect 26056 13388 26108 13394
rect 25780 13330 25832 13336
rect 25792 12782 25820 13330
rect 25976 13258 26004 13359
rect 26056 13330 26108 13336
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 26146 12880 26202 12889
rect 26146 12815 26148 12824
rect 26200 12815 26202 12824
rect 26148 12786 26200 12792
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 26148 12640 26200 12646
rect 25608 12406 25728 12434
rect 26068 12600 26148 12628
rect 25502 12336 25558 12345
rect 25502 12271 25558 12280
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 10266 25544 11018
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25410 9616 25466 9625
rect 25410 9551 25466 9560
rect 25228 9036 25280 9042
rect 25148 8996 25228 9024
rect 25148 8906 25176 8996
rect 25228 8978 25280 8984
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25424 7002 25452 7346
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25412 6996 25464 7002
rect 25412 6938 25464 6944
rect 25516 5574 25544 7142
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25240 4554 25268 4762
rect 25228 4548 25280 4554
rect 25228 4490 25280 4496
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25332 4214 25360 4422
rect 25320 4208 25372 4214
rect 25320 4150 25372 4156
rect 25516 2825 25544 5510
rect 25502 2816 25558 2825
rect 25502 2751 25558 2760
rect 25608 2106 25636 12406
rect 26068 11830 26096 12600
rect 26148 12582 26200 12588
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 26160 11778 26188 11834
rect 26160 11750 26280 11778
rect 25780 11620 25832 11626
rect 25780 11562 25832 11568
rect 25792 11082 25820 11562
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 25780 11076 25832 11082
rect 25780 11018 25832 11024
rect 26160 10742 26188 11154
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 26252 10266 26280 11750
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 26436 10198 26464 10474
rect 26424 10192 26476 10198
rect 26424 10134 26476 10140
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 25976 9178 26004 9318
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25976 7410 26004 8910
rect 26056 8288 26108 8294
rect 26056 8230 26108 8236
rect 26068 8090 26096 8230
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26148 7948 26200 7954
rect 26148 7890 26200 7896
rect 26160 7546 26188 7890
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 26056 6860 26108 6866
rect 26160 6848 26188 7482
rect 26528 7478 26556 15286
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26620 14346 26648 14554
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26620 13394 26648 13806
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 26608 12776 26660 12782
rect 26606 12744 26608 12753
rect 26660 12744 26662 12753
rect 26606 12679 26662 12688
rect 26804 12434 26832 16118
rect 27172 15502 27200 16458
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 26976 15428 27028 15434
rect 26976 15370 27028 15376
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26712 12406 26832 12434
rect 26516 7472 26568 7478
rect 26516 7414 26568 7420
rect 26108 6820 26188 6848
rect 26332 6860 26384 6866
rect 26056 6802 26108 6808
rect 26332 6802 26384 6808
rect 26344 6746 26372 6802
rect 26252 6730 26372 6746
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 26240 6724 26372 6730
rect 26292 6718 26372 6724
rect 26240 6666 26292 6672
rect 25700 5710 25728 6666
rect 25780 6656 25832 6662
rect 25780 6598 25832 6604
rect 25792 5794 25820 6598
rect 25792 5766 26188 5794
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25884 3126 25912 5766
rect 26160 5642 26188 5766
rect 26148 5636 26200 5642
rect 26148 5578 26200 5584
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26068 5030 26096 5510
rect 26424 5092 26476 5098
rect 26424 5034 26476 5040
rect 26056 5024 26108 5030
rect 26056 4966 26108 4972
rect 26068 4690 26096 4966
rect 26056 4684 26108 4690
rect 26056 4626 26108 4632
rect 26068 4146 26096 4626
rect 26332 4548 26384 4554
rect 26332 4490 26384 4496
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26068 3602 26096 4082
rect 26240 4072 26292 4078
rect 26240 4014 26292 4020
rect 26056 3596 26108 3602
rect 26056 3538 26108 3544
rect 26252 3398 26280 4014
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26160 3194 26188 3334
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 25964 2644 26016 2650
rect 25964 2586 26016 2592
rect 25976 2530 26004 2586
rect 25792 2502 26004 2530
rect 26344 2514 26372 4490
rect 26436 3398 26464 5034
rect 26528 4162 26556 7414
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 26620 5846 26648 6190
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26528 4146 26648 4162
rect 26528 4140 26660 4146
rect 26528 4134 26608 4140
rect 26608 4082 26660 4088
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26436 3126 26464 3334
rect 26712 3126 26740 12406
rect 26896 11762 26924 14826
rect 26988 12345 27016 15370
rect 27264 15026 27292 15846
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27356 14958 27384 16186
rect 27436 15904 27488 15910
rect 27436 15846 27488 15852
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27448 13258 27476 15846
rect 27540 15484 27568 16662
rect 27632 16114 27660 16730
rect 27816 16522 27844 17546
rect 27804 16516 27856 16522
rect 27804 16458 27856 16464
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 27988 15700 28040 15706
rect 27988 15642 28040 15648
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27612 15496 27664 15502
rect 27540 15456 27612 15484
rect 27612 15438 27664 15444
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27540 15162 27568 15302
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27632 14226 27660 15438
rect 27724 14550 27752 15506
rect 27896 15428 27948 15434
rect 27816 15388 27896 15416
rect 27712 14544 27764 14550
rect 27712 14486 27764 14492
rect 27816 14362 27844 15388
rect 27896 15370 27948 15376
rect 28000 15026 28028 15642
rect 28080 15632 28132 15638
rect 28080 15574 28132 15580
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 27724 14346 27844 14362
rect 27908 14346 27936 14554
rect 27988 14544 28040 14550
rect 27988 14486 28040 14492
rect 28000 14346 28028 14486
rect 27712 14340 27844 14346
rect 27764 14334 27844 14340
rect 27896 14340 27948 14346
rect 27712 14282 27764 14288
rect 27896 14282 27948 14288
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 27632 14198 27936 14226
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27712 13864 27764 13870
rect 27712 13806 27764 13812
rect 27528 13796 27580 13802
rect 27528 13738 27580 13744
rect 27540 13410 27568 13738
rect 27724 13433 27752 13806
rect 27710 13424 27766 13433
rect 27540 13382 27660 13410
rect 27526 13288 27582 13297
rect 27436 13252 27488 13258
rect 27526 13223 27528 13232
rect 27436 13194 27488 13200
rect 27580 13223 27582 13232
rect 27528 13194 27580 13200
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 26974 12336 27030 12345
rect 26974 12271 27030 12280
rect 27172 11898 27200 12854
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 27632 12730 27660 13382
rect 27710 13359 27766 13368
rect 27448 12434 27476 12718
rect 27632 12714 27752 12730
rect 27632 12708 27764 12714
rect 27632 12702 27712 12708
rect 27712 12650 27764 12656
rect 27264 12406 27476 12434
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 26884 11756 26936 11762
rect 26884 11698 26936 11704
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26988 10198 27016 10542
rect 26976 10192 27028 10198
rect 26976 10134 27028 10140
rect 26790 9752 26846 9761
rect 26790 9687 26846 9696
rect 26804 9654 26832 9687
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27080 3913 27108 9522
rect 27172 9382 27200 9522
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 27264 8537 27292 12406
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 27356 12102 27384 12174
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27724 11830 27752 12242
rect 27816 11898 27844 14010
rect 27908 12322 27936 14198
rect 28092 14113 28120 15574
rect 28078 14104 28134 14113
rect 28078 14039 28134 14048
rect 28184 13802 28212 16458
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28276 15065 28304 15302
rect 28262 15056 28318 15065
rect 28262 14991 28318 15000
rect 28552 14414 28580 18702
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 28184 13410 28212 13738
rect 28448 13728 28500 13734
rect 28448 13670 28500 13676
rect 28092 13382 28212 13410
rect 28460 13394 28488 13670
rect 28448 13388 28500 13394
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 28000 12442 28028 13126
rect 28092 12850 28120 13382
rect 28448 13330 28500 13336
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28184 13002 28212 13194
rect 28184 12974 28396 13002
rect 28264 12912 28316 12918
rect 28264 12854 28316 12860
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 27988 12436 28040 12442
rect 27988 12378 28040 12384
rect 28078 12336 28134 12345
rect 27908 12294 28028 12322
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 27804 11892 27856 11898
rect 27804 11834 27856 11840
rect 27712 11824 27764 11830
rect 27618 11792 27674 11801
rect 27528 11756 27580 11762
rect 27712 11766 27764 11772
rect 27618 11727 27674 11736
rect 27528 11698 27580 11704
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27250 8528 27306 8537
rect 27250 8463 27306 8472
rect 27264 7478 27292 8463
rect 27448 8362 27476 9522
rect 27540 8430 27568 11698
rect 27632 11694 27660 11727
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27724 11218 27752 11766
rect 27804 11756 27856 11762
rect 27908 11744 27936 12174
rect 27856 11716 27936 11744
rect 27804 11698 27856 11704
rect 27816 11558 27844 11698
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 27712 11212 27764 11218
rect 27712 11154 27764 11160
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27632 10470 27660 10950
rect 27724 10606 27752 11154
rect 27896 10736 27948 10742
rect 27896 10678 27948 10684
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27710 10160 27766 10169
rect 27710 10095 27766 10104
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27632 9178 27660 9998
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27356 6866 27384 7346
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27160 6112 27212 6118
rect 27160 6054 27212 6060
rect 27172 5778 27200 6054
rect 27250 5944 27306 5953
rect 27250 5879 27306 5888
rect 27264 5846 27292 5879
rect 27252 5840 27304 5846
rect 27252 5782 27304 5788
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 27172 5234 27200 5714
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 27172 4690 27200 5170
rect 27160 4684 27212 4690
rect 27160 4626 27212 4632
rect 27448 4078 27476 8298
rect 27528 6384 27580 6390
rect 27528 6326 27580 6332
rect 27540 5166 27568 6326
rect 27632 5642 27660 9114
rect 27620 5636 27672 5642
rect 27620 5578 27672 5584
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27724 4570 27752 10095
rect 27908 9654 27936 10678
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27896 7336 27948 7342
rect 28000 7290 28028 12294
rect 28078 12271 28134 12280
rect 28092 10742 28120 12271
rect 28080 10736 28132 10742
rect 28080 10678 28132 10684
rect 28276 10266 28304 12854
rect 28368 12442 28396 12974
rect 28356 12436 28408 12442
rect 28356 12378 28408 12384
rect 28552 11880 28580 14350
rect 28632 14340 28684 14346
rect 28632 14282 28684 14288
rect 28644 13530 28672 14282
rect 28736 13784 28764 14962
rect 28828 14074 28856 36518
rect 32312 36168 32364 36174
rect 32312 36110 32364 36116
rect 32324 31482 32352 36110
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29748 17678 29776 19790
rect 30392 18290 30420 24142
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 33152 20058 33180 20810
rect 33140 20052 33192 20058
rect 33140 19994 33192 20000
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29012 14414 29040 16594
rect 33612 15706 33640 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35820 35894 35848 37198
rect 36268 36916 36320 36922
rect 36268 36858 36320 36864
rect 36280 36825 36308 36858
rect 36266 36816 36322 36825
rect 35992 36780 36044 36786
rect 36266 36751 36322 36760
rect 35992 36722 36044 36728
rect 35728 35866 35848 35894
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35440 34944 35492 34950
rect 35440 34886 35492 34892
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34532 17882 34560 18702
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 33600 15700 33652 15706
rect 33600 15642 33652 15648
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 29000 14408 29052 14414
rect 29000 14350 29052 14356
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 29000 14068 29052 14074
rect 29000 14010 29052 14016
rect 28816 13796 28868 13802
rect 28736 13756 28816 13784
rect 28816 13738 28868 13744
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 28632 12232 28684 12238
rect 28630 12200 28632 12209
rect 28684 12200 28686 12209
rect 28630 12135 28686 12144
rect 28828 12102 28856 13738
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28460 11852 28580 11880
rect 28460 10538 28488 11852
rect 28540 11756 28592 11762
rect 28540 11698 28592 11704
rect 28552 11150 28580 11698
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28552 10985 28580 11086
rect 28538 10976 28594 10985
rect 28538 10911 28594 10920
rect 28632 10668 28684 10674
rect 28632 10610 28684 10616
rect 28448 10532 28500 10538
rect 28448 10474 28500 10480
rect 28264 10260 28316 10266
rect 28264 10202 28316 10208
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28184 8498 28212 9114
rect 28264 9104 28316 9110
rect 28264 9046 28316 9052
rect 28276 8566 28304 9046
rect 28264 8560 28316 8566
rect 28264 8502 28316 8508
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 27948 7284 28028 7290
rect 27896 7278 28028 7284
rect 27908 7262 28028 7278
rect 28000 6662 28028 7262
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 28092 5778 28120 6598
rect 28080 5772 28132 5778
rect 28080 5714 28132 5720
rect 27632 4554 27752 4570
rect 27620 4548 27752 4554
rect 27672 4542 27752 4548
rect 27620 4490 27672 4496
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27066 3904 27122 3913
rect 27066 3839 27122 3848
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26424 3120 26476 3126
rect 26424 3062 26476 3068
rect 26700 3120 26752 3126
rect 26700 3062 26752 3068
rect 26804 2650 26832 3538
rect 27080 3466 27108 3839
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26804 2514 26832 2586
rect 26332 2508 26384 2514
rect 25596 2100 25648 2106
rect 25596 2042 25648 2048
rect 25044 1964 25096 1970
rect 25044 1906 25096 1912
rect 25792 800 25820 2502
rect 26332 2450 26384 2456
rect 26792 2508 26844 2514
rect 26792 2450 26844 2456
rect 25872 2372 25924 2378
rect 25872 2314 25924 2320
rect 25884 1970 25912 2314
rect 25872 1964 25924 1970
rect 25872 1906 25924 1912
rect 27724 800 27752 3334
rect 28368 2650 28396 9998
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 28460 8838 28488 9318
rect 28644 8838 28672 10610
rect 28828 9500 28856 12038
rect 28920 11354 28948 13670
rect 29012 11354 29040 14010
rect 29104 13569 29132 14894
rect 30840 14884 30892 14890
rect 30840 14826 30892 14832
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29552 14408 29604 14414
rect 29552 14350 29604 14356
rect 29368 13932 29420 13938
rect 29368 13874 29420 13880
rect 29090 13560 29146 13569
rect 29090 13495 29146 13504
rect 29184 13320 29236 13326
rect 29184 13262 29236 13268
rect 29196 12782 29224 13262
rect 29184 12776 29236 12782
rect 29184 12718 29236 12724
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 29104 12442 29132 12650
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29196 11762 29224 12718
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 28908 11348 28960 11354
rect 28908 11290 28960 11296
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28736 9472 28856 9500
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28448 7200 28500 7206
rect 28448 7142 28500 7148
rect 28460 4214 28488 7142
rect 28448 4208 28500 4214
rect 28448 4150 28500 4156
rect 28448 4072 28500 4078
rect 28448 4014 28500 4020
rect 28460 3534 28488 4014
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28538 3496 28594 3505
rect 28538 3431 28594 3440
rect 28552 3398 28580 3431
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28356 2644 28408 2650
rect 28356 2586 28408 2592
rect 28368 1902 28396 2586
rect 28644 2582 28672 8774
rect 28736 8022 28764 9472
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 28736 5846 28764 7958
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 28920 7342 28948 7482
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 28724 5840 28776 5846
rect 28724 5782 28776 5788
rect 29012 5370 29040 10610
rect 29196 9602 29224 11698
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29104 9574 29224 9602
rect 29104 8090 29132 9574
rect 29184 9444 29236 9450
rect 29184 9386 29236 9392
rect 29196 9042 29224 9386
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29196 8838 29224 8978
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29092 8084 29144 8090
rect 29092 8026 29144 8032
rect 29196 7954 29224 8774
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 29196 7750 29224 7890
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 29196 7342 29224 7686
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29196 6662 29224 7278
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 29288 6254 29316 10542
rect 29380 9178 29408 13874
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29368 6928 29420 6934
rect 29368 6870 29420 6876
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 29184 6112 29236 6118
rect 29184 6054 29236 6060
rect 29090 5944 29146 5953
rect 29090 5879 29092 5888
rect 29144 5879 29146 5888
rect 29092 5850 29144 5856
rect 29000 5364 29052 5370
rect 29000 5306 29052 5312
rect 29012 4214 29040 5306
rect 29092 5228 29144 5234
rect 29092 5170 29144 5176
rect 29104 5030 29132 5170
rect 29196 5166 29224 6054
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 29000 4208 29052 4214
rect 29000 4150 29052 4156
rect 28908 4072 28960 4078
rect 29104 4026 29132 4694
rect 28960 4020 29132 4026
rect 28908 4014 29132 4020
rect 29184 4072 29236 4078
rect 29184 4014 29236 4020
rect 28920 3998 29132 4014
rect 29196 3738 29224 4014
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29090 3632 29146 3641
rect 29090 3567 29146 3576
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 2922 28948 3334
rect 28998 3088 29054 3097
rect 28998 3023 29054 3032
rect 29012 2990 29040 3023
rect 29000 2984 29052 2990
rect 29000 2926 29052 2932
rect 28908 2916 28960 2922
rect 28908 2858 28960 2864
rect 29104 2854 29132 3567
rect 29196 3058 29224 3674
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 29288 2650 29316 6190
rect 29380 4486 29408 6870
rect 29368 4480 29420 4486
rect 29368 4422 29420 4428
rect 29472 3924 29500 9998
rect 29564 6934 29592 14350
rect 29736 14272 29788 14278
rect 29736 14214 29788 14220
rect 29748 14074 29776 14214
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29828 12164 29880 12170
rect 29828 12106 29880 12112
rect 29840 11898 29868 12106
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29552 6928 29604 6934
rect 29552 6870 29604 6876
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29564 6118 29592 6598
rect 29656 6186 29684 7822
rect 29644 6180 29696 6186
rect 29644 6122 29696 6128
rect 29552 6112 29604 6118
rect 29604 6060 29684 6066
rect 29552 6054 29684 6060
rect 29564 6038 29684 6054
rect 29656 5710 29684 6038
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29656 5030 29684 5646
rect 29644 5024 29696 5030
rect 29644 4966 29696 4972
rect 29656 4078 29684 4966
rect 29748 4758 29776 11698
rect 30024 10810 30052 14486
rect 30852 14074 30880 14826
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 33428 13938 33456 15438
rect 34624 14278 34652 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18970 35388 26318
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34612 14272 34664 14278
rect 34612 14214 34664 14220
rect 33416 13932 33468 13938
rect 33416 13874 33468 13880
rect 30104 11144 30156 11150
rect 30104 11086 30156 11092
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 29840 5030 29868 5510
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29736 4752 29788 4758
rect 29736 4694 29788 4700
rect 29932 4622 29960 7822
rect 30116 5234 30144 11086
rect 31484 11076 31536 11082
rect 31484 11018 31536 11024
rect 31024 9648 31076 9654
rect 31024 9590 31076 9596
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30300 7750 30328 8298
rect 30288 7744 30340 7750
rect 30288 7686 30340 7692
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30392 5302 30420 6394
rect 30484 6254 30512 8842
rect 30932 7268 30984 7274
rect 30932 7210 30984 7216
rect 30748 6656 30800 6662
rect 30748 6598 30800 6604
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30472 6112 30524 6118
rect 30576 6066 30604 6258
rect 30524 6060 30604 6066
rect 30472 6054 30604 6060
rect 30484 6038 30604 6054
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 30484 5234 30512 6038
rect 30760 5302 30788 6598
rect 30564 5296 30616 5302
rect 30564 5238 30616 5244
rect 30748 5296 30800 5302
rect 30748 5238 30800 5244
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29656 3942 29684 4014
rect 29644 3936 29696 3942
rect 29472 3896 29592 3924
rect 29368 3052 29420 3058
rect 29420 3012 29500 3040
rect 29368 2994 29420 3000
rect 29276 2644 29328 2650
rect 29276 2586 29328 2592
rect 28632 2576 28684 2582
rect 28632 2518 28684 2524
rect 29472 2514 29500 3012
rect 29564 2650 29592 3896
rect 29644 3878 29696 3884
rect 30116 3670 30144 5170
rect 30484 4690 30512 5170
rect 30472 4684 30524 4690
rect 30472 4626 30524 4632
rect 30576 4049 30604 5238
rect 30748 5160 30800 5166
rect 30748 5102 30800 5108
rect 30760 4554 30788 5102
rect 30748 4548 30800 4554
rect 30748 4490 30800 4496
rect 30562 4040 30618 4049
rect 30562 3975 30618 3984
rect 30104 3664 30156 3670
rect 30104 3606 30156 3612
rect 29920 3528 29972 3534
rect 29918 3496 29920 3505
rect 29972 3496 29974 3505
rect 30944 3466 30972 7210
rect 31036 5846 31064 9590
rect 31392 9104 31444 9110
rect 31392 9046 31444 9052
rect 31208 8084 31260 8090
rect 31208 8026 31260 8032
rect 31220 7410 31248 8026
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31116 6656 31168 6662
rect 31116 6598 31168 6604
rect 31024 5840 31076 5846
rect 31024 5782 31076 5788
rect 31128 5710 31156 6598
rect 31404 6458 31432 9046
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 31496 5914 31524 11018
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32312 9444 32364 9450
rect 32312 9386 32364 9392
rect 32324 9178 32352 9386
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32324 8566 32352 9114
rect 31576 8560 31628 8566
rect 31576 8502 31628 8508
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 31588 6118 31616 8502
rect 31760 8356 31812 8362
rect 31760 8298 31812 8304
rect 31772 7478 31800 8298
rect 31864 8090 31892 8502
rect 32324 8106 32352 8502
rect 31852 8084 31904 8090
rect 32324 8078 32444 8106
rect 31852 8026 31904 8032
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 32036 7744 32088 7750
rect 32036 7686 32088 7692
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 31772 7262 31984 7290
rect 31576 6112 31628 6118
rect 31576 6054 31628 6060
rect 31484 5908 31536 5914
rect 31484 5850 31536 5856
rect 31116 5704 31168 5710
rect 31116 5646 31168 5652
rect 31496 4758 31524 5850
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 31680 5302 31708 5646
rect 31772 5574 31800 7262
rect 31956 7206 31984 7262
rect 31852 7200 31904 7206
rect 31852 7142 31904 7148
rect 31944 7200 31996 7206
rect 31944 7142 31996 7148
rect 31864 6798 31892 7142
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 31864 6322 31892 6734
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 32048 5914 32076 7686
rect 32036 5908 32088 5914
rect 32036 5850 32088 5856
rect 31760 5568 31812 5574
rect 31760 5510 31812 5516
rect 31668 5296 31720 5302
rect 31668 5238 31720 5244
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 31484 4752 31536 4758
rect 31484 4694 31536 4700
rect 31772 4622 31800 5170
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 31484 4480 31536 4486
rect 31484 4422 31536 4428
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31220 4026 31248 4082
rect 31128 3998 31248 4026
rect 31128 3505 31156 3998
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31114 3496 31170 3505
rect 29918 3431 29974 3440
rect 30932 3460 30984 3466
rect 31114 3431 31116 3440
rect 30932 3402 30984 3408
rect 31168 3431 31170 3440
rect 31116 3402 31168 3408
rect 29736 3120 29788 3126
rect 29736 3062 29788 3068
rect 29748 2990 29776 3062
rect 29736 2984 29788 2990
rect 29736 2926 29788 2932
rect 29644 2848 29696 2854
rect 31116 2848 31168 2854
rect 29644 2790 29696 2796
rect 31114 2816 31116 2825
rect 31168 2816 31170 2825
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 29460 2508 29512 2514
rect 29460 2450 29512 2456
rect 29564 2446 29592 2586
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 28356 1896 28408 1902
rect 28356 1838 28408 1844
rect 29656 800 29684 2790
rect 31114 2751 31170 2760
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 2038 29960 2314
rect 29920 2032 29972 2038
rect 29920 1974 29972 1980
rect 31220 1902 31248 3878
rect 31390 3768 31446 3777
rect 31390 3703 31392 3712
rect 31444 3703 31446 3712
rect 31392 3674 31444 3680
rect 31496 3058 31524 4422
rect 31576 4072 31628 4078
rect 31628 4020 31708 4026
rect 31576 4014 31708 4020
rect 31588 3998 31708 4014
rect 31576 3664 31628 3670
rect 31574 3632 31576 3641
rect 31628 3632 31630 3641
rect 31574 3567 31630 3576
rect 31574 3224 31630 3233
rect 31680 3194 31708 3998
rect 31772 3777 31800 4558
rect 32036 4480 32088 4486
rect 32036 4422 32088 4428
rect 32048 4010 32076 4422
rect 32036 4004 32088 4010
rect 32036 3946 32088 3952
rect 31758 3768 31814 3777
rect 31758 3703 31814 3712
rect 32048 3602 32076 3946
rect 32036 3596 32088 3602
rect 32036 3538 32088 3544
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 31772 3233 31800 3470
rect 32036 3392 32088 3398
rect 32036 3334 32088 3340
rect 31758 3224 31814 3233
rect 31574 3159 31576 3168
rect 31628 3159 31630 3168
rect 31668 3188 31720 3194
rect 31576 3130 31628 3136
rect 32048 3194 32076 3334
rect 31758 3159 31814 3168
rect 32036 3188 32088 3194
rect 31668 3130 31720 3136
rect 31772 3058 31800 3159
rect 32036 3130 32088 3136
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 32140 2446 32168 7754
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32324 7410 32352 7686
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32416 6662 32444 8078
rect 32784 7834 32812 9454
rect 32864 9376 32916 9382
rect 32864 9318 32916 9324
rect 32876 9178 32904 9318
rect 32864 9172 32916 9178
rect 32864 9114 32916 9120
rect 32876 7954 32904 9114
rect 33140 9104 33192 9110
rect 33140 9046 33192 9052
rect 32864 7948 32916 7954
rect 32864 7890 32916 7896
rect 32784 7806 32904 7834
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 32600 6458 32628 6802
rect 32784 6798 32812 7346
rect 32876 6866 32904 7806
rect 32956 6996 33008 7002
rect 32956 6938 33008 6944
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32784 6610 32812 6734
rect 32784 6582 32904 6610
rect 32588 6452 32640 6458
rect 32588 6394 32640 6400
rect 32772 6452 32824 6458
rect 32772 6394 32824 6400
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32692 6118 32720 6258
rect 32588 6112 32640 6118
rect 32588 6054 32640 6060
rect 32680 6112 32732 6118
rect 32680 6054 32732 6060
rect 32600 5914 32628 6054
rect 32588 5908 32640 5914
rect 32588 5850 32640 5856
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 32324 4146 32352 5714
rect 32692 5642 32720 6054
rect 32680 5636 32732 5642
rect 32680 5578 32732 5584
rect 32402 5264 32458 5273
rect 32402 5199 32404 5208
rect 32456 5199 32458 5208
rect 32404 5170 32456 5176
rect 32588 5092 32640 5098
rect 32588 5034 32640 5040
rect 32600 4690 32628 5034
rect 32588 4684 32640 4690
rect 32588 4626 32640 4632
rect 32692 4622 32720 5578
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 32680 4276 32732 4282
rect 32680 4218 32732 4224
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32692 3738 32720 4218
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 32508 3194 32536 3674
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32310 3088 32366 3097
rect 32310 3023 32312 3032
rect 32364 3023 32366 3032
rect 32312 2994 32364 3000
rect 32784 2582 32812 6394
rect 32876 6322 32904 6582
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 32876 5302 32904 6258
rect 32968 5914 32996 6938
rect 33048 6860 33100 6866
rect 33048 6802 33100 6808
rect 32956 5908 33008 5914
rect 32956 5850 33008 5856
rect 33060 5370 33088 6802
rect 33152 5778 33180 9046
rect 33428 8022 33456 13874
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34152 8288 34204 8294
rect 34152 8230 34204 8236
rect 33416 8016 33468 8022
rect 33416 7958 33468 7964
rect 34164 7750 34192 8230
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 34164 7410 34192 7686
rect 34152 7404 34204 7410
rect 34152 7346 34204 7352
rect 33232 6792 33284 6798
rect 33232 6734 33284 6740
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33244 6662 33272 6734
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33600 6656 33652 6662
rect 33600 6598 33652 6604
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33140 5568 33192 5574
rect 33140 5510 33192 5516
rect 33048 5364 33100 5370
rect 33048 5306 33100 5312
rect 32864 5296 32916 5302
rect 32864 5238 32916 5244
rect 32876 4282 32904 5238
rect 33046 5128 33102 5137
rect 33046 5063 33048 5072
rect 33100 5063 33102 5072
rect 33048 5034 33100 5040
rect 33048 4820 33100 4826
rect 33048 4762 33100 4768
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 32876 4146 32904 4218
rect 33060 4146 33088 4762
rect 32864 4140 32916 4146
rect 32864 4082 32916 4088
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 32772 2576 32824 2582
rect 32772 2518 32824 2524
rect 31392 2440 31444 2446
rect 31312 2400 31392 2428
rect 31208 1896 31260 1902
rect 31208 1838 31260 1844
rect 30944 870 31064 898
rect 30944 800 30972 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 15474 200 15530 800
rect 17406 200 17462 800
rect 18694 200 18750 800
rect 20626 200 20682 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 27710 200 27766 800
rect 29642 200 29698 800
rect 30930 200 30986 800
rect 31036 762 31064 870
rect 31312 762 31340 2400
rect 31392 2382 31444 2388
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 31484 2372 31536 2378
rect 31484 2314 31536 2320
rect 31496 2106 31524 2314
rect 31484 2100 31536 2106
rect 31484 2042 31536 2048
rect 32876 800 32904 2382
rect 33152 2038 33180 5510
rect 33244 5234 33272 6598
rect 33520 6390 33548 6598
rect 33612 6458 33640 6598
rect 33600 6452 33652 6458
rect 33600 6394 33652 6400
rect 33508 6384 33560 6390
rect 33508 6326 33560 6332
rect 33704 6322 33732 6734
rect 33692 6316 33744 6322
rect 33692 6258 33744 6264
rect 33784 5704 33836 5710
rect 33784 5646 33836 5652
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 33796 5370 33824 5646
rect 33784 5364 33836 5370
rect 33784 5306 33836 5312
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 33508 5228 33560 5234
rect 33508 5170 33560 5176
rect 33520 5098 33548 5170
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 33520 4622 33548 5034
rect 33796 4622 33824 5306
rect 34072 5234 34100 5646
rect 34060 5228 34112 5234
rect 34060 5170 34112 5176
rect 34072 5098 34100 5170
rect 34060 5092 34112 5098
rect 34060 5034 34112 5040
rect 33508 4616 33560 4622
rect 33230 4584 33286 4593
rect 33508 4558 33560 4564
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33230 4519 33232 4528
rect 33284 4519 33286 4528
rect 33232 4490 33284 4496
rect 33324 4480 33376 4486
rect 33324 4422 33376 4428
rect 33336 4146 33364 4422
rect 33324 4140 33376 4146
rect 33324 4082 33376 4088
rect 33336 3534 33364 4082
rect 33520 3602 33548 4558
rect 33796 4146 33824 4558
rect 33876 4480 33928 4486
rect 33876 4422 33928 4428
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 33796 3942 33824 4082
rect 33692 3936 33744 3942
rect 33692 3878 33744 3884
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33508 3596 33560 3602
rect 33508 3538 33560 3544
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 33244 3058 33272 3470
rect 33704 3126 33732 3878
rect 33692 3120 33744 3126
rect 33692 3062 33744 3068
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 33140 2032 33192 2038
rect 33140 1974 33192 1980
rect 33888 1970 33916 4422
rect 34256 2446 34284 8774
rect 34532 8362 34560 8910
rect 34520 8356 34572 8362
rect 34520 8298 34572 8304
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34532 6866 34560 7890
rect 34520 6860 34572 6866
rect 34520 6802 34572 6808
rect 34520 6724 34572 6730
rect 34520 6666 34572 6672
rect 34532 6458 34560 6666
rect 34520 6452 34572 6458
rect 34520 6394 34572 6400
rect 34520 6248 34572 6254
rect 34520 6190 34572 6196
rect 34532 5556 34560 6190
rect 34440 5528 34560 5556
rect 34440 5370 34468 5528
rect 34428 5364 34480 5370
rect 34428 5306 34480 5312
rect 34624 2650 34652 14214
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35452 11694 35480 34886
rect 35532 33516 35584 33522
rect 35532 33458 35584 33464
rect 35544 33318 35572 33458
rect 35532 33312 35584 33318
rect 35532 33254 35584 33260
rect 35544 17066 35572 33254
rect 35624 30252 35676 30258
rect 35624 30194 35676 30200
rect 35636 30054 35664 30194
rect 35624 30048 35676 30054
rect 35624 29990 35676 29996
rect 35636 17134 35664 29990
rect 35728 21350 35756 35866
rect 35808 26512 35860 26518
rect 35808 26454 35860 26460
rect 35820 25945 35848 26454
rect 35806 25936 35862 25945
rect 35806 25871 35862 25880
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 36004 21146 36032 36722
rect 36740 36378 36768 39200
rect 36728 36372 36780 36378
rect 36728 36314 36780 36320
rect 36084 35692 36136 35698
rect 36084 35634 36136 35640
rect 36096 35290 36124 35634
rect 36268 35488 36320 35494
rect 36266 35456 36268 35465
rect 36320 35456 36322 35465
rect 36266 35391 36322 35400
rect 36084 35284 36136 35290
rect 36084 35226 36136 35232
rect 36266 33416 36322 33425
rect 36266 33351 36268 33360
rect 36320 33351 36322 33360
rect 36268 33322 36320 33328
rect 36452 31884 36504 31890
rect 36452 31826 36504 31832
rect 36360 31816 36412 31822
rect 36360 31758 36412 31764
rect 36372 31414 36400 31758
rect 36360 31408 36412 31414
rect 36358 31376 36360 31385
rect 36412 31376 36414 31385
rect 36358 31311 36414 31320
rect 36268 30048 36320 30054
rect 36266 30016 36268 30025
rect 36320 30016 36322 30025
rect 36266 29951 36322 29960
rect 36268 28076 36320 28082
rect 36268 28018 36320 28024
rect 36280 27985 36308 28018
rect 36266 27976 36322 27985
rect 36266 27911 36322 27920
rect 36176 27872 36228 27878
rect 36176 27814 36228 27820
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35992 21140 36044 21146
rect 35992 21082 36044 21088
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 35728 20262 35756 20878
rect 35716 20256 35768 20262
rect 35716 20198 35768 20204
rect 35624 17128 35676 17134
rect 35624 17070 35676 17076
rect 35532 17060 35584 17066
rect 35532 17002 35584 17008
rect 35728 16574 35756 20198
rect 36096 19514 36124 22578
rect 36084 19508 36136 19514
rect 36084 19450 36136 19456
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 35544 16546 35756 16574
rect 35544 15366 35572 16546
rect 35532 15360 35584 15366
rect 35532 15302 35584 15308
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9376 34848 9382
rect 34796 9318 34848 9324
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34716 7274 34744 7414
rect 34704 7268 34756 7274
rect 34704 7210 34756 7216
rect 34716 6798 34744 7210
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34716 6254 34744 6734
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34704 6112 34756 6118
rect 34704 6054 34756 6060
rect 34716 4214 34744 6054
rect 34704 4208 34756 4214
rect 34704 4150 34756 4156
rect 34704 4072 34756 4078
rect 34704 4014 34756 4020
rect 34716 3738 34744 4014
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34808 3126 34836 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35348 8356 35400 8362
rect 35348 8298 35400 8304
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 7478 35388 8298
rect 35440 8288 35492 8294
rect 35440 8230 35492 8236
rect 35452 7954 35480 8230
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 35544 7834 35572 15302
rect 36096 15162 36124 17138
rect 36084 15156 36136 15162
rect 36084 15098 36136 15104
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 36004 13326 36032 14962
rect 35992 13320 36044 13326
rect 35992 13262 36044 13268
rect 35624 9920 35676 9926
rect 35624 9862 35676 9868
rect 35452 7806 35572 7834
rect 35348 7472 35400 7478
rect 35348 7414 35400 7420
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35452 6914 35480 7806
rect 35532 7404 35584 7410
rect 35532 7346 35584 7352
rect 35544 7002 35572 7346
rect 35532 6996 35584 7002
rect 35532 6938 35584 6944
rect 35360 6886 35480 6914
rect 35072 6792 35124 6798
rect 35072 6734 35124 6740
rect 35084 6390 35112 6734
rect 35072 6384 35124 6390
rect 35072 6326 35124 6332
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35360 3670 35388 6886
rect 35544 6458 35572 6938
rect 35532 6452 35584 6458
rect 35532 6394 35584 6400
rect 35440 6384 35492 6390
rect 35440 6326 35492 6332
rect 35452 5710 35480 6326
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 35452 5370 35480 5646
rect 35440 5364 35492 5370
rect 35440 5306 35492 5312
rect 35452 4826 35480 5306
rect 35440 4820 35492 4826
rect 35440 4762 35492 4768
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 35348 3664 35400 3670
rect 35348 3606 35400 3612
rect 35452 3602 35480 3878
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 34794 2952 34850 2961
rect 34794 2887 34796 2896
rect 34848 2887 34850 2896
rect 34796 2858 34848 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 34244 2440 34296 2446
rect 34244 2382 34296 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 33876 1964 33928 1970
rect 33876 1906 33928 1912
rect 34808 800 34836 2382
rect 35360 2145 35388 3062
rect 35636 2446 35664 9862
rect 35898 8936 35954 8945
rect 35898 8871 35900 8880
rect 35952 8871 35954 8880
rect 35900 8842 35952 8848
rect 35912 4622 35940 8842
rect 36004 6914 36032 13262
rect 36188 12442 36216 27814
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36372 23905 36400 24142
rect 36358 23896 36414 23905
rect 36358 23831 36360 23840
rect 36412 23831 36414 23840
rect 36360 23802 36412 23808
rect 36266 22536 36322 22545
rect 36266 22471 36268 22480
rect 36320 22471 36322 22480
rect 36268 22442 36320 22448
rect 36268 20800 36320 20806
rect 36268 20742 36320 20748
rect 36280 20505 36308 20742
rect 36266 20496 36322 20505
rect 36266 20431 36322 20440
rect 36268 18624 36320 18630
rect 36268 18566 36320 18572
rect 36280 18465 36308 18566
rect 36266 18456 36322 18465
rect 36266 18391 36322 18400
rect 36266 17096 36322 17105
rect 36266 17031 36268 17040
rect 36320 17031 36322 17040
rect 36268 17002 36320 17008
rect 36360 15904 36412 15910
rect 36360 15846 36412 15852
rect 36372 15502 36400 15846
rect 36360 15496 36412 15502
rect 36360 15438 36412 15444
rect 36372 15065 36400 15438
rect 36358 15056 36414 15065
rect 36358 14991 36414 15000
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 36280 13025 36308 13126
rect 36266 13016 36322 13025
rect 36266 12951 36322 12960
rect 36176 12436 36228 12442
rect 36176 12378 36228 12384
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 36096 8634 36124 11086
rect 36268 11076 36320 11082
rect 36268 11018 36320 11024
rect 36280 10985 36308 11018
rect 36266 10976 36322 10985
rect 36266 10911 36322 10920
rect 36360 10056 36412 10062
rect 36360 9998 36412 10004
rect 36372 9654 36400 9998
rect 36360 9648 36412 9654
rect 36358 9616 36360 9625
rect 36412 9616 36414 9625
rect 36358 9551 36414 9560
rect 36176 9376 36228 9382
rect 36176 9318 36228 9324
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 36004 6886 36124 6914
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 36004 3398 36032 3946
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 2650 36032 3334
rect 36096 3058 36124 6886
rect 36188 3534 36216 9318
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36280 6914 36308 8298
rect 36360 7880 36412 7886
rect 36360 7822 36412 7828
rect 36372 7585 36400 7822
rect 36358 7576 36414 7585
rect 36358 7511 36360 7520
rect 36412 7511 36414 7520
rect 36360 7482 36412 7488
rect 36464 7478 36492 31826
rect 36544 10464 36596 10470
rect 36544 10406 36596 10412
rect 36452 7472 36504 7478
rect 36452 7414 36504 7420
rect 36280 6886 36400 6914
rect 36372 5710 36400 6886
rect 36360 5704 36412 5710
rect 36360 5646 36412 5652
rect 36372 5545 36400 5646
rect 36358 5536 36414 5545
rect 36358 5471 36414 5480
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 36280 4185 36308 4422
rect 36266 4176 36322 4185
rect 36266 4111 36322 4120
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 36188 2938 36216 3470
rect 36556 3346 36584 10406
rect 36372 3318 36584 3346
rect 36372 2990 36400 3318
rect 36096 2910 36216 2938
rect 36360 2984 36412 2990
rect 36360 2926 36412 2932
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35346 2136 35402 2145
rect 35346 2071 35402 2080
rect 36096 800 36124 2910
rect 31036 734 31340 762
rect 32862 200 32918 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 36372 105 36400 2926
rect 36358 96 36414 105
rect 36358 31 36414 40
<< via2 >>
rect 2778 38120 2834 38176
rect 1674 36760 1730 36816
rect 1674 34720 1730 34776
rect 1674 32680 1730 32736
rect 1674 31320 1730 31376
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1674 29280 1730 29336
rect 1674 27276 1676 27296
rect 1676 27276 1728 27296
rect 1728 27276 1730 27296
rect 1674 27240 1730 27276
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1582 23860 1638 23896
rect 1582 23840 1584 23860
rect 1584 23840 1636 23860
rect 1636 23840 1638 23860
rect 1582 21800 1638 21856
rect 1582 19796 1584 19816
rect 1584 19796 1636 19816
rect 1636 19796 1638 19816
rect 1582 19760 1638 19796
rect 1582 18420 1638 18456
rect 1582 18400 1584 18420
rect 1584 18400 1636 18420
rect 1636 18400 1638 18420
rect 1674 16396 1676 16416
rect 1676 16396 1728 16416
rect 1728 16396 1730 16416
rect 1674 16360 1730 16396
rect 1674 14320 1730 14376
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 1674 12280 1730 12336
rect 1674 10956 1676 10976
rect 1676 10956 1728 10976
rect 1728 10956 1730 10976
rect 1674 10920 1730 10956
rect 1674 8880 1730 8936
rect 1674 6840 1730 6896
rect 1674 5516 1676 5536
rect 1676 5516 1728 5536
rect 1728 5516 1730 5536
rect 1674 5480 1730 5516
rect 1674 3440 1730 3496
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 17222 3440 17278 3496
rect 14830 2896 14886 2952
rect 16670 2896 16726 2952
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19338 11736 19394 11792
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20074 11736 20130 11792
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19338 10124 19394 10160
rect 19338 10104 19340 10124
rect 19340 10104 19392 10124
rect 19392 10104 19394 10124
rect 19614 10548 19616 10568
rect 19616 10548 19668 10568
rect 19668 10548 19670 10568
rect 19614 10512 19670 10548
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19522 8472 19578 8528
rect 19890 8508 19892 8528
rect 19892 8508 19944 8528
rect 19944 8508 19946 8528
rect 19890 8472 19946 8508
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20718 11736 20774 11792
rect 20442 10512 20498 10568
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 1674 1400 1730 1456
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20994 5208 21050 5264
rect 21454 12164 21510 12200
rect 21454 12144 21456 12164
rect 21456 12144 21508 12164
rect 21508 12144 21510 12164
rect 21270 10920 21326 10976
rect 22190 13524 22246 13560
rect 22190 13504 22192 13524
rect 22192 13504 22244 13524
rect 22244 13504 22246 13524
rect 21914 9560 21970 9616
rect 21822 9016 21878 9072
rect 22098 8356 22154 8392
rect 22098 8336 22100 8356
rect 22100 8336 22152 8356
rect 22152 8336 22154 8356
rect 22006 6316 22062 6352
rect 22006 6296 22008 6316
rect 22008 6296 22060 6316
rect 22060 6296 22062 6316
rect 22742 14068 22798 14104
rect 22742 14048 22744 14068
rect 22744 14048 22796 14068
rect 22796 14048 22798 14068
rect 22742 13504 22798 13560
rect 22650 12688 22706 12744
rect 23202 12688 23258 12744
rect 23018 12280 23074 12336
rect 23478 11736 23534 11792
rect 23754 12824 23810 12880
rect 23018 9968 23074 10024
rect 22374 8336 22430 8392
rect 21822 5072 21878 5128
rect 23294 10548 23296 10568
rect 23296 10548 23348 10568
rect 23348 10548 23350 10568
rect 23294 10512 23350 10548
rect 35530 38800 35586 38856
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 25134 13232 25190 13288
rect 24030 11076 24086 11112
rect 24030 11056 24032 11076
rect 24032 11056 24084 11076
rect 24084 11056 24086 11076
rect 23846 9968 23902 10024
rect 23478 6296 23534 6352
rect 23294 4528 23350 4584
rect 25318 15000 25374 15056
rect 24766 9696 24822 9752
rect 24950 9560 25006 9616
rect 23754 3984 23810 4040
rect 24306 3884 24308 3904
rect 24308 3884 24360 3904
rect 24360 3884 24362 3904
rect 24306 3848 24362 3884
rect 24766 3032 24822 3088
rect 24858 2760 24914 2816
rect 25962 13368 26018 13424
rect 26146 12844 26202 12880
rect 26146 12824 26148 12844
rect 26148 12824 26200 12844
rect 26200 12824 26202 12844
rect 25502 12280 25558 12336
rect 25410 9560 25466 9616
rect 25502 2760 25558 2816
rect 26606 12724 26608 12744
rect 26608 12724 26660 12744
rect 26660 12724 26662 12744
rect 26606 12688 26662 12724
rect 27526 13252 27582 13288
rect 27526 13232 27528 13252
rect 27528 13232 27580 13252
rect 27580 13232 27582 13252
rect 26974 12280 27030 12336
rect 27710 13368 27766 13424
rect 26790 9696 26846 9752
rect 28078 14048 28134 14104
rect 28262 15000 28318 15056
rect 27618 11736 27674 11792
rect 27250 8472 27306 8528
rect 27710 10104 27766 10160
rect 27250 5888 27306 5944
rect 28078 12280 28134 12336
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 36266 36760 36322 36816
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 28630 12180 28632 12200
rect 28632 12180 28684 12200
rect 28684 12180 28686 12200
rect 28630 12144 28686 12180
rect 28538 10920 28594 10976
rect 27066 3848 27122 3904
rect 29090 13504 29146 13560
rect 28538 3440 28594 3496
rect 29090 5908 29146 5944
rect 29090 5888 29092 5908
rect 29092 5888 29144 5908
rect 29144 5888 29146 5908
rect 29090 3576 29146 3632
rect 28998 3032 29054 3088
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 30562 3984 30618 4040
rect 29918 3476 29920 3496
rect 29920 3476 29972 3496
rect 29972 3476 29974 3496
rect 29918 3440 29974 3476
rect 31114 3460 31170 3496
rect 31114 3440 31116 3460
rect 31116 3440 31168 3460
rect 31168 3440 31170 3460
rect 31114 2796 31116 2816
rect 31116 2796 31168 2816
rect 31168 2796 31170 2816
rect 31114 2760 31170 2796
rect 31390 3732 31446 3768
rect 31390 3712 31392 3732
rect 31392 3712 31444 3732
rect 31444 3712 31446 3732
rect 31574 3612 31576 3632
rect 31576 3612 31628 3632
rect 31628 3612 31630 3632
rect 31574 3576 31630 3612
rect 31574 3188 31630 3224
rect 31758 3712 31814 3768
rect 31574 3168 31576 3188
rect 31576 3168 31628 3188
rect 31628 3168 31630 3188
rect 31758 3168 31814 3224
rect 32402 5228 32458 5264
rect 32402 5208 32404 5228
rect 32404 5208 32456 5228
rect 32456 5208 32458 5228
rect 32310 3052 32366 3088
rect 32310 3032 32312 3052
rect 32312 3032 32364 3052
rect 32364 3032 32366 3052
rect 33046 5092 33102 5128
rect 33046 5072 33048 5092
rect 33048 5072 33100 5092
rect 33100 5072 33102 5092
rect 33230 4548 33286 4584
rect 33230 4528 33232 4548
rect 33232 4528 33284 4548
rect 33284 4528 33286 4548
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35806 25880 35862 25936
rect 36266 35436 36268 35456
rect 36268 35436 36320 35456
rect 36320 35436 36322 35456
rect 36266 35400 36322 35436
rect 36266 33380 36322 33416
rect 36266 33360 36268 33380
rect 36268 33360 36320 33380
rect 36320 33360 36322 33380
rect 36358 31356 36360 31376
rect 36360 31356 36412 31376
rect 36412 31356 36414 31376
rect 36358 31320 36414 31356
rect 36266 29996 36268 30016
rect 36268 29996 36320 30016
rect 36320 29996 36322 30016
rect 36266 29960 36322 29996
rect 36266 27920 36322 27976
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34794 2916 34850 2952
rect 34794 2896 34796 2916
rect 34796 2896 34848 2916
rect 34848 2896 34850 2916
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35898 8900 35954 8936
rect 35898 8880 35900 8900
rect 35900 8880 35952 8900
rect 35952 8880 35954 8900
rect 36358 23860 36414 23896
rect 36358 23840 36360 23860
rect 36360 23840 36412 23860
rect 36412 23840 36414 23860
rect 36266 22500 36322 22536
rect 36266 22480 36268 22500
rect 36268 22480 36320 22500
rect 36320 22480 36322 22500
rect 36266 20440 36322 20496
rect 36266 18400 36322 18456
rect 36266 17060 36322 17096
rect 36266 17040 36268 17060
rect 36268 17040 36320 17060
rect 36320 17040 36322 17060
rect 36358 15000 36414 15056
rect 36266 12960 36322 13016
rect 36266 10920 36322 10976
rect 36358 9596 36360 9616
rect 36360 9596 36412 9616
rect 36412 9596 36414 9616
rect 36358 9560 36414 9596
rect 36358 7540 36414 7576
rect 36358 7520 36360 7540
rect 36360 7520 36412 7540
rect 36412 7520 36414 7540
rect 36358 5480 36414 5536
rect 36266 4120 36322 4176
rect 35346 2080 35402 2136
rect 36358 40 36414 96
<< metal3 >>
rect 35525 38858 35591 38861
rect 37200 38858 37800 38888
rect 35525 38856 37800 38858
rect 35525 38800 35530 38856
rect 35586 38800 37800 38856
rect 35525 38798 37800 38800
rect 35525 38795 35591 38798
rect 37200 38768 37800 38798
rect 200 38178 800 38208
rect 2773 38178 2839 38181
rect 200 38176 2839 38178
rect 200 38120 2778 38176
rect 2834 38120 2839 38176
rect 200 38118 2839 38120
rect 200 38088 800 38118
rect 2773 38115 2839 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 1669 36818 1735 36821
rect 200 36816 1735 36818
rect 200 36760 1674 36816
rect 1730 36760 1735 36816
rect 200 36758 1735 36760
rect 200 36728 800 36758
rect 1669 36755 1735 36758
rect 36261 36818 36327 36821
rect 37200 36818 37800 36848
rect 36261 36816 37800 36818
rect 36261 36760 36266 36816
rect 36322 36760 37800 36816
rect 36261 36758 37800 36760
rect 36261 36755 36327 36758
rect 37200 36728 37800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 36261 35458 36327 35461
rect 37200 35458 37800 35488
rect 36261 35456 37800 35458
rect 36261 35400 36266 35456
rect 36322 35400 37800 35456
rect 36261 35398 37800 35400
rect 36261 35395 36327 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 37200 35368 37800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1669 34778 1735 34781
rect 200 34776 1735 34778
rect 200 34720 1674 34776
rect 1730 34720 1735 34776
rect 200 34718 1735 34720
rect 200 34688 800 34718
rect 1669 34715 1735 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 36261 33418 36327 33421
rect 37200 33418 37800 33448
rect 36261 33416 37800 33418
rect 36261 33360 36266 33416
rect 36322 33360 37800 33416
rect 36261 33358 37800 33360
rect 36261 33355 36327 33358
rect 37200 33328 37800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1669 32738 1735 32741
rect 200 32736 1735 32738
rect 200 32680 1674 32736
rect 1730 32680 1735 32736
rect 200 32678 1735 32680
rect 200 32648 800 32678
rect 1669 32675 1735 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1669 31378 1735 31381
rect 200 31376 1735 31378
rect 200 31320 1674 31376
rect 1730 31320 1735 31376
rect 200 31318 1735 31320
rect 200 31288 800 31318
rect 1669 31315 1735 31318
rect 36353 31378 36419 31381
rect 37200 31378 37800 31408
rect 36353 31376 37800 31378
rect 36353 31320 36358 31376
rect 36414 31320 37800 31376
rect 36353 31318 37800 31320
rect 36353 31315 36419 31318
rect 37200 31288 37800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 36261 30018 36327 30021
rect 37200 30018 37800 30048
rect 36261 30016 37800 30018
rect 36261 29960 36266 30016
rect 36322 29960 37800 30016
rect 36261 29958 37800 29960
rect 36261 29955 36327 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 37200 29928 37800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1669 29338 1735 29341
rect 200 29336 1735 29338
rect 200 29280 1674 29336
rect 1730 29280 1735 29336
rect 200 29278 1735 29280
rect 200 29248 800 29278
rect 1669 29275 1735 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 36261 27978 36327 27981
rect 37200 27978 37800 28008
rect 36261 27976 37800 27978
rect 36261 27920 36266 27976
rect 36322 27920 37800 27976
rect 36261 27918 37800 27920
rect 36261 27915 36327 27918
rect 37200 27888 37800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1669 27298 1735 27301
rect 200 27296 1735 27298
rect 200 27240 1674 27296
rect 1730 27240 1735 27296
rect 200 27238 1735 27240
rect 200 27208 800 27238
rect 1669 27235 1735 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 35801 25938 35867 25941
rect 37200 25938 37800 25968
rect 35801 25936 37800 25938
rect 35801 25880 35806 25936
rect 35862 25880 37800 25936
rect 35801 25878 37800 25880
rect 35801 25875 35867 25878
rect 37200 25848 37800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25168 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1577 23898 1643 23901
rect 200 23896 1643 23898
rect 200 23840 1582 23896
rect 1638 23840 1643 23896
rect 200 23838 1643 23840
rect 200 23808 800 23838
rect 1577 23835 1643 23838
rect 36353 23898 36419 23901
rect 37200 23898 37800 23928
rect 36353 23896 37800 23898
rect 36353 23840 36358 23896
rect 36414 23840 37800 23896
rect 36353 23838 37800 23840
rect 36353 23835 36419 23838
rect 37200 23808 37800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 36261 22538 36327 22541
rect 37200 22538 37800 22568
rect 36261 22536 37800 22538
rect 36261 22480 36266 22536
rect 36322 22480 37800 22536
rect 36261 22478 37800 22480
rect 36261 22475 36327 22478
rect 37200 22448 37800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 200 21858 800 21888
rect 1577 21858 1643 21861
rect 200 21856 1643 21858
rect 200 21800 1582 21856
rect 1638 21800 1643 21856
rect 200 21798 1643 21800
rect 200 21768 800 21798
rect 1577 21795 1643 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 36261 20498 36327 20501
rect 37200 20498 37800 20528
rect 36261 20496 37800 20498
rect 36261 20440 36266 20496
rect 36322 20440 37800 20496
rect 36261 20438 37800 20440
rect 36261 20435 36327 20438
rect 37200 20408 37800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1577 19818 1643 19821
rect 200 19816 1643 19818
rect 200 19760 1582 19816
rect 1638 19760 1643 19816
rect 200 19758 1643 19760
rect 200 19728 800 19758
rect 1577 19755 1643 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 1577 18458 1643 18461
rect 200 18456 1643 18458
rect 200 18400 1582 18456
rect 1638 18400 1643 18456
rect 200 18398 1643 18400
rect 200 18368 800 18398
rect 1577 18395 1643 18398
rect 36261 18458 36327 18461
rect 37200 18458 37800 18488
rect 36261 18456 37800 18458
rect 36261 18400 36266 18456
rect 36322 18400 37800 18456
rect 36261 18398 37800 18400
rect 36261 18395 36327 18398
rect 37200 18368 37800 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 36261 17098 36327 17101
rect 37200 17098 37800 17128
rect 36261 17096 37800 17098
rect 36261 17040 36266 17096
rect 36322 17040 37800 17096
rect 36261 17038 37800 17040
rect 36261 17035 36327 17038
rect 37200 17008 37800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 200 16418 800 16448
rect 1669 16418 1735 16421
rect 200 16416 1735 16418
rect 200 16360 1674 16416
rect 1730 16360 1735 16416
rect 200 16358 1735 16360
rect 200 16328 800 16358
rect 1669 16355 1735 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 25313 15058 25379 15061
rect 28257 15058 28323 15061
rect 25313 15056 28323 15058
rect 25313 15000 25318 15056
rect 25374 15000 28262 15056
rect 28318 15000 28323 15056
rect 25313 14998 28323 15000
rect 25313 14995 25379 14998
rect 28257 14995 28323 14998
rect 36353 15058 36419 15061
rect 37200 15058 37800 15088
rect 36353 15056 37800 15058
rect 36353 15000 36358 15056
rect 36414 15000 37800 15056
rect 36353 14998 37800 15000
rect 36353 14995 36419 14998
rect 37200 14968 37800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1669 14378 1735 14381
rect 200 14376 1735 14378
rect 200 14320 1674 14376
rect 1730 14320 1735 14376
rect 200 14318 1735 14320
rect 200 14288 800 14318
rect 1669 14315 1735 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 22737 14106 22803 14109
rect 28073 14106 28139 14109
rect 22737 14104 28139 14106
rect 22737 14048 22742 14104
rect 22798 14048 28078 14104
rect 28134 14048 28139 14104
rect 22737 14046 28139 14048
rect 22737 14043 22803 14046
rect 28073 14043 28139 14046
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 22185 13562 22251 13565
rect 22737 13562 22803 13565
rect 29085 13562 29151 13565
rect 22185 13560 29151 13562
rect 22185 13504 22190 13560
rect 22246 13504 22742 13560
rect 22798 13504 29090 13560
rect 29146 13504 29151 13560
rect 22185 13502 29151 13504
rect 22185 13499 22251 13502
rect 22737 13499 22803 13502
rect 29085 13499 29151 13502
rect 25957 13426 26023 13429
rect 27705 13426 27771 13429
rect 25957 13424 27771 13426
rect 25957 13368 25962 13424
rect 26018 13368 27710 13424
rect 27766 13368 27771 13424
rect 25957 13366 27771 13368
rect 25957 13363 26023 13366
rect 27705 13363 27771 13366
rect 25129 13290 25195 13293
rect 27521 13290 27587 13293
rect 25129 13288 27587 13290
rect 25129 13232 25134 13288
rect 25190 13232 27526 13288
rect 27582 13232 27587 13288
rect 25129 13230 27587 13232
rect 25129 13227 25195 13230
rect 27521 13227 27587 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 36261 13018 36327 13021
rect 37200 13018 37800 13048
rect 36261 13016 37800 13018
rect 36261 12960 36266 13016
rect 36322 12960 37800 13016
rect 36261 12958 37800 12960
rect 36261 12955 36327 12958
rect 37200 12928 37800 12958
rect 23749 12882 23815 12885
rect 26141 12882 26207 12885
rect 23749 12880 26207 12882
rect 23749 12824 23754 12880
rect 23810 12824 26146 12880
rect 26202 12824 26207 12880
rect 23749 12822 26207 12824
rect 23749 12819 23815 12822
rect 26141 12819 26207 12822
rect 22645 12746 22711 12749
rect 23197 12746 23263 12749
rect 26601 12746 26667 12749
rect 22645 12744 26667 12746
rect 22645 12688 22650 12744
rect 22706 12688 23202 12744
rect 23258 12688 26606 12744
rect 26662 12688 26667 12744
rect 22645 12686 26667 12688
rect 22645 12683 22711 12686
rect 23197 12683 23263 12686
rect 26601 12683 26667 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 23013 12338 23079 12341
rect 25497 12338 25563 12341
rect 23013 12336 25563 12338
rect 23013 12280 23018 12336
rect 23074 12280 25502 12336
rect 25558 12280 25563 12336
rect 23013 12278 25563 12280
rect 23013 12275 23079 12278
rect 25497 12275 25563 12278
rect 26969 12338 27035 12341
rect 28073 12338 28139 12341
rect 26969 12336 28139 12338
rect 26969 12280 26974 12336
rect 27030 12280 28078 12336
rect 28134 12280 28139 12336
rect 26969 12278 28139 12280
rect 26969 12275 27035 12278
rect 28073 12275 28139 12278
rect 21449 12202 21515 12205
rect 28625 12202 28691 12205
rect 21449 12200 28691 12202
rect 21449 12144 21454 12200
rect 21510 12144 28630 12200
rect 28686 12144 28691 12200
rect 21449 12142 28691 12144
rect 21449 12139 21515 12142
rect 28625 12139 28691 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 19333 11794 19399 11797
rect 20069 11794 20135 11797
rect 20713 11794 20779 11797
rect 19333 11792 20779 11794
rect 19333 11736 19338 11792
rect 19394 11736 20074 11792
rect 20130 11736 20718 11792
rect 20774 11736 20779 11792
rect 19333 11734 20779 11736
rect 19333 11731 19399 11734
rect 20069 11731 20135 11734
rect 20713 11731 20779 11734
rect 23473 11794 23539 11797
rect 27613 11794 27679 11797
rect 23473 11792 27679 11794
rect 23473 11736 23478 11792
rect 23534 11736 27618 11792
rect 27674 11736 27679 11792
rect 23473 11734 27679 11736
rect 23473 11731 23539 11734
rect 27613 11731 27679 11734
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 24025 11114 24091 11117
rect 24710 11114 24716 11116
rect 24025 11112 24716 11114
rect 24025 11056 24030 11112
rect 24086 11056 24716 11112
rect 24025 11054 24716 11056
rect 24025 11051 24091 11054
rect 24710 11052 24716 11054
rect 24780 11052 24786 11116
rect 200 10978 800 11008
rect 1669 10978 1735 10981
rect 200 10976 1735 10978
rect 200 10920 1674 10976
rect 1730 10920 1735 10976
rect 200 10918 1735 10920
rect 200 10888 800 10918
rect 1669 10915 1735 10918
rect 21265 10978 21331 10981
rect 28533 10978 28599 10981
rect 21265 10976 28599 10978
rect 21265 10920 21270 10976
rect 21326 10920 28538 10976
rect 28594 10920 28599 10976
rect 21265 10918 28599 10920
rect 21265 10915 21331 10918
rect 28533 10915 28599 10918
rect 36261 10978 36327 10981
rect 37200 10978 37800 11008
rect 36261 10976 37800 10978
rect 36261 10920 36266 10976
rect 36322 10920 37800 10976
rect 36261 10918 37800 10920
rect 36261 10915 36327 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 37200 10888 37800 10918
rect 19570 10847 19886 10848
rect 19609 10570 19675 10573
rect 20437 10570 20503 10573
rect 23289 10570 23355 10573
rect 19609 10568 23355 10570
rect 19609 10512 19614 10568
rect 19670 10512 20442 10568
rect 20498 10512 23294 10568
rect 23350 10512 23355 10568
rect 19609 10510 23355 10512
rect 19609 10507 19675 10510
rect 20437 10507 20503 10510
rect 23289 10507 23355 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19333 10162 19399 10165
rect 27705 10162 27771 10165
rect 19333 10160 27771 10162
rect 19333 10104 19338 10160
rect 19394 10104 27710 10160
rect 27766 10104 27771 10160
rect 19333 10102 27771 10104
rect 19333 10099 19399 10102
rect 27705 10099 27771 10102
rect 23013 10026 23079 10029
rect 23841 10026 23907 10029
rect 23013 10024 23907 10026
rect 23013 9968 23018 10024
rect 23074 9968 23846 10024
rect 23902 9968 23907 10024
rect 23013 9966 23907 9968
rect 23013 9963 23079 9966
rect 23841 9963 23907 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 24761 9754 24827 9757
rect 26785 9754 26851 9757
rect 24761 9752 26851 9754
rect 24761 9696 24766 9752
rect 24822 9696 26790 9752
rect 26846 9696 26851 9752
rect 24761 9694 26851 9696
rect 24761 9691 24827 9694
rect 26785 9691 26851 9694
rect 21909 9618 21975 9621
rect 24945 9618 25011 9621
rect 25405 9618 25471 9621
rect 21909 9616 25471 9618
rect 21909 9560 21914 9616
rect 21970 9560 24950 9616
rect 25006 9560 25410 9616
rect 25466 9560 25471 9616
rect 21909 9558 25471 9560
rect 21909 9555 21975 9558
rect 24945 9555 25011 9558
rect 25405 9555 25471 9558
rect 36353 9618 36419 9621
rect 37200 9618 37800 9648
rect 36353 9616 37800 9618
rect 36353 9560 36358 9616
rect 36414 9560 37800 9616
rect 36353 9558 37800 9560
rect 36353 9555 36419 9558
rect 37200 9528 37800 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 21817 9074 21883 9077
rect 21817 9072 22110 9074
rect 21817 9016 21822 9072
rect 21878 9016 22110 9072
rect 21817 9014 22110 9016
rect 21817 9011 21883 9014
rect 200 8938 800 8968
rect 1669 8938 1735 8941
rect 200 8936 1735 8938
rect 200 8880 1674 8936
rect 1730 8880 1735 8936
rect 200 8878 1735 8880
rect 22050 8938 22110 9014
rect 35893 8938 35959 8941
rect 22050 8936 35959 8938
rect 22050 8880 35898 8936
rect 35954 8880 35959 8936
rect 22050 8878 35959 8880
rect 200 8848 800 8878
rect 1669 8875 1735 8878
rect 35893 8875 35959 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 19517 8530 19583 8533
rect 19885 8530 19951 8533
rect 27245 8530 27311 8533
rect 19517 8528 27311 8530
rect 19517 8472 19522 8528
rect 19578 8472 19890 8528
rect 19946 8472 27250 8528
rect 27306 8472 27311 8528
rect 19517 8470 27311 8472
rect 19517 8467 19583 8470
rect 19885 8467 19951 8470
rect 27245 8467 27311 8470
rect 22093 8394 22159 8397
rect 22369 8394 22435 8397
rect 22093 8392 22435 8394
rect 22093 8336 22098 8392
rect 22154 8336 22374 8392
rect 22430 8336 22435 8392
rect 22093 8334 22435 8336
rect 22093 8331 22159 8334
rect 22369 8331 22435 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 36353 7578 36419 7581
rect 37200 7578 37800 7608
rect 36353 7576 37800 7578
rect 36353 7520 36358 7576
rect 36414 7520 37800 7576
rect 36353 7518 37800 7520
rect 36353 7515 36419 7518
rect 37200 7488 37800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1669 6898 1735 6901
rect 200 6896 1735 6898
rect 200 6840 1674 6896
rect 1730 6840 1735 6896
rect 200 6838 1735 6840
rect 200 6808 800 6838
rect 1669 6835 1735 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 22001 6354 22067 6357
rect 23473 6354 23539 6357
rect 22001 6352 23539 6354
rect 22001 6296 22006 6352
rect 22062 6296 23478 6352
rect 23534 6296 23539 6352
rect 22001 6294 23539 6296
rect 22001 6291 22067 6294
rect 23473 6291 23539 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 27245 5946 27311 5949
rect 29085 5946 29151 5949
rect 27245 5944 29151 5946
rect 27245 5888 27250 5944
rect 27306 5888 29090 5944
rect 29146 5888 29151 5944
rect 27245 5886 29151 5888
rect 27245 5883 27311 5886
rect 29085 5883 29151 5886
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 36353 5538 36419 5541
rect 37200 5538 37800 5568
rect 36353 5536 37800 5538
rect 36353 5480 36358 5536
rect 36414 5480 37800 5536
rect 36353 5478 37800 5480
rect 36353 5475 36419 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 37200 5448 37800 5478
rect 19570 5407 19886 5408
rect 20989 5266 21055 5269
rect 32397 5266 32463 5269
rect 20989 5264 32463 5266
rect 20989 5208 20994 5264
rect 21050 5208 32402 5264
rect 32458 5208 32463 5264
rect 20989 5206 32463 5208
rect 20989 5203 21055 5206
rect 32397 5203 32463 5206
rect 21817 5130 21883 5133
rect 33041 5130 33107 5133
rect 21817 5128 33107 5130
rect 21817 5072 21822 5128
rect 21878 5072 33046 5128
rect 33102 5072 33107 5128
rect 21817 5070 33107 5072
rect 21817 5067 21883 5070
rect 33041 5067 33107 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 23289 4586 23355 4589
rect 33225 4586 33291 4589
rect 23289 4584 33291 4586
rect 23289 4528 23294 4584
rect 23350 4528 33230 4584
rect 33286 4528 33291 4584
rect 23289 4526 33291 4528
rect 23289 4523 23355 4526
rect 33225 4523 33291 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 36261 4178 36327 4181
rect 37200 4178 37800 4208
rect 36261 4176 37800 4178
rect 36261 4120 36266 4176
rect 36322 4120 37800 4176
rect 36261 4118 37800 4120
rect 36261 4115 36327 4118
rect 37200 4088 37800 4118
rect 23749 4042 23815 4045
rect 30557 4042 30623 4045
rect 23749 4040 30623 4042
rect 23749 3984 23754 4040
rect 23810 3984 30562 4040
rect 30618 3984 30623 4040
rect 23749 3982 30623 3984
rect 23749 3979 23815 3982
rect 30557 3979 30623 3982
rect 24301 3906 24367 3909
rect 27061 3906 27127 3909
rect 24301 3904 27127 3906
rect 24301 3848 24306 3904
rect 24362 3848 27066 3904
rect 27122 3848 27127 3904
rect 24301 3846 27127 3848
rect 24301 3843 24367 3846
rect 27061 3843 27127 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 31385 3770 31451 3773
rect 31753 3770 31819 3773
rect 31385 3768 31819 3770
rect 31385 3712 31390 3768
rect 31446 3712 31758 3768
rect 31814 3712 31819 3768
rect 31385 3710 31819 3712
rect 31385 3707 31451 3710
rect 31753 3707 31819 3710
rect 29085 3634 29151 3637
rect 31569 3634 31635 3637
rect 29085 3632 31635 3634
rect 29085 3576 29090 3632
rect 29146 3576 31574 3632
rect 31630 3576 31635 3632
rect 29085 3574 31635 3576
rect 29085 3571 29151 3574
rect 31569 3571 31635 3574
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 17217 3498 17283 3501
rect 28533 3498 28599 3501
rect 17217 3496 28599 3498
rect 17217 3440 17222 3496
rect 17278 3440 28538 3496
rect 28594 3440 28599 3496
rect 17217 3438 28599 3440
rect 17217 3435 17283 3438
rect 28533 3435 28599 3438
rect 29913 3498 29979 3501
rect 31109 3498 31175 3501
rect 29913 3496 31175 3498
rect 29913 3440 29918 3496
rect 29974 3440 31114 3496
rect 31170 3440 31175 3496
rect 29913 3438 31175 3440
rect 29913 3435 29979 3438
rect 31109 3435 31175 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 24710 3164 24716 3228
rect 24780 3226 24786 3228
rect 31569 3226 31635 3229
rect 31753 3226 31819 3229
rect 24780 3166 31402 3226
rect 24780 3164 24786 3166
rect 24761 3090 24827 3093
rect 28993 3090 29059 3093
rect 24761 3088 29059 3090
rect 24761 3032 24766 3088
rect 24822 3032 28998 3088
rect 29054 3032 29059 3088
rect 24761 3030 29059 3032
rect 31342 3090 31402 3166
rect 31569 3224 31819 3226
rect 31569 3168 31574 3224
rect 31630 3168 31758 3224
rect 31814 3168 31819 3224
rect 31569 3166 31819 3168
rect 31569 3163 31635 3166
rect 31753 3163 31819 3166
rect 32305 3090 32371 3093
rect 31342 3088 32371 3090
rect 31342 3032 32310 3088
rect 32366 3032 32371 3088
rect 31342 3030 32371 3032
rect 24761 3027 24827 3030
rect 28993 3027 29059 3030
rect 32305 3027 32371 3030
rect 14825 2954 14891 2957
rect 16665 2954 16731 2957
rect 34789 2954 34855 2957
rect 14825 2952 34855 2954
rect 14825 2896 14830 2952
rect 14886 2896 16670 2952
rect 16726 2896 34794 2952
rect 34850 2896 34855 2952
rect 14825 2894 34855 2896
rect 14825 2891 14891 2894
rect 16665 2891 16731 2894
rect 34789 2891 34855 2894
rect 24853 2818 24919 2821
rect 25497 2818 25563 2821
rect 31109 2818 31175 2821
rect 24853 2816 31175 2818
rect 24853 2760 24858 2816
rect 24914 2760 25502 2816
rect 25558 2760 31114 2816
rect 31170 2760 31175 2816
rect 24853 2758 31175 2760
rect 24853 2755 24919 2758
rect 25497 2755 25563 2758
rect 31109 2755 31175 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 35341 2138 35407 2141
rect 37200 2138 37800 2168
rect 35341 2136 37800 2138
rect 35341 2080 35346 2136
rect 35402 2080 37800 2136
rect 35341 2078 37800 2080
rect 35341 2075 35407 2078
rect 37200 2048 37800 2078
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 36353 98 36419 101
rect 37200 98 37800 128
rect 36353 96 37800 98
rect 36353 40 36358 96
rect 36414 40 37800 96
rect 36353 38 37800 40
rect 36353 35 36419 38
rect 37200 8 37800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 24716 11052 24780 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 24716 3164 24780 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 24715 11116 24781 11117
rect 24715 11052 24716 11116
rect 24780 11052 24781 11116
rect 24715 11051 24781 11052
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 24718 3229 24778 11051
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 24715 3228 24781 3229
rect 24715 3164 24716 3228
rect 24780 3164 24781 3228
rect 24715 3163 24781 3164
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17112 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1667941163
transform -1 0 29900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1667941163
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1667941163
transform -1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1667941163
transform -1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1667941163
transform -1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1667941163
transform -1 0 26680 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1667941163
transform -1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1667941163
transform -1 0 30452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1667941163
transform 1 0 19504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1667941163
transform -1 0 20976 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1667941163
transform -1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1667941163
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1667941163
transform -1 0 24104 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1667941163
transform -1 0 25208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1667941163
transform -1 0 17664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1667941163
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1667941163
transform -1 0 6716 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1667941163
transform -1 0 25300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1667941163
transform -1 0 29900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1667941163
transform 1 0 21344 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1667941163
transform -1 0 23736 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1667941163
transform -1 0 28060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1667941163
transform 1 0 25944 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1667941163
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A
timestamp 1667941163
transform -1 0 9936 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform 1 0 32108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1667941163
transform -1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1667941163
transform -1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 22816 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform -1 0 35604 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1667941163
transform 1 0 23460 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1667941163
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1667941163
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1667941163
transform 1 0 29716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1667941163
transform -1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A
timestamp 1667941163
transform -1 0 16836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1667941163
transform -1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform -1 0 15916 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1667941163
transform -1 0 33764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1667941163
transform -1 0 34316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1667941163
transform 1 0 30728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 34224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1667941163
transform 1 0 34868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1667941163
transform 1 0 33672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1667941163
transform 1 0 34868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1667941163
transform -1 0 35604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1667941163
transform 1 0 32200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1667941163
transform -1 0 34960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1667941163
transform 1 0 34868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A
timestamp 1667941163
transform 1 0 33580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1667941163
transform 1 0 35696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1667941163
transform 1 0 35328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1667941163
transform 1 0 32752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1667941163
transform 1 0 34776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A
timestamp 1667941163
transform 1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform -1 0 33212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1667941163
transform -1 0 36248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform 1 0 35512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1667941163
transform -1 0 36064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1667941163
transform 1 0 30544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform 1 0 34132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform -1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1667941163
transform 1 0 31648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1667941163
transform -1 0 36432 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform 1 0 31372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1667941163
transform 1 0 34868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1667941163
transform 1 0 30544 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1667941163
transform 1 0 31096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform -1 0 36064 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A
timestamp 1667941163
transform 1 0 32476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform 1 0 35328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1667941163
transform -1 0 34408 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A
timestamp 1667941163
transform -1 0 33856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1667941163
transform 1 0 31648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform 1 0 31648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1667941163
transform 1 0 15180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 1667941163
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__CLK
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__D
timestamp 1667941163
transform 1 0 25392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__CLK
timestamp 1667941163
transform 1 0 35420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__CLK
timestamp 1667941163
transform 1 0 25760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__CLK
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__D
timestamp 1667941163
transform 1 0 29624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__CLK
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__CLK
timestamp 1667941163
transform 1 0 26772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__CLK
timestamp 1667941163
transform 1 0 34224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__D
timestamp 1667941163
transform -1 0 35052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__CLK
timestamp 1667941163
transform 1 0 25944 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__CLK
timestamp 1667941163
transform 1 0 28520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__CLK
timestamp 1667941163
transform 1 0 26220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__CLK
timestamp 1667941163
transform 1 0 28980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__CLK
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__CLK
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__D
timestamp 1667941163
transform -1 0 23276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__CLK
timestamp 1667941163
transform 1 0 23828 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__D
timestamp 1667941163
transform -1 0 23460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__CLK
timestamp 1667941163
transform 1 0 27968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__D
timestamp 1667941163
transform -1 0 26864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__CLK
timestamp 1667941163
transform 1 0 25668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__CLK
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__CLK
timestamp 1667941163
transform -1 0 36340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__CLK
timestamp 1667941163
transform 1 0 26404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__D
timestamp 1667941163
transform 1 0 28980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__CLK
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__CLK
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__CLK
timestamp 1667941163
transform 1 0 26496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__CLK
timestamp 1667941163
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__CLK
timestamp 1667941163
transform 1 0 29992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__CLK
timestamp 1667941163
transform 1 0 29532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__CLK
timestamp 1667941163
transform 1 0 29716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__CLK
timestamp 1667941163
transform 1 0 28612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__CLK
timestamp 1667941163
transform 1 0 29072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__CLK
timestamp 1667941163
transform 1 0 26496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__CLK
timestamp 1667941163
transform 1 0 28980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__CLK
timestamp 1667941163
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__CLK
timestamp 1667941163
transform 1 0 25208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__CLK
timestamp 1667941163
transform 1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__CLK
timestamp 1667941163
transform 1 0 30360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__CLK
timestamp 1667941163
transform 1 0 23552 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__CLK
timestamp 1667941163
transform 1 0 25944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__CLK
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__CLK
timestamp 1667941163
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__CLK
timestamp 1667941163
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1667941163
transform 1 0 12696 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform -1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform -1 0 7360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform 1 0 17112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1667941163
transform -1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform -1 0 30544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform -1 0 27416 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform -1 0 23460 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform -1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1667941163
transform 1 0 35696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform -1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1667941163
transform -1 0 28244 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1667941163
transform -1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1667941163
transform -1 0 5520 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1667941163
transform -1 0 4784 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1667941163
transform -1 0 24012 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform -1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform -1 0 35512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform 1 0 12328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1667941163
transform -1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1667941163
transform -1 0 30544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1667941163
transform -1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1667941163
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 36432 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 36432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 35696 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 1748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 36432 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 4876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 18400 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform 1 0 21344 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 35328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 35052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 36432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 35052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 24564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform 1 0 16192 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 1748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 31280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 35696 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 24288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 2392 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 36432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 11868 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 36432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 25024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 6808 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 1748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 13156 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 23644 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output46_A
timestamp 1667941163
transform 1 0 35512 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1667941163
transform 1 0 28796 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1667941163
transform 1 0 35512 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1667941163
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1667941163
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1667941163
transform -1 0 34132 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1667941163
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1667941163
transform 1 0 18216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1667941163
transform 1 0 35880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1667941163
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1667941163
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 1667941163
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1667941163
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1667941163
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1667941163
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1667941163
transform 1 0 20608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1667941163
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_383
timestamp 1667941163
transform 1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_21
timestamp 1667941163
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1667941163
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1667941163
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_118
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1667941163
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_133
timestamp 1667941163
transform 1 0 13340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1667941163
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_150
timestamp 1667941163
transform 1 0 14904 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp 1667941163
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_173
timestamp 1667941163
transform 1 0 17020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_185
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_201
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1667941163
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1667941163
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_238
timestamp 1667941163
transform 1 0 23000 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_246
timestamp 1667941163
transform 1 0 23736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1667941163
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1667941163
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_327
timestamp 1667941163
transform 1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1667941163
transform 1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_350
timestamp 1667941163
transform 1 0 33304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_357
timestamp 1667941163
transform 1 0 33948 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1667941163
transform 1 0 34684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1667941163
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1667941163
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_103
timestamp 1667941163
transform 1 0 10580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_115
timestamp 1667941163
transform 1 0 11684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_127
timestamp 1667941163
transform 1 0 12788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1667941163
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_155
timestamp 1667941163
transform 1 0 15364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_167
timestamp 1667941163
transform 1 0 16468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1667941163
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1667941163
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_186
timestamp 1667941163
transform 1 0 18216 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1667941163
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1667941163
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1667941163
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1667941163
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_299
timestamp 1667941163
transform 1 0 28612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1667941163
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1667941163
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 1667941163
transform 1 0 32200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_352
timestamp 1667941163
transform 1 0 33488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1667941163
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1667941163
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_375
timestamp 1667941163
transform 1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_379
timestamp 1667941163
transform 1 0 35972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_384
timestamp 1667941163
transform 1 0 36432 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1667941163
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1667941163
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1667941163
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1667941163
transform 1 0 18032 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_192
timestamp 1667941163
transform 1 0 18768 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_196
timestamp 1667941163
transform 1 0 19136 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_208
timestamp 1667941163
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_248
timestamp 1667941163
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1667941163
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp 1667941163
transform 1 0 27324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_306
timestamp 1667941163
transform 1 0 29256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1667941163
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1667941163
transform 1 0 32568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_356
timestamp 1667941163
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_362
timestamp 1667941163
transform 1 0 34408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1667941163
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_374
timestamp 1667941163
transform 1 0 35512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_380
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_131
timestamp 1667941163
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_145
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_155
timestamp 1667941163
transform 1 0 15364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1667941163
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1667941163
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_179
timestamp 1667941163
transform 1 0 17572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1667941163
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1667941163
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1667941163
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1667941163
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1667941163
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_263
timestamp 1667941163
transform 1 0 25300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_269
timestamp 1667941163
transform 1 0 25852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_281
timestamp 1667941163
transform 1 0 26956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1667941163
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1667941163
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_337
timestamp 1667941163
transform 1 0 32108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_344
timestamp 1667941163
transform 1 0 32752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_351
timestamp 1667941163
transform 1 0 33396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_358
timestamp 1667941163
transform 1 0 34040 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_369
timestamp 1667941163
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_375
timestamp 1667941163
transform 1 0 35604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_379
timestamp 1667941163
transform 1 0 35972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_384
timestamp 1667941163
transform 1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1667941163
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1667941163
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_188
timestamp 1667941163
transform 1 0 18400 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1667941163
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_204
timestamp 1667941163
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_229
timestamp 1667941163
transform 1 0 22172 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_239
timestamp 1667941163
transform 1 0 23092 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1667941163
transform 1 0 23460 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_246
timestamp 1667941163
transform 1 0 23736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_252
timestamp 1667941163
transform 1 0 24288 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_260
timestamp 1667941163
transform 1 0 25024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_266
timestamp 1667941163
transform 1 0 25576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_272
timestamp 1667941163
transform 1 0 26128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_303
timestamp 1667941163
transform 1 0 28980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_311
timestamp 1667941163
transform 1 0 29716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_320
timestamp 1667941163
transform 1 0 30544 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_327
timestamp 1667941163
transform 1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1667941163
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_342
timestamp 1667941163
transform 1 0 32568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_356
timestamp 1667941163
transform 1 0 33856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_362
timestamp 1667941163
transform 1 0 34408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_368
timestamp 1667941163
transform 1 0 34960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_374
timestamp 1667941163
transform 1 0 35512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_380
timestamp 1667941163
transform 1 0 36064 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_171
timestamp 1667941163
transform 1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1667941163
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_185
timestamp 1667941163
transform 1 0 18124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1667941163
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1667941163
transform 1 0 20240 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_237
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_243
timestamp 1667941163
transform 1 0 23460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1667941163
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_257
timestamp 1667941163
transform 1 0 24748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_263
timestamp 1667941163
transform 1 0 25300 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_266
timestamp 1667941163
transform 1 0 25576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_272
timestamp 1667941163
transform 1 0 26128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_280
timestamp 1667941163
transform 1 0 26864 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_284
timestamp 1667941163
transform 1 0 27232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1667941163
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_338
timestamp 1667941163
transform 1 0 32200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_352
timestamp 1667941163
transform 1 0 33488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1667941163
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1667941163
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_384
timestamp 1667941163
transform 1 0 36432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_10
timestamp 1667941163
transform 1 0 2024 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_22
timestamp 1667941163
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_34
timestamp 1667941163
transform 1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1667941163
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1667941163
transform 1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1667941163
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_198
timestamp 1667941163
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_248
timestamp 1667941163
transform 1 0 23920 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_254
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_285
timestamp 1667941163
transform 1 0 27324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_310
timestamp 1667941163
transform 1 0 29624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_316
timestamp 1667941163
transform 1 0 30176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_322
timestamp 1667941163
transform 1 0 30728 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_330
timestamp 1667941163
transform 1 0 31464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1667941163
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_344
timestamp 1667941163
transform 1 0 32752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_351
timestamp 1667941163
transform 1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_358
timestamp 1667941163
transform 1 0 34040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_365
timestamp 1667941163
transform 1 0 34684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_372
timestamp 1667941163
transform 1 0 35328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_378
timestamp 1667941163
transform 1 0 35880 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_384
timestamp 1667941163
transform 1 0 36432 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_90
timestamp 1667941163
transform 1 0 9384 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_102
timestamp 1667941163
transform 1 0 10488 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_114
timestamp 1667941163
transform 1 0 11592 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_126
timestamp 1667941163
transform 1 0 12696 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_173
timestamp 1667941163
transform 1 0 17020 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_179
timestamp 1667941163
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1667941163
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1667941163
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_208
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_237
timestamp 1667941163
transform 1 0 22908 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1667941163
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_257
timestamp 1667941163
transform 1 0 24748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_263
timestamp 1667941163
transform 1 0 25300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1667941163
transform 1 0 27600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1667941163
transform 1 0 28152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_300
timestamp 1667941163
transform 1 0 28704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1667941163
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_313
timestamp 1667941163
transform 1 0 29900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_324
timestamp 1667941163
transform 1 0 30912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_328
timestamp 1667941163
transform 1 0 31280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_331
timestamp 1667941163
transform 1 0 31556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_340
timestamp 1667941163
transform 1 0 32384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_347
timestamp 1667941163
transform 1 0 33028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_354
timestamp 1667941163
transform 1 0 33672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1667941163
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_370
timestamp 1667941163
transform 1 0 35144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_376
timestamp 1667941163
transform 1 0 35696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_382
timestamp 1667941163
transform 1 0 36248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 1667941163
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1667941163
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1667941163
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1667941163
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_248
timestamp 1667941163
transform 1 0 23920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_270
timestamp 1667941163
transform 1 0 25944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_274
timestamp 1667941163
transform 1 0 26312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_306
timestamp 1667941163
transform 1 0 29256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_312
timestamp 1667941163
transform 1 0 29808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_322
timestamp 1667941163
transform 1 0 30728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_328
timestamp 1667941163
transform 1 0 31280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1667941163
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_343
timestamp 1667941163
transform 1 0 32660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_350
timestamp 1667941163
transform 1 0 33304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_357
timestamp 1667941163
transform 1 0 33948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_363
timestamp 1667941163
transform 1 0 34500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_369
timestamp 1667941163
transform 1 0 35052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_375
timestamp 1667941163
transform 1 0 35604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_381
timestamp 1667941163
transform 1 0 36156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_384
timestamp 1667941163
transform 1 0 36432 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1667941163
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1667941163
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_207
timestamp 1667941163
transform 1 0 20148 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1667941163
transform 1 0 22816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1667941163
transform 1 0 25392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1667941163
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1667941163
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_313
timestamp 1667941163
transform 1 0 29900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_325
timestamp 1667941163
transform 1 0 31004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_328
timestamp 1667941163
transform 1 0 31280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1667941163
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_340
timestamp 1667941163
transform 1 0 32384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_349
timestamp 1667941163
transform 1 0 33212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_355
timestamp 1667941163
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1667941163
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_369
timestamp 1667941163
transform 1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_373
timestamp 1667941163
transform 1 0 35420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_384
timestamp 1667941163
transform 1 0 36432 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp 1667941163
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_290
timestamp 1667941163
transform 1 0 27784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_314
timestamp 1667941163
transform 1 0 29992 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_320
timestamp 1667941163
transform 1 0 30544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1667941163
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_343
timestamp 1667941163
transform 1 0 32660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_350
timestamp 1667941163
transform 1 0 33304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_356
timestamp 1667941163
transform 1 0 33856 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_362
timestamp 1667941163
transform 1 0 34408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_366
timestamp 1667941163
transform 1 0 34776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_369
timestamp 1667941163
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_375
timestamp 1667941163
transform 1 0 35604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_381
timestamp 1667941163
transform 1 0 36156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 1667941163
transform 1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1667941163
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1667941163
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1667941163
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_275
timestamp 1667941163
transform 1 0 26404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_299
timestamp 1667941163
transform 1 0 28612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1667941163
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_337
timestamp 1667941163
transform 1 0 32108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_340
timestamp 1667941163
transform 1 0 32384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_346
timestamp 1667941163
transform 1 0 32936 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_352
timestamp 1667941163
transform 1 0 33488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_355
timestamp 1667941163
transform 1 0 33764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1667941163
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_369
timestamp 1667941163
transform 1 0 35052 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_380
timestamp 1667941163
transform 1 0 36064 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1667941163
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1667941163
transform 1 0 18400 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1667941163
transform 1 0 19504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1667941163
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_247
timestamp 1667941163
transform 1 0 23828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_271
timestamp 1667941163
transform 1 0 26036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1667941163
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_299
timestamp 1667941163
transform 1 0 28612 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_345
timestamp 1667941163
transform 1 0 32844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_353
timestamp 1667941163
transform 1 0 33580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_356
timestamp 1667941163
transform 1 0 33856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_362
timestamp 1667941163
transform 1 0 34408 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_372
timestamp 1667941163
transform 1 0 35328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_378
timestamp 1667941163
transform 1 0 35880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_384
timestamp 1667941163
transform 1 0 36432 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_72
timestamp 1667941163
transform 1 0 7728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1667941163
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1667941163
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1667941163
transform 1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_214
timestamp 1667941163
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_231
timestamp 1667941163
transform 1 0 22356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_244
timestamp 1667941163
transform 1 0 23552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_259
timestamp 1667941163
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 1667941163
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1667941163
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1667941163
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_298
timestamp 1667941163
transform 1 0 28520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1667941163
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_369
timestamp 1667941163
transform 1 0 35052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_373
timestamp 1667941163
transform 1 0 35420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_384
timestamp 1667941163
transform 1 0 36432 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_175
timestamp 1667941163
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1667941163
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1667941163
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1667941163
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1667941163
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1667941163
transform 1 0 23184 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_257
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_263
timestamp 1667941163
transform 1 0 25300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1667941163
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_296
timestamp 1667941163
transform 1 0 28336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1667941163
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_310
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_381
timestamp 1667941163
transform 1 0 36156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_384
timestamp 1667941163
transform 1 0 36432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1667941163
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_169
timestamp 1667941163
transform 1 0 16652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1667941163
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_212
timestamp 1667941163
transform 1 0 20608 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1667941163
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1667941163
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_273
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_294
timestamp 1667941163
transform 1 0 28152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_373
timestamp 1667941163
transform 1 0 35420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_376
timestamp 1667941163
transform 1 0 35696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_384
timestamp 1667941163
transform 1 0 36432 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_79
timestamp 1667941163
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_91
timestamp 1667941163
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1667941163
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_150
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1667941163
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 1667941163
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1667941163
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1667941163
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1667941163
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_236
timestamp 1667941163
transform 1 0 22816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_243
timestamp 1667941163
transform 1 0 23460 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1667941163
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1667941163
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1667941163
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1667941163
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_314
timestamp 1667941163
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_326
timestamp 1667941163
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1667941163
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_73
timestamp 1667941163
transform 1 0 7820 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1667941163
transform 1 0 12880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1667941163
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_182
timestamp 1667941163
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_207
timestamp 1667941163
transform 1 0 20148 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_214
timestamp 1667941163
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1667941163
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1667941163
transform 1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_286
timestamp 1667941163
transform 1 0 27416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_293
timestamp 1667941163
transform 1 0 28060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_300
timestamp 1667941163
transform 1 0 28704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1667941163
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_313
timestamp 1667941163
transform 1 0 29900 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_319
timestamp 1667941163
transform 1 0 30452 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_331
timestamp 1667941163
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_343
timestamp 1667941163
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1667941163
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_385
timestamp 1667941163
transform 1 0 36524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1667941163
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_22
timestamp 1667941163
transform 1 0 3128 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_34
timestamp 1667941163
transform 1 0 4232 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1667941163
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1667941163
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1667941163
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_202
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_213
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1667941163
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_244
timestamp 1667941163
transform 1 0 23552 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1667941163
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_267
timestamp 1667941163
transform 1 0 25668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1667941163
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1667941163
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_307
timestamp 1667941163
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_313
timestamp 1667941163
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1667941163
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1667941163
transform 1 0 16836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_174
timestamp 1667941163
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1667941163
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_225
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_232
timestamp 1667941163
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_236
timestamp 1667941163
transform 1 0 22816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_258
timestamp 1667941163
transform 1 0 24840 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1667941163
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1667941163
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_299
timestamp 1667941163
transform 1 0 28612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_314
timestamp 1667941163
transform 1 0 29992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_320
timestamp 1667941163
transform 1 0 30544 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_328
timestamp 1667941163
transform 1 0 31280 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_334
timestamp 1667941163
transform 1 0 31832 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_346
timestamp 1667941163
transform 1 0 32936 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_358
timestamp 1667941163
transform 1 0 34040 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_384
timestamp 1667941163
transform 1 0 36432 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1667941163
transform 1 0 17204 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1667941163
transform 1 0 19504 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1667941163
transform 1 0 19872 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_214
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1667941163
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_236
timestamp 1667941163
transform 1 0 22816 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1667941163
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_260
timestamp 1667941163
transform 1 0 25024 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_270
timestamp 1667941163
transform 1 0 25944 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_296
timestamp 1667941163
transform 1 0 28336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_304
timestamp 1667941163
transform 1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_311
timestamp 1667941163
transform 1 0 29716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_318
timestamp 1667941163
transform 1 0 30360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1667941163
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1667941163
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1667941163
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1667941163
transform 1 0 20148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_211
timestamp 1667941163
transform 1 0 20516 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1667941163
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_238
timestamp 1667941163
transform 1 0 23000 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_264
timestamp 1667941163
transform 1 0 25392 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_273
timestamp 1667941163
transform 1 0 26220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1667941163
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1667941163
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_320
timestamp 1667941163
transform 1 0 30544 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_332
timestamp 1667941163
transform 1 0 31648 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_344
timestamp 1667941163
transform 1 0 32752 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_356
timestamp 1667941163
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_385
timestamp 1667941163
transform 1 0 36524 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_176
timestamp 1667941163
transform 1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1667941163
transform 1 0 17940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1667941163
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1667941163
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1667941163
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1667941163
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_255
timestamp 1667941163
transform 1 0 24564 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1667941163
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1667941163
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_300
timestamp 1667941163
transform 1 0 28704 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_307
timestamp 1667941163
transform 1 0 29348 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_313
timestamp 1667941163
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_325
timestamp 1667941163
transform 1 0 31004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1667941163
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_377
timestamp 1667941163
transform 1 0 35788 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_381
timestamp 1667941163
transform 1 0 36156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_185
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_188
timestamp 1667941163
transform 1 0 18400 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1667941163
transform 1 0 19596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1667941163
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1667941163
transform 1 0 22724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1667941163
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_266
timestamp 1667941163
transform 1 0 25576 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1667941163
transform 1 0 26312 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1667941163
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_291
timestamp 1667941163
transform 1 0 27876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_298
timestamp 1667941163
transform 1 0 28520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1667941163
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_329
timestamp 1667941163
transform 1 0 31372 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_339
timestamp 1667941163
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1667941163
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_373
timestamp 1667941163
transform 1 0 35420 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_384
timestamp 1667941163
transform 1 0 36432 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1667941163
transform 1 0 11960 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_124
timestamp 1667941163
transform 1 0 12512 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_136
timestamp 1667941163
transform 1 0 13616 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_148
timestamp 1667941163
transform 1 0 14720 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1667941163
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_204
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_216
timestamp 1667941163
transform 1 0 20976 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1667941163
transform 1 0 23184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_247
timestamp 1667941163
transform 1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_262
timestamp 1667941163
transform 1 0 25208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1667941163
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_299
timestamp 1667941163
transform 1 0 28612 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_311
timestamp 1667941163
transform 1 0 29716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_323
timestamp 1667941163
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_381
timestamp 1667941163
transform 1 0 36156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_384
timestamp 1667941163
transform 1 0 36432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1667941163
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1667941163
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1667941163
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_217
timestamp 1667941163
transform 1 0 21068 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_223
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1667941163
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_232
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1667941163
transform 1 0 23276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1667941163
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_258
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_280
timestamp 1667941163
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_287
timestamp 1667941163
transform 1 0 27508 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1667941163
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1667941163
transform 1 0 36524 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1667941163
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1667941163
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1667941163
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_239
timestamp 1667941163
transform 1 0 23092 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1667941163
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_264
timestamp 1667941163
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_271
timestamp 1667941163
transform 1 0 26036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_379
timestamp 1667941163
transform 1 0 35972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_384
timestamp 1667941163
transform 1 0 36432 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1667941163
transform 1 0 20700 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_216
timestamp 1667941163
transform 1 0 20976 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1667941163
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1667941163
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1667941163
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_259
timestamp 1667941163
transform 1 0 24932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_266
timestamp 1667941163
transform 1 0 25576 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_272
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_278
timestamp 1667941163
transform 1 0 26680 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_290
timestamp 1667941163
transform 1 0 27784 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1667941163
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_351
timestamp 1667941163
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1667941163
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_7
timestamp 1667941163
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_19
timestamp 1667941163
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1667941163
transform 1 0 22172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 1667941163
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_243
timestamp 1667941163
transform 1 0 23460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_247
timestamp 1667941163
transform 1 0 23828 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_250
timestamp 1667941163
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_262
timestamp 1667941163
transform 1 0 25208 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1667941163
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_286
timestamp 1667941163
transform 1 0 27416 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_298
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_310
timestamp 1667941163
transform 1 0 29624 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_322
timestamp 1667941163
transform 1 0 30728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1667941163
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_9
timestamp 1667941163
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1667941163
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_241
timestamp 1667941163
transform 1 0 23276 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_327
timestamp 1667941163
transform 1 0 31188 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_339
timestamp 1667941163
transform 1 0 32292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_351
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_384
timestamp 1667941163
transform 1 0 36432 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_7
timestamp 1667941163
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_19
timestamp 1667941163
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1667941163
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1667941163
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_368
timestamp 1667941163
transform 1 0 34960 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_374
timestamp 1667941163
transform 1 0 35512 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_314
timestamp 1667941163
transform 1 0 29992 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_320
timestamp 1667941163
transform 1 0 30544 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_332
timestamp 1667941163
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_344
timestamp 1667941163
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1667941163
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_385
timestamp 1667941163
transform 1 0 36524 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_378
timestamp 1667941163
transform 1 0 35880 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_90
timestamp 1667941163
transform 1 0 9384 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_96
timestamp 1667941163
transform 1 0 9936 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_108
timestamp 1667941163
transform 1 0 11040 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_120
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1667941163
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_376
timestamp 1667941163
transform 1 0 35696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_384
timestamp 1667941163
transform 1 0 36432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1667941163
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_19
timestamp 1667941163
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1667941163
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_189
timestamp 1667941163
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1667941163
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_202
timestamp 1667941163
transform 1 0 19688 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1667941163
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_385
timestamp 1667941163
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_379
timestamp 1667941163
transform 1 0 35972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_384
timestamp 1667941163
transform 1 0 36432 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_37
timestamp 1667941163
transform 1 0 4508 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1667941163
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_48
timestamp 1667941163
transform 1 0 5520 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_60
timestamp 1667941163
transform 1 0 6624 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_72
timestamp 1667941163
transform 1 0 7728 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_385
timestamp 1667941163
transform 1 0 36524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_7
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_19
timestamp 1667941163
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_31
timestamp 1667941163
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_43
timestamp 1667941163
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_68
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_80
timestamp 1667941163
transform 1 0 8464 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_92
timestamp 1667941163
transform 1 0 9568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1667941163
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_122
timestamp 1667941163
transform 1 0 12328 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_128
timestamp 1667941163
transform 1 0 12880 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_140
timestamp 1667941163
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1667941163
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_381
timestamp 1667941163
transform 1 0 36156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_384
timestamp 1667941163
transform 1 0 36432 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_373
timestamp 1667941163
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_384
timestamp 1667941163
transform 1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1667941163
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1667941163
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_385
timestamp 1667941163
transform 1 0 36524 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1667941163
transform 1 0 26864 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_286
timestamp 1667941163
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_298
timestamp 1667941163
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_384
timestamp 1667941163
transform 1 0 36432 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1667941163
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_385
timestamp 1667941163
transform 1 0 36524 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_376
timestamp 1667941163
transform 1 0 35696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_384
timestamp 1667941163
transform 1 0 36432 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_385
timestamp 1667941163
transform 1 0 36524 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1667941163
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_49
timestamp 1667941163
transform 1 0 5612 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_55
timestamp 1667941163
transform 1 0 6164 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_61
timestamp 1667941163
transform 1 0 6716 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_73
timestamp 1667941163
transform 1 0 7820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 1667941163
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_117
timestamp 1667941163
transform 1 0 11868 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_385
timestamp 1667941163
transform 1 0 36524 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_376
timestamp 1667941163
transform 1 0 35696 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_384
timestamp 1667941163
transform 1 0 36432 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_10
timestamp 1667941163
transform 1 0 2024 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1667941163
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_385
timestamp 1667941163
transform 1 0 36524 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_7
timestamp 1667941163
transform 1 0 1748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_11
timestamp 1667941163
transform 1 0 2116 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_17
timestamp 1667941163
transform 1 0 2668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_29
timestamp 1667941163
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_41
timestamp 1667941163
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1667941163
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_201
timestamp 1667941163
transform 1 0 19596 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_206
timestamp 1667941163
transform 1 0 20056 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_218
timestamp 1667941163
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_240
timestamp 1667941163
transform 1 0 23184 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_246
timestamp 1667941163
transform 1 0 23736 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_258
timestamp 1667941163
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1667941163
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_285
timestamp 1667941163
transform 1 0 27324 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_289
timestamp 1667941163
transform 1 0 27692 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_295
timestamp 1667941163
transform 1 0 28244 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_307
timestamp 1667941163
transform 1 0 29348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_319
timestamp 1667941163
transform 1 0 30452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_331
timestamp 1667941163
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_381
timestamp 1667941163
transform 1 0 36156 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_384
timestamp 1667941163
transform 1 0 36432 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1667941163
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_34
timestamp 1667941163
transform 1 0 4232 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_40
timestamp 1667941163
transform 1 0 4784 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_52
timestamp 1667941163
transform 1 0 5888 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_64
timestamp 1667941163
transform 1 0 6992 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_76
timestamp 1667941163
transform 1 0 8096 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_373
timestamp 1667941163
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_384
timestamp 1667941163
transform 1 0 36432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1667941163
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_19
timestamp 1667941163
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1667941163
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_43
timestamp 1667941163
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1667941163
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_385
timestamp 1667941163
transform 1 0 36524 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_376
timestamp 1667941163
transform 1 0 35696 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_384
timestamp 1667941163
transform 1 0 36432 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_385
timestamp 1667941163
transform 1 0 36524 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1667941163
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1667941163
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_375
timestamp 1667941163
transform 1 0 35604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_383
timestamp 1667941163
transform 1 0 36340 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_379
timestamp 1667941163
transform 1 0 35972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_384
timestamp 1667941163
transform 1 0 36432 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_14
timestamp 1667941163
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_384
timestamp 1667941163
transform 1 0 36432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_31
timestamp 1667941163
transform 1 0 3956 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_177
timestamp 1667941163
transform 1 0 17388 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_182
timestamp 1667941163
transform 1 0 17848 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_190
timestamp 1667941163
transform 1 0 18584 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_194
timestamp 1667941163
transform 1 0 18952 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_206
timestamp 1667941163
transform 1 0 20056 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1667941163
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_236
timestamp 1667941163
transform 1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_243
timestamp 1667941163
transform 1 0 23460 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_255
timestamp 1667941163
transform 1 0 24564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_267
timestamp 1667941163
transform 1 0 25668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_303
timestamp 1667941163
transform 1 0 28980 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_315
timestamp 1667941163
transform 1 0 30084 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_327
timestamp 1667941163
transform 1 0 31188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_359
timestamp 1667941163
transform 1 0 34132 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_371
timestamp 1667941163
transform 1 0 35236 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_379
timestamp 1667941163
transform 1 0 35972 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_384
timestamp 1667941163
transform 1 0 36432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_14
timestamp 1667941163
transform 1 0 2392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 1667941163
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_76
timestamp 1667941163
transform 1 0 8096 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_93
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_99
timestamp 1667941163
transform 1 0 10212 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_117
timestamp 1667941163
transform 1 0 11868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_131
timestamp 1667941163
transform 1 0 13156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_135
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1667941163
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_163
timestamp 1667941163
transform 1 0 16100 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_174
timestamp 1667941163
transform 1 0 17112 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_215
timestamp 1667941163
transform 1 0 20884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_219
timestamp 1667941163
transform 1 0 21252 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_239
timestamp 1667941163
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_271
timestamp 1667941163
transform 1 0 26036 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_295
timestamp 1667941163
transform 1 0 28244 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_327
timestamp 1667941163
transform 1 0 31188 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 36892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 36892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 36892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 36892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 36892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 36892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 36892 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 36892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 36892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 36892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 36892 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 36892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 36892 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 36892 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 36892 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 36892 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 36892 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 36892 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 36892 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 36892 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 36892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 36892 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1667941163
transform 1 0 28428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1667941163
transform 1 0 27140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1667941163
transform 1 0 27784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1667941163
transform -1 0 16928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1667941163
transform -1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1667941163
transform 1 0 28520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1667941163
transform -1 0 24104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1667941163
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1667941163
transform -1 0 18952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1667941163
transform -1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1667941163
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1667941163
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1667941163
transform -1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1667941163
transform -1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1667941163
transform -1 0 17572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1667941163
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1667941163
transform -1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1667941163
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1667941163
transform -1 0 29716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1667941163
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1667941163
transform -1 0 28060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1667941163
transform -1 0 29348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1667941163
transform 1 0 29072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1667941163
transform 1 0 29716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1667941163
transform -1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1667941163
transform -1 0 27416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1667941163
transform -1 0 28980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1667941163
transform -1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1667941163
transform 1 0 22172 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1667941163
transform 1 0 19596 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1667941163
transform 1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1667941163
transform -1 0 28704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1667941163
transform -1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1667941163
transform -1 0 24840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1667941163
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1667941163
transform -1 0 18952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1667941163
transform -1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1667941163
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1667941163
transform 1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1667941163
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1667941163
transform 1 0 27600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1667941163
transform 1 0 26404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1667941163
transform -1 0 28060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1667941163
transform -1 0 28704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1667941163
transform -1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1667941163
transform -1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1667941163
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1667941163
transform 1 0 30360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1667941163
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1667941163
transform 1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1667941163
transform -1 0 27416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1667941163
transform -1 0 28520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1667941163
transform -1 0 25392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1667941163
transform -1 0 23552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1667941163
transform -1 0 23920 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1667941163
transform -1 0 29624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1667941163
transform -1 0 27508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1667941163
transform -1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1667941163
transform -1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1667941163
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1667941163
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1667941163
transform -1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1667941163
transform -1 0 17848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1667941163
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1667941163
transform -1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1667941163
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1667941163
transform 1 0 20516 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1667941163
transform 1 0 26036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform -1 0 6164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform -1 0 31004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform -1 0 24656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform -1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform 1 0 9108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform -1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform 1 0 33120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _225_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform 1 0 27784 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform -1 0 25576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform -1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform -1 0 27416 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _233_
timestamp 1667941163
transform -1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 11960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform -1 0 31832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform 1 0 30912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 31740 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform -1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _245_
timestamp 1667941163
transform 1 0 35972 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _246_
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform -1 0 29992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _249_
timestamp 1667941163
transform -1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform -1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 17204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _256_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 34040 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform -1 0 31188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 32200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform -1 0 32568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform -1 0 33304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 35328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform -1 0 33488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _267_
timestamp 1667941163
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform -1 0 34684 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform -1 0 33212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform -1 0 32752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform -1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform -1 0 31832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 32752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform -1 0 33488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform -1 0 35144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform -1 0 35144 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _278_
timestamp 1667941163
transform 1 0 14812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform -1 0 33396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform -1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform -1 0 33304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform -1 0 33948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform -1 0 33856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform -1 0 32384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform -1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform -1 0 31832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _289_
timestamp 1667941163
transform 1 0 13892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform -1 0 31832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform -1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform -1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform -1 0 33396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform -1 0 34132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform -1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform -1 0 34132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform -1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform -1 0 33028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _302_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 1667941163
transform 1 0 29348 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _305_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20884 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _306_
timestamp 1667941163
transform 1 0 19596 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _307_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 29256 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 1667941163
transform -1 0 31556 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _311_
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _312_
timestamp 1667941163
transform 1 0 25668 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _313_
timestamp 1667941163
transform 1 0 27324 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1667941163
transform 1 0 20884 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _317_
timestamp 1667941163
transform 1 0 20792 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _318_
timestamp 1667941163
transform 1 0 24564 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _319_
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1667941163
transform 1 0 27324 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1667941163
transform 1 0 26772 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _323_
timestamp 1667941163
transform 1 0 20792 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _324_
timestamp 1667941163
transform -1 0 23920 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _325_
timestamp 1667941163
transform 1 0 27324 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1667941163
transform -1 0 29256 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1667941163
transform -1 0 31556 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _329_
timestamp 1667941163
transform 1 0 26312 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _330_
timestamp 1667941163
transform 1 0 24288 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _331_
timestamp 1667941163
transform -1 0 29624 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 1667941163
transform -1 0 26128 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1667941163
transform 1 0 20884 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _335_
timestamp 1667941163
transform -1 0 22908 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _336_
timestamp 1667941163
transform -1 0 23920 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _337_
timestamp 1667941163
transform -1 0 29992 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _338_
timestamp 1667941163
transform -1 0 28980 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _340_
timestamp 1667941163
transform 1 0 22080 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _341_
timestamp 1667941163
transform 1 0 24196 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _342_
timestamp 1667941163
transform -1 0 21528 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _343_
timestamp 1667941163
transform -1 0 23828 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _351_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1748 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1667941163
transform 1 0 26956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1667941163
transform -1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1667941163
transform -1 0 36156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1667941163
transform -1 0 17848 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1667941163
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _357_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1667941163
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _360_
timestamp 1667941163
transform -1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _361_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _362_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _363_
timestamp 1667941163
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _365_
timestamp 1667941163
transform -1 0 23644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1667941163
transform 1 0 4048 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1667941163
transform -1 0 29992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1667941163
transform -1 0 26864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _369_
timestamp 1667941163
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1667941163
transform 1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1667941163
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1667941163
transform -1 0 35696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _373_
timestamp 1667941163
transform -1 0 26312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _374_
timestamp 1667941163
transform -1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1667941163
transform -1 0 27692 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _376_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1667941163
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1667941163
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1667941163
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1667941163
transform -1 0 22816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1667941163
transform -1 0 23460 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _382_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1667941163
transform -1 0 34960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _384_
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1667941163
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _387_
timestamp 1667941163
transform -1 0 29992 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1667941163
transform -1 0 33672 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _389_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24012 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _390_
timestamp 1667941163
transform 1 0 20976 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _391_
timestamp 1667941163
transform -1 0 24104 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _392_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _393__87 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18584 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _393_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _394_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _395_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18492 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _396_
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _397_
timestamp 1667941163
transform -1 0 26496 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _398_
timestamp 1667941163
transform 1 0 18400 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _399_
timestamp 1667941163
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _400_
timestamp 1667941163
transform -1 0 24748 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _401_
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _402__88
timestamp 1667941163
transform -1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _402_
timestamp 1667941163
transform -1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _403_
timestamp 1667941163
transform 1 0 20056 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _404_
timestamp 1667941163
transform 1 0 27232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _405_
timestamp 1667941163
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _406_
timestamp 1667941163
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _407_
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _408_
timestamp 1667941163
transform 1 0 23460 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _409_
timestamp 1667941163
transform 1 0 27508 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _410_
timestamp 1667941163
transform -1 0 24748 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _411_
timestamp 1667941163
transform -1 0 26312 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _412_
timestamp 1667941163
transform -1 0 26220 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _413_
timestamp 1667941163
transform -1 0 21804 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _414_
timestamp 1667941163
transform -1 0 25300 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _415_
timestamp 1667941163
transform -1 0 28612 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _416__89
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _416_
timestamp 1667941163
transform -1 0 25484 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _417_
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _418_
timestamp 1667941163
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _419_
timestamp 1667941163
transform -1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _420_
timestamp 1667941163
transform 1 0 18768 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _421_
timestamp 1667941163
transform 1 0 20056 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _422_
timestamp 1667941163
transform -1 0 26864 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _423_
timestamp 1667941163
transform 1 0 19596 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _424_
timestamp 1667941163
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _425_
timestamp 1667941163
transform 1 0 25760 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _426_
timestamp 1667941163
transform 1 0 27784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _427_
timestamp 1667941163
transform 1 0 22080 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _428__90
timestamp 1667941163
transform 1 0 25760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _428_
timestamp 1667941163
transform -1 0 25208 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _429_
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _430_
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _431_
timestamp 1667941163
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _432_
timestamp 1667941163
transform -1 0 22724 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _433_
timestamp 1667941163
transform 1 0 25668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _434_
timestamp 1667941163
transform -1 0 27416 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _435_
timestamp 1667941163
transform -1 0 22816 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _436_
timestamp 1667941163
transform 1 0 20976 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _437_
timestamp 1667941163
transform 1 0 25576 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _438_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _439_
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _440_
timestamp 1667941163
transform -1 0 25576 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _440__91
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _441_
timestamp 1667941163
transform -1 0 23736 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _442_
timestamp 1667941163
transform -1 0 22540 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _443_
timestamp 1667941163
transform 1 0 23644 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _444_
timestamp 1667941163
transform -1 0 26220 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _445_
timestamp 1667941163
transform 1 0 26956 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _446_
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _447_
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _448_
timestamp 1667941163
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _449_
timestamp 1667941163
transform -1 0 18492 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _450_
timestamp 1667941163
transform 1 0 19596 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _451_
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _452_
timestamp 1667941163
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _452__92
timestamp 1667941163
transform 1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _453_
timestamp 1667941163
transform -1 0 19320 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _454_
timestamp 1667941163
transform -1 0 20148 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _455_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _456_
timestamp 1667941163
transform -1 0 22816 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _457_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _458_
timestamp 1667941163
transform 1 0 19412 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _459_
timestamp 1667941163
transform 1 0 20424 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _460_
timestamp 1667941163
transform -1 0 25668 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _461_
timestamp 1667941163
transform -1 0 20608 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _462_
timestamp 1667941163
transform 1 0 17204 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _462__93
timestamp 1667941163
transform 1 0 17296 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _463_
timestamp 1667941163
transform -1 0 23736 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _464_
timestamp 1667941163
transform 1 0 22172 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _465_
timestamp 1667941163
transform -1 0 27416 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _466_
timestamp 1667941163
transform 1 0 22724 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _467_
timestamp 1667941163
transform -1 0 23184 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _468_
timestamp 1667941163
transform 1 0 21528 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _469_
timestamp 1667941163
transform -1 0 25944 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 36432 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1667941163
transform -1 0 36432 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform -1 0 36432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 35512 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform -1 0 36432 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform -1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform -1 0 17848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform -1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1667941163
transform -1 0 36432 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform -1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform 1 0 2024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform -1 0 17112 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform -1 0 36432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1667941163
transform -1 0 36432 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1667941163
transform -1 0 24104 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform -1 0 1840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1667941163
transform -1 0 36432 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform -1 0 11224 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform -1 0 36432 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 26312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform -1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1667941163
transform -1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 36064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 36064 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform -1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform -1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 36064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 28796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform 1 0 34868 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform 1 0 36064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform -1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform -1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform 1 0 36064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 3128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 36064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 33948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 36064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 36064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 36064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 36064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 36064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform -1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 36064 0 1 18496
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 0 nsew signal tristate
flabel metal3 s 37200 25848 37800 25968 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 1 nsew signal tristate
flabel metal3 s 37200 35368 37800 35488 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 2 nsew signal tristate
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
port 3 nsew signal tristate
flabel metal3 s 37200 31288 37800 31408 0 FreeSans 480 0 0 0 ccff_head
port 4 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal3 s 37200 7488 37800 7608 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 37200 27888 37800 28008 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 37200 38768 37800 38888 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 37200 23808 37800 23928 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 17406 39200 17462 39800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal3 s 37200 2048 37800 2168 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal3 s 37200 14968 37800 15088 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal3 s 37200 29928 37800 30048 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal3 s 37200 17008 37800 17128 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 37200 12928 37800 13048 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal2 s 15474 200 15530 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal3 s 37200 33328 37800 33448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal3 s 37200 10888 37800 11008 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal3 s 37200 5448 37800 5568 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal3 s 37200 8 37800 128 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal3 s 37200 9528 37800 9648 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal3 s 37200 36728 37800 36848 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal3 s 37200 4088 37800 4208 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal3 s 37200 20408 37800 20528 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal3 s 200 16328 800 16448 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal3 s 37200 22448 37800 22568 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 pReset
port 82 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 prog_clk
port 83 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 84 nsew signal tristate
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 85 nsew signal tristate
flabel metal3 s 37200 18368 37800 18488 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 86 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 87 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 87 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 88 nsew ground bidirectional
rlabel metal1 18998 37536 18998 37536 0 vccd1
rlabel metal1 18998 36992 18998 36992 0 vssd1
rlabel metal2 33902 3196 33902 3196 0 _000_
rlabel metal2 33718 3502 33718 3502 0 _001_
rlabel metal1 30820 5202 30820 5202 0 _002_
rlabel metal2 32062 6800 32062 6800 0 _003_
rlabel via2 32430 5219 32430 5219 0 _004_
rlabel metal2 31786 7888 31786 7888 0 _005_
rlabel metal1 34960 6086 34960 6086 0 _006_
rlabel metal1 33626 6834 33626 6834 0 _007_
rlabel metal1 30873 3434 30873 3434 0 _008_
rlabel metal1 33166 5882 33166 5882 0 _009_
rlabel metal2 34546 6562 34546 6562 0 _010_
rlabel metal1 29355 4590 29355 4590 0 _011_
rlabel metal2 32614 6630 32614 6630 0 _012_
rlabel metal2 31050 7718 31050 7718 0 _013_
rlabel metal2 33074 4454 33074 4454 0 _014_
rlabel metal1 30774 4998 30774 4998 0 _015_
rlabel metal2 32614 4862 32614 4862 0 _016_
rlabel via2 31602 3621 31602 3621 0 _017_
rlabel metal2 33166 3774 33166 3774 0 _018_
rlabel metal2 32798 4488 32798 4488 0 _019_
rlabel metal1 29401 8874 29401 8874 0 _020_
rlabel metal1 32384 4114 32384 4114 0 _021_
rlabel metal2 30406 5848 30406 5848 0 _022_
rlabel metal2 31878 7276 31878 7276 0 _023_
rlabel metal1 31878 7412 31878 7412 0 _024_
rlabel metal2 30774 4828 30774 4828 0 _025_
rlabel metal2 31142 6154 31142 6154 0 _026_
rlabel metal1 28711 7854 28711 7854 0 _027_
rlabel metal1 31556 6426 31556 6426 0 _028_
rlabel metal2 33534 6494 33534 6494 0 _029_
rlabel metal1 31602 3026 31602 3026 0 _030_
rlabel metal1 32844 3162 32844 3162 0 _031_
rlabel metal2 32062 3264 32062 3264 0 _032_
rlabel via2 33074 5083 33074 5083 0 _033_
rlabel via2 33258 4539 33258 4539 0 _034_
rlabel metal1 33396 5814 33396 5814 0 _035_
rlabel metal2 29762 3026 29762 3026 0 _036_
rlabel metal1 32867 3434 32867 3434 0 _037_
rlabel metal2 32706 3978 32706 3978 0 _038_
rlabel metal2 32798 8653 32798 8653 0 _039_
rlabel metal1 14996 5066 14996 5066 0 _040_
rlabel metal2 21482 4318 21482 4318 0 _041_
rlabel metal1 32522 5236 32522 5236 0 _042_
rlabel metal2 31786 4471 31786 4471 0 _043_
rlabel metal2 31878 6528 31878 6528 0 _044_
rlabel metal2 31786 3111 31786 3111 0 _045_
rlabel via2 26174 12835 26174 12835 0 _046_
rlabel metal1 20930 13226 20930 13226 0 _047_
rlabel metal1 23322 7514 23322 7514 0 _048_
rlabel metal1 19642 6664 19642 6664 0 _049_
rlabel metal1 20976 12954 20976 12954 0 _050_
rlabel metal1 18906 13498 18906 13498 0 _051_
rlabel metal2 18170 10472 18170 10472 0 _052_
rlabel metal2 19090 7582 19090 7582 0 _053_
rlabel metal2 26128 12614 26128 12614 0 _054_
rlabel metal1 18262 8534 18262 8534 0 _055_
rlabel metal1 17894 12818 17894 12818 0 _056_
rlabel metal1 24610 8058 24610 8058 0 _057_
rlabel metal2 28106 11509 28106 11509 0 _058_
rlabel metal1 23046 17544 23046 17544 0 _059_
rlabel metal2 20746 8500 20746 8500 0 _060_
rlabel metal1 27876 12886 27876 12886 0 _061_
rlabel metal1 26680 14994 26680 14994 0 _062_
rlabel metal1 23598 14484 23598 14484 0 _063_
rlabel metal1 23736 16626 23736 16626 0 _064_
rlabel metal1 24288 14926 24288 14926 0 _065_
rlabel metal1 29026 14008 29026 14008 0 _066_
rlabel metal1 24518 17272 24518 17272 0 _067_
rlabel metal1 26128 16082 26128 16082 0 _068_
rlabel metal1 27554 14450 27554 14450 0 _069_
rlabel metal1 21574 14280 21574 14280 0 _070_
rlabel metal1 27002 10234 27002 10234 0 _071_
rlabel metal2 28290 12988 28290 12988 0 _072_
rlabel metal1 26588 15062 26588 15062 0 _073_
rlabel metal1 19826 15130 19826 15130 0 _074_
rlabel metal1 20976 14994 20976 14994 0 _075_
rlabel metal2 18170 11492 18170 11492 0 _076_
rlabel metal2 18998 9996 18998 9996 0 _077_
rlabel metal1 19780 10710 19780 10710 0 _078_
rlabel metal2 26634 16728 26634 16728 0 _079_
rlabel metal1 20010 14994 20010 14994 0 _080_
rlabel metal2 18446 9180 18446 9180 0 _081_
rlabel metal1 27512 9962 27512 9962 0 _082_
rlabel metal1 29026 14518 29026 14518 0 _083_
rlabel metal1 23000 15062 23000 15062 0 _084_
rlabel metal1 27968 14926 27968 14926 0 _085_
rlabel metal2 18814 11560 18814 11560 0 _086_
rlabel metal2 19642 5882 19642 5882 0 _087_
rlabel metal2 20884 15402 20884 15402 0 _088_
rlabel metal1 22402 13498 22402 13498 0 _089_
rlabel metal1 25898 10744 25898 10744 0 _090_
rlabel metal1 29992 14042 29992 14042 0 _091_
rlabel metal2 24702 11560 24702 11560 0 _092_
rlabel metal1 21666 11016 21666 11016 0 _093_
rlabel metal2 29854 12002 29854 12002 0 _094_
rlabel metal2 27922 10166 27922 10166 0 _095_
rlabel metal1 29095 11594 29095 11594 0 _096_
rlabel metal1 28382 15130 28382 15130 0 _097_
rlabel metal1 23506 13192 23506 13192 0 _098_
rlabel metal1 22310 12104 22310 12104 0 _099_
rlabel metal1 24610 12886 24610 12886 0 _100_
rlabel metal2 27738 13617 27738 13617 0 _101_
rlabel metal1 27600 11050 27600 11050 0 _102_
rlabel metal1 22448 14586 22448 14586 0 _103_
rlabel metal1 20746 13974 20746 13974 0 _104_
rlabel metal1 24150 14586 24150 14586 0 _105_
rlabel metal1 17848 6834 17848 6834 0 _106_
rlabel metal1 19872 5338 19872 5338 0 _107_
rlabel metal2 19182 12988 19182 12988 0 _108_
rlabel metal2 17618 12002 17618 12002 0 _109_
rlabel metal2 18630 6052 18630 6052 0 _110_
rlabel metal1 19366 7854 19366 7854 0 _111_
rlabel metal1 18354 12614 18354 12614 0 _112_
rlabel metal1 22402 12886 22402 12886 0 _113_
rlabel metal1 19090 10234 19090 10234 0 _114_
rlabel metal2 17526 11696 17526 11696 0 _115_
rlabel metal1 18400 6766 18400 6766 0 _116_
rlabel metal1 26312 12886 26312 12886 0 _117_
rlabel metal1 20378 8840 20378 8840 0 _118_
rlabel metal2 16790 5032 16790 5032 0 _119_
rlabel metal1 27784 11662 27784 11662 0 _120_
rlabel metal2 23966 9554 23966 9554 0 _121_
rlabel metal1 27600 13158 27600 13158 0 _122_
rlabel metal1 26404 9418 26404 9418 0 _123_
rlabel metal1 26220 9622 26220 9622 0 _124_
rlabel metal2 21758 9826 21758 9826 0 _125_
rlabel metal1 26772 14042 26772 14042 0 _126_
rlabel metal3 1188 31348 1188 31348 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
rlabel metal3 36532 25908 36532 25908 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
rlabel via2 36294 35445 36294 35445 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal3 1188 14348 1188 14348 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
rlabel via2 36386 31365 36386 31365 0 ccff_head
rlabel metal2 13570 1520 13570 1520 0 ccff_tail
rlabel via2 36386 7531 36386 7531 0 chanx_left_in[0]
rlabel metal1 8464 2278 8464 2278 0 chanx_left_in[10]
rlabel metal2 36294 27999 36294 27999 0 chanx_left_in[11]
rlabel metal1 19182 2414 19182 2414 0 chanx_left_in[12]
rlabel metal2 1610 21913 1610 21913 0 chanx_left_in[13]
rlabel metal2 35558 38063 35558 38063 0 chanx_left_in[14]
rlabel via2 36386 23851 36386 23851 0 chanx_left_in[15]
rlabel metal1 36248 3502 36248 3502 0 chanx_left_in[16]
rlabel metal1 5290 37230 5290 37230 0 chanx_left_in[17]
rlabel metal1 17572 37230 17572 37230 0 chanx_left_in[18]
rlabel metal1 21344 37434 21344 37434 0 chanx_left_in[1]
rlabel metal1 34914 3094 34914 3094 0 chanx_left_in[2]
rlabel metal1 35282 2414 35282 2414 0 chanx_left_in[3]
rlabel metal2 36386 15249 36386 15249 0 chanx_left_in[4]
rlabel metal1 34040 2414 34040 2414 0 chanx_left_in[5]
rlabel metal1 24610 37230 24610 37230 0 chanx_left_in[6]
rlabel metal1 2070 37230 2070 37230 0 chanx_left_in[7]
rlabel metal1 16721 37230 16721 37230 0 chanx_left_in[8]
rlabel via2 1610 23851 1610 23851 0 chanx_left_in[9]
rlabel via2 36294 30005 36294 30005 0 chanx_left_out[0]
rlabel metal3 1188 1428 1188 1428 0 chanx_left_out[10]
rlabel metal3 1188 29308 1188 29308 0 chanx_left_out[11]
rlabel metal1 28474 37094 28474 37094 0 chanx_left_out[12]
rlabel metal3 1188 3468 1188 3468 0 chanx_left_out[13]
rlabel metal1 34960 36890 34960 36890 0 chanx_left_out[14]
rlabel via2 36294 17051 36294 17051 0 chanx_left_out[15]
rlabel metal1 19504 37094 19504 37094 0 chanx_left_out[16]
rlabel metal1 22678 2822 22678 2822 0 chanx_left_out[17]
rlabel metal3 1188 36788 1188 36788 0 chanx_left_out[18]
rlabel metal1 26910 37094 26910 37094 0 chanx_left_out[1]
rlabel metal2 36294 13073 36294 13073 0 chanx_left_out[2]
rlabel metal1 1472 37434 1472 37434 0 chanx_left_out[3]
rlabel metal1 30176 2822 30176 2822 0 chanx_left_out[4]
rlabel metal2 15502 1520 15502 1520 0 chanx_left_out[5]
rlabel metal3 1188 6868 1188 6868 0 chanx_left_out[6]
rlabel via2 36294 33371 36294 33371 0 chanx_left_out[7]
rlabel metal3 1188 8908 1188 8908 0 chanx_left_out[8]
rlabel metal2 3266 1520 3266 1520 0 chanx_left_out[9]
rlabel metal1 10442 2346 10442 2346 0 chanx_right_in[0]
rlabel metal1 32246 2414 32246 2414 0 chanx_right_in[10]
rlabel metal2 36294 10999 36294 10999 0 chanx_right_in[11]
rlabel metal2 36386 5593 36386 5593 0 chanx_right_in[12]
rlabel metal1 24104 3570 24104 3570 0 chanx_right_in[13]
rlabel metal1 2530 36346 2530 36346 0 chanx_right_in[14]
rlabel metal2 36386 1513 36386 1513 0 chanx_right_in[15]
rlabel metal1 10764 37298 10764 37298 0 chanx_right_in[16]
rlabel via2 36386 9605 36386 9605 0 chanx_right_in[17]
rlabel via2 1610 25245 1610 25245 0 chanx_right_in[18]
rlabel metal2 26450 4080 26450 4080 0 chanx_right_in[1]
rlabel via2 1610 18411 1610 18411 0 chanx_right_in[2]
rlabel metal2 7130 38260 7130 38260 0 chanx_right_in[3]
rlabel metal1 14306 37230 14306 37230 0 chanx_right_in[4]
rlabel metal2 1702 32759 1702 32759 0 chanx_right_in[5]
rlabel metal1 2346 2380 2346 2380 0 chanx_right_in[6]
rlabel via2 1610 19805 1610 19805 0 chanx_right_in[7]
rlabel metal1 12512 37230 12512 37230 0 chanx_right_in[8]
rlabel metal1 22770 37230 22770 37230 0 chanx_right_in[9]
rlabel metal1 33626 37094 33626 37094 0 chanx_right_out[0]
rlabel metal3 1188 27268 1188 27268 0 chanx_right_out[10]
rlabel metal2 5198 1520 5198 1520 0 chanx_right_out[11]
rlabel metal2 1334 1520 1334 1520 0 chanx_right_out[12]
rlabel metal1 36524 36346 36524 36346 0 chanx_right_out[13]
rlabel metal3 1188 5508 1188 5508 0 chanx_right_out[14]
rlabel metal2 17434 1520 17434 1520 0 chanx_right_out[15]
rlabel metal2 36294 36839 36294 36839 0 chanx_right_out[16]
rlabel metal2 36294 4301 36294 4301 0 chanx_right_out[17]
rlabel metal3 1188 10948 1188 10948 0 chanx_right_out[18]
rlabel metal2 36294 20621 36294 20621 0 chanx_right_out[1]
rlabel metal2 6486 1520 6486 1520 0 chanx_right_out[2]
rlabel metal2 11638 1520 11638 1520 0 chanx_right_out[3]
rlabel via2 1702 16405 1702 16405 0 chanx_right_out[4]
rlabel via2 36294 22491 36294 22491 0 chanx_right_out[5]
rlabel metal2 20654 1520 20654 1520 0 chanx_right_out[6]
rlabel metal1 32154 37094 32154 37094 0 chanx_right_out[7]
rlabel metal1 29808 37094 29808 37094 0 chanx_right_out[8]
rlabel metal1 4048 37094 4048 37094 0 chanx_right_out[9]
rlabel metal2 17802 10336 17802 10336 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal1 19872 13158 19872 13158 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal2 20286 6494 20286 6494 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal2 24794 5457 24794 5457 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal1 18078 7820 18078 7820 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal1 18262 10098 18262 10098 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal1 29302 14382 29302 14382 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel metal1 27738 6630 27738 6630 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal1 34822 3706 34822 3706 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel metal1 29946 3638 29946 3638 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal1 28980 5338 28980 5338 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal1 27922 2618 27922 2618 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal1 21666 2618 21666 2618 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal1 24426 9486 24426 9486 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal2 24058 7786 24058 7786 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal2 27094 6494 27094 6494 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal2 17250 6205 17250 6205 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal1 21390 2890 21390 2890 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal1 20286 16626 20286 16626 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal1 19044 14994 19044 14994 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal1 20562 17136 20562 17136 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal2 19090 10268 19090 10268 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal2 23782 8398 23782 8398 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 27646 7820 27646 7820 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal1 29348 13702 29348 13702 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal1 20792 5610 20792 5610 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal1 18170 13362 18170 13362 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal1 29256 2550 29256 2550 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal1 30544 2618 30544 2618 0 mem_top_ipin_1.DFFR_4_.Q
rlabel metal1 29210 2618 29210 2618 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal2 21850 14144 21850 14144 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal1 28658 12784 28658 12784 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal1 29670 13838 29670 13838 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal2 31510 8466 31510 8466 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal2 29762 8228 29762 8228 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal1 27738 9554 27738 9554 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal1 17802 6766 17802 6766 0 mem_top_ipin_3.DFFR_0_.Q
rlabel metal1 18216 13294 18216 13294 0 mem_top_ipin_3.DFFR_1_.Q
rlabel metal1 20976 8806 20976 8806 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal1 22632 3638 22632 3638 0 mem_top_ipin_3.DFFR_3_.Q
rlabel via2 22034 6307 22034 6307 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal2 30866 14450 30866 14450 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal2 23414 13872 23414 13872 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 24656 13838 24656 13838 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal2 18538 7514 18538 7514 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 19136 6290 19136 6290 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal1 21022 7956 21022 7956 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal1 18078 12750 18078 12750 0 mux_bottom_ipin_0.INVTX1_6_.out
rlabel metal1 17848 14042 17848 14042 0 mux_bottom_ipin_0.INVTX1_7_.out
rlabel metal1 23414 13804 23414 13804 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19090 8296 19090 8296 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 19458 14144 19458 14144 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 6348 29614 6348 29614 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 25898 16252 25898 16252 0 mux_bottom_ipin_1.INVTX1_2_.out
rlabel metal1 27692 15878 27692 15878 0 mux_bottom_ipin_1.INVTX1_3_.out
rlabel metal1 23276 14994 23276 14994 0 mux_bottom_ipin_1.INVTX1_4_.out
rlabel metal2 21390 16796 21390 16796 0 mux_bottom_ipin_1.INVTX1_5_.out
rlabel metal2 24610 17374 24610 17374 0 mux_bottom_ipin_1.INVTX1_6_.out
rlabel metal1 19136 5338 19136 5338 0 mux_bottom_ipin_1.INVTX1_7_.out
rlabel metal1 24794 14246 24794 14246 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23690 14858 23690 14858 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal3 24656 12716 24656 12716 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 32453 17646 32453 17646 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 18768 8942 18768 8942 0 mux_bottom_ipin_2.INVTX1_2_.out
rlabel metal1 19458 11628 19458 11628 0 mux_bottom_ipin_2.INVTX1_3_.out
rlabel metal1 24150 12274 24150 12274 0 mux_bottom_ipin_2.INVTX1_4_.out
rlabel metal1 21850 11152 21850 11152 0 mux_bottom_ipin_2.INVTX1_5_.out
rlabel metal1 26082 13838 26082 13838 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 21574 9078 21574 9078 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 7958 10030 7958 10030 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 18814 7514 18814 7514 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal1 14674 29478 14674 29478 0 mux_top_ipin_0.INVTX1_3_.out
rlabel metal2 9246 18462 9246 18462 0 mux_top_ipin_0.INVTX1_4_.out
rlabel metal2 20746 15810 20746 15810 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal2 26726 17340 26726 17340 0 mux_top_ipin_0.INVTX1_6_.out
rlabel metal1 30084 13226 30084 13226 0 mux_top_ipin_0.INVTX1_7_.out
rlabel metal1 20102 10574 20102 10574 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20700 15062 20700 15062 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal3 26358 13260 26358 13260 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 2300 31314 2300 31314 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22356 15538 22356 15538 0 mux_top_ipin_1.INVTX1_2_.out
rlabel metal1 23552 11866 23552 11866 0 mux_top_ipin_1.INVTX1_3_.out
rlabel metal1 19780 11662 19780 11662 0 mux_top_ipin_1.INVTX1_4_.out
rlabel metal2 17894 4828 17894 4828 0 mux_top_ipin_1.INVTX1_5_.out
rlabel metal1 27508 14314 27508 14314 0 mux_top_ipin_1.INVTX1_6_.out
rlabel metal1 19964 31110 19964 31110 0 mux_top_ipin_1.INVTX1_7_.out
rlabel metal1 21850 15402 21850 15402 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20286 5678 20286 5678 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 24426 15402 24426 15402 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 28566 16558 28566 16558 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 26082 13430 26082 13430 0 mux_top_ipin_2.INVTX1_2_.out
rlabel metal1 19734 13974 19734 13974 0 mux_top_ipin_2.INVTX1_3_.out
rlabel metal1 23184 16014 23184 16014 0 mux_top_ipin_2.INVTX1_6_.out
rlabel metal1 25438 10234 25438 10234 0 mux_top_ipin_2.INVTX1_7_.out
rlabel metal2 24334 14042 24334 14042 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 22954 13532 22954 13532 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 25208 15538 25208 15538 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 35949 35054 35949 35054 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 21390 12818 21390 12818 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19366 7718 19366 7718 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19826 12614 19826 12614 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 2806 12818 2806 12818 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 36294 31858 36294 31858 0 net1
rlabel metal2 5566 27676 5566 27676 0 net10
rlabel metal1 17296 37298 17296 37298 0 net11
rlabel metal1 23920 37366 23920 37366 0 net12
rlabel via2 34822 2907 34822 2907 0 net13
rlabel metal1 17986 4726 17986 4726 0 net14
rlabel metal1 12466 16014 12466 16014 0 net15
rlabel metal1 34178 2618 34178 2618 0 net16
rlabel metal2 24886 36589 24886 36589 0 net17
rlabel metal2 23230 36958 23230 36958 0 net18
rlabel metal1 22586 36788 22586 36788 0 net19
rlabel metal1 35995 7922 35995 7922 0 net2
rlabel metal1 3266 24174 3266 24174 0 net20
rlabel metal2 10626 2108 10626 2108 0 net21
rlabel metal1 32614 2380 32614 2380 0 net22
rlabel metal2 36110 9860 36110 9860 0 net23
rlabel metal1 34638 5746 34638 5746 0 net24
rlabel metal1 10534 3468 10534 3468 0 net25
rlabel metal1 1794 36040 1794 36040 0 net26
rlabel metal2 36110 4963 36110 4963 0 net27
rlabel metal1 19090 36754 19090 36754 0 net28
rlabel metal1 27186 10064 27186 10064 0 net29
rlabel metal1 5198 23086 5198 23086 0 net3
rlabel metal2 1886 23086 1886 23086 0 net30
rlabel metal1 27508 26282 27508 26282 0 net31
rlabel metal1 2300 18666 2300 18666 0 net32
rlabel metal2 7498 36992 7498 36992 0 net33
rlabel metal1 16146 12342 16146 12342 0 net34
rlabel metal1 9844 32742 9844 32742 0 net35
rlabel metal2 1978 6528 1978 6528 0 net36
rlabel metal2 21390 18836 21390 18836 0 net37
rlabel metal1 6831 23698 6831 23698 0 net38
rlabel metal1 22724 37298 22724 37298 0 net39
rlabel metal2 36202 20128 36202 20128 0 net4
rlabel metal1 11546 37434 11546 37434 0 net40
rlabel metal1 1932 31450 1932 31450 0 net41
rlabel metal2 35374 22644 35374 22644 0 net42
rlabel metal2 36110 35462 36110 35462 0 net43
rlabel metal1 2162 12954 2162 12954 0 net44
rlabel metal1 14582 2448 14582 2448 0 net45
rlabel metal2 35650 30124 35650 30124 0 net46
rlabel metal1 4393 3026 4393 3026 0 net47
rlabel metal1 1932 29614 1932 29614 0 net48
rlabel metal1 28796 37230 28796 37230 0 net49
rlabel metal1 19274 2618 19274 2618 0 net5
rlabel metal1 4393 3502 4393 3502 0 net50
rlabel metal1 22678 36720 22678 36720 0 net51
rlabel metal2 36110 16150 36110 16150 0 net52
rlabel metal2 18906 37060 18906 37060 0 net53
rlabel metal1 23046 3026 23046 3026 0 net54
rlabel metal1 1840 36754 1840 36754 0 net55
rlabel metal1 27002 37230 27002 37230 0 net56
rlabel metal1 36110 13328 36110 13328 0 net57
rlabel metal1 3588 36890 3588 36890 0 net58
rlabel via2 32338 3043 32338 3043 0 net59
rlabel metal1 27784 31314 27784 31314 0 net6
rlabel metal1 16652 2414 16652 2414 0 net60
rlabel metal1 1840 6426 1840 6426 0 net61
rlabel metal2 35558 33388 35558 33388 0 net62
rlabel metal1 4508 9146 4508 9146 0 net63
rlabel metal1 4508 2414 4508 2414 0 net64
rlabel metal1 33810 36550 33810 36550 0 net65
rlabel metal1 4232 23290 4232 23290 0 net66
rlabel metal2 5566 6970 5566 6970 0 net67
rlabel metal2 4646 2652 4646 2652 0 net68
rlabel metal1 34224 36142 34224 36142 0 net69
rlabel metal2 35834 36555 35834 36555 0 net7
rlabel metal1 2116 5678 2116 5678 0 net70
rlabel metal2 18354 2176 18354 2176 0 net71
rlabel metal1 36064 36754 36064 36754 0 net72
rlabel metal1 36018 4590 36018 4590 0 net73
rlabel metal2 1886 11594 1886 11594 0 net74
rlabel metal1 35995 20910 35995 20910 0 net75
rlabel metal1 10534 2448 10534 2448 0 net76
rlabel metal1 12236 2414 12236 2414 0 net77
rlabel metal2 11730 16388 11730 16388 0 net78
rlabel metal2 36110 21046 36110 21046 0 net79
rlabel metal1 33258 24174 33258 24174 0 net8
rlabel metal2 21022 2587 21022 2587 0 net80
rlabel metal1 24978 36584 24978 36584 0 net81
rlabel metal1 25070 36652 25070 36652 0 net82
rlabel metal2 4002 34612 4002 34612 0 net83
rlabel metal2 5658 11560 5658 11560 0 net84
rlabel metal1 4370 29818 4370 29818 0 net85
rlabel metal1 33902 17850 33902 17850 0 net86
rlabel metal1 19320 14450 19320 14450 0 net87
rlabel metal2 23138 17952 23138 17952 0 net88
rlabel metal2 25346 14977 25346 14977 0 net89
rlabel metal1 35742 3638 35742 3638 0 net9
rlabel metal1 25438 16150 25438 16150 0 net90
rlabel metal1 26772 15130 26772 15130 0 net91
rlabel metal2 18170 12036 18170 12036 0 net92
rlabel metal2 17342 4896 17342 4896 0 net93
rlabel metal1 9154 37230 9154 37230 0 pReset
rlabel metal2 36018 2992 36018 2992 0 prog_clk
rlabel metal3 1188 12308 1188 12308 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
rlabel metal3 1188 34748 1188 34748 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel metal2 36294 18513 36294 18513 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
<< properties >>
string FIXED_BBOX 0 0 38000 40000
<< end >>
