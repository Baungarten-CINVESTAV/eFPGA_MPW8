magic
tech sky130A
magscale 1 2
timestamp 1672417963
<< viali >>
rect 2513 27557 2547 27591
rect 3249 27557 3283 27591
rect 3985 27557 4019 27591
rect 7849 27557 7883 27591
rect 10609 27557 10643 27591
rect 13645 27557 13679 27591
rect 15117 27557 15151 27591
rect 17049 27557 17083 27591
rect 18337 27557 18371 27591
rect 19441 27557 19475 27591
rect 20913 27557 20947 27591
rect 24593 27557 24627 27591
rect 27997 27557 28031 27591
rect 2329 27421 2363 27455
rect 3433 27421 3467 27455
rect 4169 27421 4203 27455
rect 5457 27421 5491 27455
rect 6745 27421 6779 27455
rect 8033 27421 8067 27455
rect 9321 27421 9355 27455
rect 10425 27421 10459 27455
rect 11897 27421 11931 27455
rect 12541 27421 12575 27455
rect 13461 27421 13495 27455
rect 14289 27421 14323 27455
rect 14933 27421 14967 27455
rect 15853 27421 15887 27455
rect 16865 27421 16899 27455
rect 18153 27421 18187 27455
rect 19625 27421 19659 27455
rect 20085 27421 20119 27455
rect 20729 27421 20763 27455
rect 22845 27421 22879 27455
rect 23305 27421 23339 27455
rect 24777 27421 24811 27455
rect 25421 27421 25455 27455
rect 26065 27421 26099 27455
rect 27353 27421 27387 27455
rect 27813 27421 27847 27455
rect 1685 27353 1719 27387
rect 1869 27353 1903 27387
rect 5273 27285 5307 27319
rect 6561 27285 6595 27319
rect 9137 27285 9171 27319
rect 11713 27285 11747 27319
rect 12357 27285 12391 27319
rect 14381 27285 14415 27319
rect 15669 27285 15703 27319
rect 20177 27285 20211 27319
rect 22017 27285 22051 27319
rect 22661 27285 22695 27319
rect 23397 27285 23431 27319
rect 25237 27285 25271 27319
rect 25881 27285 25915 27319
rect 27169 27285 27203 27319
rect 1777 27081 1811 27115
rect 3893 27081 3927 27115
rect 13185 27081 13219 27115
rect 27537 27081 27571 27115
rect 28273 27081 28307 27115
rect 20729 27013 20763 27047
rect 1593 26945 1627 26979
rect 2513 26945 2547 26979
rect 3157 26945 3191 26979
rect 4077 26945 4111 26979
rect 13369 26945 13403 26979
rect 14013 26945 14047 26979
rect 14473 26945 14507 26979
rect 15117 26945 15151 26979
rect 16865 26945 16899 26979
rect 17785 26945 17819 26979
rect 18613 26945 18647 26979
rect 19257 26945 19291 26979
rect 21373 26945 21407 26979
rect 22017 26945 22051 26979
rect 23305 26945 23339 26979
rect 23765 26945 23799 26979
rect 24409 26945 24443 26979
rect 25513 26945 25547 26979
rect 25973 26945 26007 26979
rect 27353 26945 27387 26979
rect 28089 26945 28123 26979
rect 11713 26877 11747 26911
rect 15301 26877 15335 26911
rect 17049 26877 17083 26911
rect 20085 26877 20119 26911
rect 20269 26877 20303 26911
rect 22201 26877 22235 26911
rect 2329 26809 2363 26843
rect 18429 26809 18463 26843
rect 2973 26741 3007 26775
rect 13829 26741 13863 26775
rect 14565 26741 14599 26775
rect 15761 26741 15795 26775
rect 17877 26741 17911 26775
rect 19073 26741 19107 26775
rect 21189 26741 21223 26775
rect 22569 26741 22603 26775
rect 23121 26741 23155 26775
rect 23857 26741 23891 26775
rect 24501 26741 24535 26775
rect 25329 26741 25363 26775
rect 26065 26741 26099 26775
rect 1593 26537 1627 26571
rect 4261 26537 4295 26571
rect 4905 26537 4939 26571
rect 10701 26537 10735 26571
rect 18797 26537 18831 26571
rect 19441 26537 19475 26571
rect 20177 26537 20211 26571
rect 20729 26537 20763 26571
rect 21373 26537 21407 26571
rect 22661 26537 22695 26571
rect 27353 26537 27387 26571
rect 28273 26537 28307 26571
rect 11345 26469 11379 26503
rect 15669 26469 15703 26503
rect 16865 26469 16899 26503
rect 23305 26469 23339 26503
rect 26065 26469 26099 26503
rect 15209 26401 15243 26435
rect 16681 26401 16715 26435
rect 1777 26333 1811 26367
rect 4169 26333 4203 26367
rect 5089 26333 5123 26367
rect 10885 26333 10919 26367
rect 11529 26333 11563 26367
rect 11989 26333 12023 26367
rect 12725 26333 12759 26367
rect 13369 26333 13403 26367
rect 14381 26333 14415 26367
rect 15025 26333 15059 26367
rect 16497 26333 16531 26367
rect 18061 26333 18095 26367
rect 18705 26333 18739 26367
rect 19625 26333 19659 26367
rect 20085 26333 20119 26367
rect 20913 26333 20947 26367
rect 21557 26333 21591 26367
rect 22201 26333 22235 26367
rect 22845 26333 22879 26367
rect 23489 26333 23523 26367
rect 25145 26333 25179 26367
rect 26249 26333 26283 26367
rect 26893 26333 26927 26367
rect 27537 26333 27571 26367
rect 28089 26333 28123 26367
rect 12817 26265 12851 26299
rect 12081 26197 12115 26231
rect 13461 26197 13495 26231
rect 18153 26197 18187 26231
rect 22017 26197 22051 26231
rect 24961 26197 24995 26231
rect 26709 26197 26743 26231
rect 4997 25993 5031 26027
rect 15117 25993 15151 26027
rect 27537 25993 27571 26027
rect 11805 25925 11839 25959
rect 11897 25925 11931 25959
rect 13369 25925 13403 25959
rect 4905 25857 4939 25891
rect 8125 25857 8159 25891
rect 10609 25857 10643 25891
rect 14565 25857 14599 25891
rect 15025 25857 15059 25891
rect 17049 25857 17083 25891
rect 17877 25857 17911 25891
rect 18521 25857 18555 25891
rect 19625 25857 19659 25891
rect 21005 25857 21039 25891
rect 22017 25857 22051 25891
rect 24409 25857 24443 25891
rect 25605 25857 25639 25891
rect 27721 25857 27755 25891
rect 28365 25857 28399 25891
rect 12081 25789 12115 25823
rect 13277 25789 13311 25823
rect 13553 25789 13587 25823
rect 15669 25789 15703 25823
rect 15853 25789 15887 25823
rect 18705 25789 18739 25823
rect 22661 25789 22695 25823
rect 22845 25789 22879 25823
rect 8217 25721 8251 25755
rect 16313 25721 16347 25755
rect 23305 25721 23339 25755
rect 10425 25653 10459 25687
rect 14381 25653 14415 25687
rect 17141 25653 17175 25687
rect 17969 25653 18003 25687
rect 18889 25653 18923 25687
rect 20821 25653 20855 25687
rect 22109 25653 22143 25687
rect 24225 25653 24259 25687
rect 25697 25653 25731 25687
rect 28181 25653 28215 25687
rect 12265 25449 12299 25483
rect 14381 25449 14415 25483
rect 17601 25449 17635 25483
rect 19901 25449 19935 25483
rect 21557 25449 21591 25483
rect 25237 25449 25271 25483
rect 27905 25449 27939 25483
rect 11713 25381 11747 25415
rect 17049 25381 17083 25415
rect 21189 25313 21223 25347
rect 21373 25313 21407 25347
rect 22845 25313 22879 25347
rect 23581 25313 23615 25347
rect 26617 25313 26651 25347
rect 11161 25245 11195 25279
rect 11621 25245 11655 25279
rect 12449 25245 12483 25279
rect 13093 25245 13127 25279
rect 13553 25245 13587 25279
rect 14565 25245 14599 25279
rect 16497 25245 16531 25279
rect 16681 25245 16715 25279
rect 17785 25245 17819 25279
rect 18429 25245 18463 25279
rect 19809 25245 19843 25279
rect 20453 25245 20487 25279
rect 22753 25245 22787 25279
rect 23397 25245 23431 25279
rect 24777 25245 24811 25279
rect 25421 25245 25455 25279
rect 25881 25245 25915 25279
rect 26525 25245 26559 25279
rect 27813 25245 27847 25279
rect 15117 25177 15151 25211
rect 15209 25177 15243 25211
rect 15761 25177 15795 25211
rect 20545 25177 20579 25211
rect 24041 25177 24075 25211
rect 25973 25177 26007 25211
rect 10333 25109 10367 25143
rect 10977 25109 11011 25143
rect 12909 25109 12943 25143
rect 13645 25109 13679 25143
rect 18245 25109 18279 25143
rect 24593 25109 24627 25143
rect 18153 24905 18187 24939
rect 17141 24837 17175 24871
rect 25421 24837 25455 24871
rect 1777 24769 1811 24803
rect 9229 24769 9263 24803
rect 9873 24769 9907 24803
rect 10517 24769 10551 24803
rect 11713 24769 11747 24803
rect 13001 24769 13035 24803
rect 13921 24769 13955 24803
rect 14105 24769 14139 24803
rect 18337 24769 18371 24803
rect 18981 24769 19015 24803
rect 19441 24769 19475 24803
rect 20269 24769 20303 24803
rect 20729 24769 20763 24803
rect 23581 24769 23615 24803
rect 25145 24769 25179 24803
rect 25881 24769 25915 24803
rect 27261 24769 27295 24803
rect 28181 24769 28215 24803
rect 10977 24701 11011 24735
rect 12817 24701 12851 24735
rect 17049 24701 17083 24735
rect 22017 24701 22051 24735
rect 22201 24701 22235 24735
rect 23765 24701 23799 24735
rect 9045 24633 9079 24667
rect 10333 24633 10367 24667
rect 17601 24633 17635 24667
rect 22661 24633 22695 24667
rect 1593 24565 1627 24599
rect 9689 24565 9723 24599
rect 11805 24565 11839 24599
rect 13461 24565 13495 24599
rect 14289 24565 14323 24599
rect 18797 24565 18831 24599
rect 19533 24565 19567 24599
rect 20085 24565 20119 24599
rect 20821 24565 20855 24599
rect 23949 24565 23983 24599
rect 25973 24565 26007 24599
rect 27353 24565 27387 24599
rect 27997 24565 28031 24599
rect 12173 24361 12207 24395
rect 13645 24361 13679 24395
rect 20177 24361 20211 24395
rect 23581 24361 23615 24395
rect 24961 24361 24995 24395
rect 27261 24361 27295 24395
rect 27905 24361 27939 24395
rect 15393 24293 15427 24327
rect 16865 24293 16899 24327
rect 21465 24293 21499 24327
rect 22937 24293 22971 24327
rect 8493 24225 8527 24259
rect 9413 24225 9447 24259
rect 10977 24225 11011 24259
rect 11621 24225 11655 24259
rect 17417 24225 17451 24259
rect 22569 24225 22603 24259
rect 24593 24225 24627 24259
rect 26065 24225 26099 24259
rect 8401 24157 8435 24191
rect 9229 24157 9263 24191
rect 12357 24157 12391 24191
rect 12817 24157 12851 24191
rect 13553 24157 13587 24191
rect 14933 24157 14967 24191
rect 15577 24157 15611 24191
rect 16129 24157 16163 24191
rect 16773 24157 16807 24191
rect 17601 24157 17635 24191
rect 18613 24157 18647 24191
rect 19441 24157 19475 24191
rect 20361 24157 20395 24191
rect 20821 24157 20855 24191
rect 21649 24157 21683 24191
rect 22385 24157 22419 24191
rect 23489 24157 23523 24191
rect 24777 24157 24811 24191
rect 26249 24157 26283 24191
rect 27169 24157 27203 24191
rect 27813 24157 27847 24191
rect 11069 24089 11103 24123
rect 18061 24089 18095 24123
rect 19533 24089 19567 24123
rect 26709 24089 26743 24123
rect 9873 24021 9907 24055
rect 12909 24021 12943 24055
rect 14749 24021 14783 24055
rect 16221 24021 16255 24055
rect 18705 24021 18739 24055
rect 20913 24021 20947 24055
rect 8033 23817 8067 23851
rect 9505 23817 9539 23851
rect 25145 23817 25179 23851
rect 25697 23817 25731 23851
rect 14749 23749 14783 23783
rect 15301 23749 15335 23783
rect 18521 23749 18555 23783
rect 19165 23749 19199 23783
rect 23305 23749 23339 23783
rect 23397 23749 23431 23783
rect 1777 23681 1811 23715
rect 8217 23681 8251 23715
rect 8861 23681 8895 23715
rect 9321 23681 9355 23715
rect 10333 23681 10367 23715
rect 11161 23681 11195 23715
rect 12173 23681 12207 23715
rect 12633 23681 12667 23715
rect 13645 23681 13679 23715
rect 15853 23681 15887 23715
rect 17049 23681 17083 23715
rect 18061 23681 18095 23715
rect 20177 23681 20211 23715
rect 20821 23681 20855 23715
rect 22293 23681 22327 23715
rect 24409 23681 24443 23715
rect 25053 23681 25087 23715
rect 25881 23681 25915 23715
rect 26525 23681 26559 23715
rect 28365 23681 28399 23715
rect 13461 23613 13495 23647
rect 14657 23613 14691 23647
rect 16129 23613 16163 23647
rect 17877 23613 17911 23647
rect 19073 23613 19107 23647
rect 19533 23613 19567 23647
rect 20913 23613 20947 23647
rect 1593 23545 1627 23579
rect 10977 23545 11011 23579
rect 11989 23545 12023 23579
rect 20269 23545 20303 23579
rect 23857 23545 23891 23579
rect 8677 23477 8711 23511
rect 12725 23477 12759 23511
rect 14105 23477 14139 23511
rect 16865 23477 16899 23511
rect 22385 23477 22419 23511
rect 24501 23477 24535 23511
rect 26341 23477 26375 23511
rect 28181 23477 28215 23511
rect 10609 23273 10643 23307
rect 14933 23273 14967 23307
rect 18705 23273 18739 23307
rect 24685 23273 24719 23307
rect 26433 23273 26467 23307
rect 10425 23137 10459 23171
rect 11345 23137 11379 23171
rect 12449 23137 12483 23171
rect 12633 23137 12667 23171
rect 14473 23137 14507 23171
rect 22661 23137 22695 23171
rect 9597 23069 9631 23103
rect 10241 23069 10275 23103
rect 11529 23069 11563 23103
rect 13737 23069 13771 23103
rect 14289 23069 14323 23103
rect 15393 23069 15427 23103
rect 17509 23069 17543 23103
rect 18153 23069 18187 23103
rect 18613 23069 18647 23103
rect 20637 23069 20671 23103
rect 21281 23069 21315 23103
rect 21925 23069 21959 23103
rect 24593 23069 24627 23103
rect 25881 23069 25915 23103
rect 26341 23069 26375 23103
rect 27997 23069 28031 23103
rect 11989 23001 12023 23035
rect 13093 23001 13127 23035
rect 16221 23001 16255 23035
rect 16313 23001 16347 23035
rect 16865 23001 16899 23035
rect 19533 23001 19567 23035
rect 19625 23001 19659 23035
rect 20177 23001 20211 23035
rect 20729 23001 20763 23035
rect 22753 23001 22787 23035
rect 23673 23001 23707 23035
rect 9689 22933 9723 22967
rect 13553 22933 13587 22967
rect 15485 22933 15519 22967
rect 17325 22933 17359 22967
rect 17969 22933 18003 22967
rect 21373 22933 21407 22967
rect 22017 22933 22051 22967
rect 25697 22933 25731 22967
rect 28089 22933 28123 22967
rect 11897 22729 11931 22763
rect 19349 22729 19383 22763
rect 13369 22661 13403 22695
rect 15761 22661 15795 22695
rect 16313 22661 16347 22695
rect 24317 22661 24351 22695
rect 8401 22593 8435 22627
rect 9045 22593 9079 22627
rect 9689 22593 9723 22627
rect 10333 22593 10367 22627
rect 11161 22593 11195 22627
rect 11805 22593 11839 22627
rect 13093 22593 13127 22627
rect 14197 22593 14231 22627
rect 15025 22593 15059 22627
rect 17049 22593 17083 22627
rect 17509 22593 17543 22627
rect 19993 22593 20027 22627
rect 20913 22593 20947 22627
rect 22017 22593 22051 22627
rect 22937 22593 22971 22627
rect 23121 22593 23155 22627
rect 24041 22593 24075 22627
rect 28089 22593 28123 22627
rect 12449 22525 12483 22559
rect 15669 22525 15703 22559
rect 18705 22525 18739 22559
rect 18889 22525 18923 22559
rect 19809 22525 19843 22559
rect 9505 22457 9539 22491
rect 10425 22457 10459 22491
rect 17601 22457 17635 22491
rect 28273 22457 28307 22491
rect 8217 22389 8251 22423
rect 8861 22389 8895 22423
rect 10977 22389 11011 22423
rect 14289 22389 14323 22423
rect 14841 22389 14875 22423
rect 16865 22389 16899 22423
rect 20177 22389 20211 22423
rect 21005 22389 21039 22423
rect 22109 22389 22143 22423
rect 23305 22389 23339 22423
rect 25789 22389 25823 22423
rect 19441 22185 19475 22219
rect 17049 22117 17083 22151
rect 11069 22049 11103 22083
rect 13277 22049 13311 22083
rect 15301 22049 15335 22083
rect 15945 22049 15979 22083
rect 16589 22049 16623 22083
rect 18245 22049 18279 22083
rect 21005 22049 21039 22083
rect 22937 22049 22971 22083
rect 1777 21981 1811 22015
rect 9505 21981 9539 22015
rect 10425 21981 10459 22015
rect 10885 21981 10919 22015
rect 11989 21981 12023 22015
rect 12173 21981 12207 22015
rect 13093 21981 13127 22015
rect 14757 21981 14791 22015
rect 16405 21981 16439 22015
rect 18705 21981 18739 22015
rect 19625 21981 19659 22015
rect 22845 21981 22879 22015
rect 23489 21981 23523 22015
rect 24777 21981 24811 22015
rect 25237 21981 25271 22015
rect 26249 21981 26283 22015
rect 15393 21913 15427 21947
rect 17601 21913 17635 21947
rect 17693 21913 17727 21947
rect 20545 21913 20579 21947
rect 20637 21913 20671 21947
rect 21741 21913 21775 21947
rect 21833 21913 21867 21947
rect 22385 21913 22419 21947
rect 25329 21913 25363 21947
rect 26525 21913 26559 21947
rect 1593 21845 1627 21879
rect 9321 21845 9355 21879
rect 10241 21845 10275 21879
rect 11529 21845 11563 21879
rect 12633 21845 12667 21879
rect 13737 21845 13771 21879
rect 14565 21845 14599 21879
rect 18797 21845 18831 21879
rect 23581 21845 23615 21879
rect 24593 21845 24627 21879
rect 27997 21845 28031 21879
rect 7389 21641 7423 21675
rect 20821 21641 20855 21675
rect 26525 21641 26559 21675
rect 15761 21573 15795 21607
rect 23029 21573 23063 21607
rect 7297 21505 7331 21539
rect 9597 21505 9631 21539
rect 10517 21505 10551 21539
rect 10977 21505 11011 21539
rect 11805 21505 11839 21539
rect 11897 21505 11931 21539
rect 13829 21505 13863 21539
rect 14657 21505 14691 21539
rect 16865 21505 16899 21539
rect 20177 21505 20211 21539
rect 22017 21505 22051 21539
rect 22753 21505 22787 21539
rect 26433 21505 26467 21539
rect 27169 21505 27203 21539
rect 28089 21505 28123 21539
rect 12449 21437 12483 21471
rect 12633 21437 12667 21471
rect 15117 21437 15151 21471
rect 15301 21437 15335 21471
rect 17969 21437 18003 21471
rect 18245 21437 18279 21471
rect 24501 21437 24535 21471
rect 9413 21369 9447 21403
rect 11069 21369 11103 21403
rect 13921 21369 13955 21403
rect 10333 21301 10367 21335
rect 12817 21301 12851 21335
rect 14473 21301 14507 21335
rect 16957 21301 16991 21335
rect 19717 21301 19751 21335
rect 20269 21301 20303 21335
rect 22109 21301 22143 21335
rect 27261 21301 27295 21335
rect 28273 21301 28307 21335
rect 11161 21097 11195 21131
rect 15117 21097 15151 21131
rect 15945 21097 15979 21131
rect 17785 21097 17819 21131
rect 20526 21097 20560 21131
rect 23121 21097 23155 21131
rect 13461 21029 13495 21063
rect 17233 21029 17267 21063
rect 22017 21029 22051 21063
rect 23673 21029 23707 21063
rect 13277 20961 13311 20995
rect 14565 20961 14599 20995
rect 14749 20961 14783 20995
rect 20269 20961 20303 20995
rect 22477 20961 22511 20995
rect 22661 20961 22695 20995
rect 26341 20961 26375 20995
rect 1777 20893 1811 20927
rect 6101 20893 6135 20927
rect 10241 20893 10275 20927
rect 11069 20893 11103 20927
rect 11989 20893 12023 20927
rect 12173 20893 12207 20927
rect 13093 20893 13127 20927
rect 16129 20893 16163 20927
rect 17969 20893 18003 20927
rect 18429 20893 18463 20927
rect 19441 20893 19475 20927
rect 23581 20893 23615 20927
rect 16681 20825 16715 20859
rect 16773 20825 16807 20859
rect 26617 20825 26651 20859
rect 28365 20825 28399 20859
rect 1593 20757 1627 20791
rect 6193 20757 6227 20791
rect 9597 20757 9631 20791
rect 10333 20757 10367 20791
rect 12633 20757 12667 20791
rect 18521 20757 18555 20791
rect 19533 20757 19567 20791
rect 10517 20553 10551 20587
rect 22017 20553 22051 20587
rect 27905 20553 27939 20587
rect 18337 20485 18371 20519
rect 8769 20417 8803 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 11161 20417 11195 20451
rect 11713 20417 11747 20451
rect 12817 20417 12851 20451
rect 14565 20417 14599 20451
rect 16037 20417 16071 20451
rect 16865 20417 16899 20451
rect 18061 20417 18095 20451
rect 20913 20417 20947 20451
rect 28089 20417 28123 20451
rect 4629 20349 4663 20383
rect 4813 20349 4847 20383
rect 11897 20349 11931 20383
rect 13461 20349 13495 20383
rect 13645 20349 13679 20383
rect 14749 20349 14783 20383
rect 20269 20349 20303 20383
rect 20453 20349 20487 20383
rect 23213 20349 23247 20383
rect 23489 20349 23523 20383
rect 25237 20349 25271 20383
rect 14105 20281 14139 20315
rect 5273 20213 5307 20247
rect 8861 20213 8895 20247
rect 10977 20213 11011 20247
rect 12357 20213 12391 20247
rect 14933 20213 14967 20247
rect 15853 20213 15887 20247
rect 16957 20213 16991 20247
rect 19809 20213 19843 20247
rect 5089 20009 5123 20043
rect 6193 20009 6227 20043
rect 11069 20009 11103 20043
rect 12909 20009 12943 20043
rect 28181 20009 28215 20043
rect 21281 19941 21315 19975
rect 15301 19873 15335 19907
rect 19533 19873 19567 19907
rect 21741 19873 21775 19907
rect 22017 19873 22051 19907
rect 24685 19873 24719 19907
rect 1777 19805 1811 19839
rect 5089 19805 5123 19839
rect 6101 19805 6135 19839
rect 9137 19805 9171 19839
rect 10517 19805 10551 19839
rect 10977 19805 11011 19839
rect 11621 19805 11655 19839
rect 13093 19805 13127 19839
rect 13737 19805 13771 19839
rect 14841 19805 14875 19839
rect 15485 19805 15519 19839
rect 17785 19805 17819 19839
rect 17877 19805 17911 19839
rect 18421 19815 18455 19849
rect 28365 19805 28399 19839
rect 15945 19737 15979 19771
rect 16681 19737 16715 19771
rect 16773 19737 16807 19771
rect 17325 19737 17359 19771
rect 19809 19737 19843 19771
rect 24961 19737 24995 19771
rect 26709 19737 26743 19771
rect 1593 19669 1627 19703
rect 9229 19669 9263 19703
rect 10333 19669 10367 19703
rect 11713 19669 11747 19703
rect 12265 19669 12299 19703
rect 13553 19669 13587 19703
rect 14657 19669 14691 19703
rect 18521 19669 18555 19703
rect 23489 19669 23523 19703
rect 6561 19465 6595 19499
rect 10333 19465 10367 19499
rect 10977 19465 11011 19499
rect 11989 19465 12023 19499
rect 13277 19465 13311 19499
rect 14381 19465 14415 19499
rect 14841 19465 14875 19499
rect 16037 19465 16071 19499
rect 17601 19465 17635 19499
rect 24133 19465 24167 19499
rect 26525 19465 26559 19499
rect 22661 19397 22695 19431
rect 6745 19329 6779 19363
rect 7573 19329 7607 19363
rect 9873 19329 9907 19363
rect 10517 19329 10551 19363
rect 11161 19329 11195 19363
rect 12173 19329 12207 19363
rect 12633 19329 12667 19363
rect 15025 19329 15059 19363
rect 15945 19329 15979 19363
rect 17509 19329 17543 19363
rect 18153 19329 18187 19363
rect 20361 19329 20395 19363
rect 22385 19329 22419 19363
rect 24777 19329 24811 19363
rect 12817 19261 12851 19295
rect 13737 19261 13771 19295
rect 13921 19261 13955 19295
rect 16865 19261 16899 19295
rect 18429 19261 18463 19295
rect 25053 19261 25087 19295
rect 7389 19125 7423 19159
rect 9689 19125 9723 19159
rect 19901 19125 19935 19159
rect 20453 19125 20487 19159
rect 9965 18921 9999 18955
rect 17785 18921 17819 18955
rect 22845 18921 22879 18955
rect 28181 18921 28215 18955
rect 7113 18785 7147 18819
rect 8493 18785 8527 18819
rect 9505 18785 9539 18819
rect 11621 18785 11655 18819
rect 12265 18785 12299 18819
rect 14841 18785 14875 18819
rect 15945 18785 15979 18819
rect 21097 18785 21131 18819
rect 24593 18785 24627 18819
rect 26617 18785 26651 18819
rect 1593 18717 1627 18751
rect 6929 18717 6963 18751
rect 8401 18717 8435 18751
rect 9321 18717 9355 18751
rect 11805 18717 11839 18751
rect 13185 18717 13219 18751
rect 15485 18717 15519 18751
rect 16129 18717 16163 18751
rect 17049 18717 17083 18751
rect 17693 18717 17727 18751
rect 18329 18719 18363 18753
rect 28365 18717 28399 18751
rect 14933 18649 14967 18683
rect 21373 18649 21407 18683
rect 24869 18649 24903 18683
rect 1777 18581 1811 18615
rect 7573 18581 7607 18615
rect 10977 18581 11011 18615
rect 13277 18581 13311 18615
rect 16589 18581 16623 18615
rect 17141 18581 17175 18615
rect 18429 18581 18463 18615
rect 8309 18377 8343 18411
rect 13737 18377 13771 18411
rect 15485 18377 15519 18411
rect 19993 18377 20027 18411
rect 14473 18309 14507 18343
rect 16957 18309 16991 18343
rect 17049 18309 17083 18343
rect 25605 18309 25639 18343
rect 4445 18241 4479 18275
rect 5273 18241 5307 18275
rect 7849 18241 7883 18275
rect 9229 18241 9263 18275
rect 9873 18241 9907 18275
rect 10517 18241 10551 18275
rect 11161 18241 11195 18275
rect 12265 18241 12299 18275
rect 13645 18241 13679 18275
rect 15025 18241 15059 18275
rect 15669 18241 15703 18275
rect 16129 18241 16163 18275
rect 16221 18241 16255 18275
rect 7665 18173 7699 18207
rect 12449 18173 12483 18207
rect 14381 18173 14415 18207
rect 17233 18173 17267 18207
rect 18245 18173 18279 18207
rect 18521 18173 18555 18207
rect 23581 18173 23615 18207
rect 23857 18173 23891 18207
rect 4261 18105 4295 18139
rect 9045 18105 9079 18139
rect 10333 18105 10367 18139
rect 5089 18037 5123 18071
rect 9689 18037 9723 18071
rect 10977 18037 11011 18071
rect 12817 18037 12851 18071
rect 7757 17833 7791 17867
rect 8401 17833 8435 17867
rect 9321 17833 9355 17867
rect 11805 17833 11839 17867
rect 27077 17833 27111 17867
rect 15209 17765 15243 17799
rect 15945 17765 15979 17799
rect 25053 17765 25087 17799
rect 10057 17697 10091 17731
rect 19441 17697 19475 17731
rect 21649 17697 21683 17731
rect 25329 17697 25363 17731
rect 25605 17697 25639 17731
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9229 17629 9263 17663
rect 9873 17629 9907 17663
rect 11345 17629 11379 17663
rect 11989 17629 12023 17663
rect 12633 17629 12667 17663
rect 13093 17629 13127 17663
rect 13277 17629 13311 17663
rect 13737 17629 13771 17663
rect 14841 17629 14875 17663
rect 15025 17629 15059 17663
rect 16129 17629 16163 17663
rect 16589 17629 16623 17663
rect 17509 17629 17543 17663
rect 18153 17629 18187 17663
rect 10517 17561 10551 17595
rect 16865 17561 16899 17595
rect 19717 17561 19751 17595
rect 21925 17561 21959 17595
rect 5825 17493 5859 17527
rect 11161 17493 11195 17527
rect 12449 17493 12483 17527
rect 17601 17493 17635 17527
rect 18245 17493 18279 17527
rect 21189 17493 21223 17527
rect 23397 17493 23431 17527
rect 6653 17289 6687 17323
rect 10977 17289 11011 17323
rect 12357 17289 12391 17323
rect 26525 17289 26559 17323
rect 7481 17221 7515 17255
rect 8585 17221 8619 17255
rect 8677 17221 8711 17255
rect 13093 17221 13127 17255
rect 13194 17221 13228 17255
rect 14933 17221 14967 17255
rect 15485 17221 15519 17255
rect 1593 17153 1627 17187
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 6837 17153 6871 17187
rect 10333 17153 10367 17187
rect 11161 17153 11195 17187
rect 11897 17153 11931 17187
rect 12541 17153 12575 17187
rect 16129 17153 16163 17187
rect 16865 17153 16899 17187
rect 18061 17153 18095 17187
rect 20269 17153 20303 17187
rect 22569 17153 22603 17187
rect 24777 17153 24811 17187
rect 28365 17153 28399 17187
rect 7389 17085 7423 17119
rect 7665 17085 7699 17119
rect 13369 17085 13403 17119
rect 14841 17085 14875 17119
rect 17141 17085 17175 17119
rect 18337 17085 18371 17119
rect 22845 17085 22879 17119
rect 24317 17085 24351 17119
rect 25053 17085 25087 17119
rect 1777 17017 1811 17051
rect 5733 17017 5767 17051
rect 9137 17017 9171 17051
rect 10149 17017 10183 17051
rect 11713 17017 11747 17051
rect 16221 16949 16255 16983
rect 19809 16949 19843 16983
rect 20361 16949 20395 16983
rect 28181 16949 28215 16983
rect 5457 16745 5491 16779
rect 7757 16745 7791 16779
rect 9689 16609 9723 16643
rect 9873 16609 9907 16643
rect 12633 16609 12667 16643
rect 12909 16609 12943 16643
rect 14289 16609 14323 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 19441 16609 19475 16643
rect 19717 16609 19751 16643
rect 21649 16609 21683 16643
rect 26341 16609 26375 16643
rect 26617 16609 26651 16643
rect 5641 16541 5675 16575
rect 6285 16541 6319 16575
rect 7021 16541 7055 16575
rect 7113 16541 7147 16575
rect 7941 16541 7975 16575
rect 8401 16541 8435 16575
rect 11529 16541 11563 16575
rect 15117 16541 15151 16575
rect 17049 16541 17083 16575
rect 17693 16541 17727 16575
rect 18337 16541 18371 16575
rect 8493 16473 8527 16507
rect 12725 16473 12759 16507
rect 21925 16473 21959 16507
rect 28365 16473 28399 16507
rect 6377 16405 6411 16439
rect 10333 16405 10367 16439
rect 11345 16405 11379 16439
rect 14933 16405 14967 16439
rect 16221 16405 16255 16439
rect 17141 16405 17175 16439
rect 17785 16405 17819 16439
rect 18429 16405 18463 16439
rect 21189 16405 21223 16439
rect 23397 16405 23431 16439
rect 12357 16201 12391 16235
rect 14197 16201 14231 16235
rect 14841 16201 14875 16235
rect 15485 16201 15519 16235
rect 9137 16133 9171 16167
rect 17509 16133 17543 16167
rect 24685 16133 24719 16167
rect 1777 16065 1811 16099
rect 4905 16065 4939 16099
rect 8401 16065 8435 16099
rect 9045 16065 9079 16099
rect 9873 16065 9907 16099
rect 12265 16065 12299 16099
rect 13093 16065 13127 16099
rect 13737 16065 13771 16099
rect 14381 16065 14415 16099
rect 15669 16065 15703 16099
rect 18153 16065 18187 16099
rect 18705 16065 18739 16099
rect 21281 16065 21315 16099
rect 22201 16065 22235 16099
rect 24409 16065 24443 16099
rect 28089 16065 28123 16099
rect 10333 15997 10367 16031
rect 10517 15997 10551 16031
rect 16129 15997 16163 16031
rect 16865 15997 16899 16031
rect 17049 15997 17083 16031
rect 18981 15997 19015 16031
rect 22477 15997 22511 16031
rect 26433 15997 26467 16031
rect 1593 15929 1627 15963
rect 8493 15929 8527 15963
rect 12909 15929 12943 15963
rect 4997 15861 5031 15895
rect 9689 15861 9723 15895
rect 10977 15861 11011 15895
rect 13553 15861 13587 15895
rect 17969 15861 18003 15895
rect 20453 15861 20487 15895
rect 21373 15861 21407 15895
rect 23949 15861 23983 15895
rect 28273 15861 28307 15895
rect 6929 15657 6963 15691
rect 11069 15657 11103 15691
rect 9873 15589 9907 15623
rect 17233 15589 17267 15623
rect 23397 15589 23431 15623
rect 6285 15521 6319 15555
rect 7941 15521 7975 15555
rect 9229 15521 9263 15555
rect 11621 15521 11655 15555
rect 17049 15521 17083 15555
rect 19441 15521 19475 15555
rect 21649 15521 21683 15555
rect 26249 15521 26283 15555
rect 26525 15521 26559 15555
rect 6469 15453 6503 15487
rect 9137 15453 9171 15487
rect 9781 15453 9815 15487
rect 10425 15453 10459 15487
rect 10609 15453 10643 15487
rect 12909 15453 12943 15487
rect 13093 15453 13127 15487
rect 15945 15453 15979 15487
rect 16865 15453 16899 15487
rect 17969 15453 18003 15487
rect 18613 15453 18647 15487
rect 8033 15385 8067 15419
rect 8585 15385 8619 15419
rect 11713 15385 11747 15419
rect 12265 15385 12299 15419
rect 14657 15385 14691 15419
rect 14749 15385 14783 15419
rect 15301 15385 15335 15419
rect 16221 15385 16255 15419
rect 19717 15385 19751 15419
rect 21925 15385 21959 15419
rect 24685 15385 24719 15419
rect 24777 15385 24811 15419
rect 25329 15385 25363 15419
rect 28273 15385 28307 15419
rect 13553 15317 13587 15351
rect 18061 15317 18095 15351
rect 18705 15317 18739 15351
rect 21189 15317 21223 15351
rect 9045 15113 9079 15147
rect 10885 15113 10919 15147
rect 15761 15113 15795 15147
rect 19993 15113 20027 15147
rect 20545 15113 20579 15147
rect 21373 15113 21407 15147
rect 24133 15113 24167 15147
rect 14473 15045 14507 15079
rect 8953 14977 8987 15011
rect 9781 14977 9815 15011
rect 10425 14977 10459 15011
rect 11069 14977 11103 15011
rect 12173 14977 12207 15011
rect 13185 14977 13219 15011
rect 13369 14977 13403 15011
rect 15945 14977 15979 15011
rect 18245 14977 18279 15011
rect 20453 14977 20487 15011
rect 21281 14977 21315 15011
rect 22385 14977 22419 15011
rect 27169 14977 27203 15011
rect 27997 14977 28031 15011
rect 12357 14909 12391 14943
rect 14381 14909 14415 14943
rect 14657 14909 14691 14943
rect 17049 14909 17083 14943
rect 17233 14909 17267 14943
rect 18521 14909 18555 14943
rect 22661 14909 22695 14943
rect 24593 14909 24627 14943
rect 24869 14909 24903 14943
rect 26617 14909 26651 14943
rect 10241 14841 10275 14875
rect 9597 14773 9631 14807
rect 13829 14773 13863 14807
rect 17417 14773 17451 14807
rect 27261 14773 27295 14807
rect 28089 14773 28123 14807
rect 9689 14569 9723 14603
rect 12633 14569 12667 14603
rect 13553 14569 13587 14603
rect 15945 14569 15979 14603
rect 23581 14569 23615 14603
rect 28181 14569 28215 14603
rect 10977 14501 11011 14535
rect 14657 14501 14691 14535
rect 18613 14501 18647 14535
rect 22937 14501 22971 14535
rect 12449 14433 12483 14467
rect 15485 14433 15519 14467
rect 17141 14433 17175 14467
rect 17877 14433 17911 14467
rect 21189 14433 21223 14467
rect 26617 14433 26651 14467
rect 1777 14365 1811 14399
rect 4905 14365 4939 14399
rect 9597 14365 9631 14399
rect 10425 14365 10459 14399
rect 11161 14365 11195 14399
rect 11621 14365 11655 14399
rect 12265 14365 12299 14399
rect 13737 14365 13771 14399
rect 14841 14365 14875 14399
rect 15301 14365 15335 14399
rect 17601 14365 17635 14399
rect 18521 14365 18555 14399
rect 19441 14365 19475 14399
rect 20085 14365 20119 14399
rect 23489 14365 23523 14399
rect 24593 14365 24627 14399
rect 28365 14365 28399 14399
rect 16497 14297 16531 14331
rect 16589 14297 16623 14331
rect 19533 14297 19567 14331
rect 21465 14297 21499 14331
rect 24869 14297 24903 14331
rect 1593 14229 1627 14263
rect 4721 14229 4755 14263
rect 10241 14229 10275 14263
rect 11713 14229 11747 14263
rect 20177 14229 20211 14263
rect 1593 14025 1627 14059
rect 5825 14025 5859 14059
rect 10149 14025 10183 14059
rect 13553 14025 13587 14059
rect 14289 14025 14323 14059
rect 15945 14025 15979 14059
rect 19901 14025 19935 14059
rect 21281 14025 21315 14059
rect 23765 14025 23799 14059
rect 8861 13957 8895 13991
rect 10977 13957 11011 13991
rect 11897 13957 11931 13991
rect 17049 13957 17083 13991
rect 17601 13957 17635 13991
rect 24869 13957 24903 13991
rect 26617 13957 26651 13991
rect 1777 13889 1811 13923
rect 4905 13889 4939 13923
rect 6009 13889 6043 13923
rect 6561 13889 6595 13923
rect 8769 13889 8803 13923
rect 9597 13889 9631 13923
rect 10333 13889 10367 13923
rect 12449 13889 12483 13923
rect 13461 13889 13495 13923
rect 14197 13889 14231 13923
rect 15025 13889 15059 13923
rect 18153 13889 18187 13923
rect 20361 13889 20395 13923
rect 21189 13889 21223 13923
rect 4721 13821 4755 13855
rect 5365 13821 5399 13855
rect 6745 13821 6779 13855
rect 11805 13821 11839 13855
rect 14841 13821 14875 13855
rect 15485 13821 15519 13855
rect 16957 13821 16991 13855
rect 20453 13821 20487 13855
rect 22017 13821 22051 13855
rect 24593 13821 24627 13855
rect 7205 13685 7239 13719
rect 9413 13685 9447 13719
rect 18410 13685 18444 13719
rect 22274 13685 22308 13719
rect 3341 13481 3375 13515
rect 8309 13481 8343 13515
rect 13737 13481 13771 13515
rect 14657 13481 14691 13515
rect 15853 13481 15887 13515
rect 24685 13481 24719 13515
rect 25789 13481 25823 13515
rect 7021 13413 7055 13447
rect 11897 13413 11931 13447
rect 18153 13413 18187 13447
rect 21189 13413 21223 13447
rect 7941 13345 7975 13379
rect 10333 13345 10367 13379
rect 11713 13345 11747 13379
rect 13093 13345 13127 13379
rect 15209 13345 15243 13379
rect 17785 13345 17819 13379
rect 19441 13345 19475 13379
rect 21741 13345 21775 13379
rect 23489 13345 23523 13379
rect 26341 13345 26375 13379
rect 26617 13345 26651 13379
rect 28365 13345 28399 13379
rect 3249 13277 3283 13311
rect 4169 13277 4203 13311
rect 4353 13277 4387 13311
rect 5273 13277 5307 13311
rect 6653 13277 6687 13311
rect 6837 13277 6871 13311
rect 7757 13277 7791 13311
rect 10241 13277 10275 13311
rect 11069 13277 11103 13311
rect 11529 13277 11563 13311
rect 13277 13277 13311 13311
rect 14565 13277 14599 13311
rect 15393 13277 15427 13311
rect 17325 13277 17359 13311
rect 17969 13277 18003 13311
rect 24593 13277 24627 13311
rect 25697 13277 25731 13311
rect 16681 13209 16715 13243
rect 16773 13209 16807 13243
rect 19717 13209 19751 13243
rect 22017 13209 22051 13243
rect 4813 13141 4847 13175
rect 5365 13141 5399 13175
rect 9597 13141 9631 13175
rect 10885 13141 10919 13175
rect 4261 12937 4295 12971
rect 5733 12937 5767 12971
rect 11989 12937 12023 12971
rect 15025 12937 15059 12971
rect 17693 12937 17727 12971
rect 24317 12937 24351 12971
rect 26525 12937 26559 12971
rect 8861 12869 8895 12903
rect 10517 12869 10551 12903
rect 10609 12869 10643 12903
rect 11161 12869 11195 12903
rect 12817 12869 12851 12903
rect 15761 12869 15795 12903
rect 19717 12869 19751 12903
rect 22845 12869 22879 12903
rect 1777 12801 1811 12835
rect 5917 12801 5951 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 12173 12801 12207 12835
rect 14013 12801 14047 12835
rect 14933 12801 14967 12835
rect 16865 12801 16899 12835
rect 17601 12801 17635 12835
rect 18429 12801 18463 12835
rect 19441 12801 19475 12835
rect 24777 12801 24811 12835
rect 28365 12801 28399 12835
rect 8033 12733 8067 12767
rect 8769 12733 8803 12767
rect 9045 12733 9079 12767
rect 12725 12733 12759 12767
rect 13001 12733 13035 12767
rect 15669 12733 15703 12767
rect 16313 12733 16347 12767
rect 18245 12733 18279 12767
rect 18889 12733 18923 12767
rect 21465 12733 21499 12767
rect 22569 12733 22603 12767
rect 6929 12665 6963 12699
rect 13829 12665 13863 12699
rect 1593 12597 1627 12631
rect 16957 12597 16991 12631
rect 25040 12597 25074 12631
rect 28181 12597 28215 12631
rect 6745 12393 6779 12427
rect 7665 12393 7699 12427
rect 9229 12393 9263 12427
rect 9873 12393 9907 12427
rect 11805 12393 11839 12427
rect 15853 12393 15887 12427
rect 18153 12393 18187 12427
rect 25329 12393 25363 12427
rect 11253 12325 11287 12359
rect 24041 12325 24075 12359
rect 13093 12257 13127 12291
rect 14565 12257 14599 12291
rect 16865 12257 16899 12291
rect 19717 12257 19751 12291
rect 24685 12257 24719 12291
rect 27997 12257 28031 12291
rect 4905 12189 4939 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 6653 12189 6687 12223
rect 7565 12189 7599 12223
rect 8585 12189 8619 12223
rect 9413 12189 9447 12223
rect 10057 12189 10091 12223
rect 11161 12189 11195 12223
rect 11989 12189 12023 12223
rect 12449 12189 12483 12223
rect 13277 12189 13311 12223
rect 16037 12189 16071 12223
rect 18061 12189 18095 12223
rect 18705 12189 18739 12223
rect 22293 12189 22327 12223
rect 24593 12189 24627 12223
rect 25237 12189 25271 12223
rect 26249 12189 26283 12223
rect 12541 12121 12575 12155
rect 14657 12121 14691 12155
rect 15209 12121 15243 12155
rect 16589 12121 16623 12155
rect 16681 12121 16715 12155
rect 19993 12121 20027 12155
rect 21741 12121 21775 12155
rect 22569 12121 22603 12155
rect 26525 12121 26559 12155
rect 6193 12053 6227 12087
rect 8401 12053 8435 12087
rect 10517 12053 10551 12087
rect 13737 12053 13771 12087
rect 18797 12053 18831 12087
rect 5733 11849 5767 11883
rect 9413 11849 9447 11883
rect 13461 11849 13495 11883
rect 15393 11849 15427 11883
rect 16129 11849 16163 11883
rect 23765 11849 23799 11883
rect 10517 11781 10551 11815
rect 10609 11781 10643 11815
rect 14013 11781 14047 11815
rect 14105 11781 14139 11815
rect 16957 11781 16991 11815
rect 22293 11781 22327 11815
rect 5917 11713 5951 11747
rect 7205 11713 7239 11747
rect 7665 11713 7699 11747
rect 9597 11713 9631 11747
rect 11713 11713 11747 11747
rect 15301 11713 15335 11747
rect 16313 11713 16347 11747
rect 16865 11713 16899 11747
rect 17693 11713 17727 11747
rect 22017 11713 22051 11747
rect 24593 11713 24627 11747
rect 8309 11645 8343 11679
rect 8493 11645 8527 11679
rect 11897 11645 11931 11679
rect 12817 11645 12851 11679
rect 13001 11645 13035 11679
rect 14289 11645 14323 11679
rect 18429 11645 18463 11679
rect 18705 11645 18739 11679
rect 20177 11645 20211 11679
rect 24869 11645 24903 11679
rect 26617 11645 26651 11679
rect 11069 11577 11103 11611
rect 7021 11509 7055 11543
rect 7757 11509 7791 11543
rect 8953 11509 8987 11543
rect 12357 11509 12391 11543
rect 17509 11509 17543 11543
rect 1593 11305 1627 11339
rect 7021 11305 7055 11339
rect 7665 11305 7699 11339
rect 10609 11305 10643 11339
rect 12541 11305 12575 11339
rect 14657 11305 14691 11339
rect 15393 11305 15427 11339
rect 23673 11305 23707 11339
rect 25053 11305 25087 11339
rect 17601 11237 17635 11271
rect 20085 11237 20119 11271
rect 8493 11169 8527 11203
rect 9229 11169 9263 11203
rect 9689 11169 9723 11203
rect 11345 11169 11379 11203
rect 14473 11169 14507 11203
rect 17141 11169 17175 11203
rect 18337 11169 18371 11203
rect 21373 11169 21407 11203
rect 23121 11169 23155 11203
rect 26341 11169 26375 11203
rect 26617 11169 26651 11203
rect 28365 11169 28399 11203
rect 1777 11101 1811 11135
rect 7205 11101 7239 11135
rect 7849 11101 7883 11135
rect 8401 11101 8435 11135
rect 10793 11101 10827 11135
rect 12449 11101 12483 11135
rect 13553 11101 13587 11135
rect 14289 11101 14323 11135
rect 15577 11101 15611 11135
rect 17785 11101 17819 11135
rect 18245 11101 18279 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 20269 11101 20303 11135
rect 23581 11101 23615 11135
rect 24961 11101 24995 11135
rect 25605 11101 25639 11135
rect 9321 11033 9355 11067
rect 11437 11033 11471 11067
rect 11989 11033 12023 11067
rect 16129 11033 16163 11067
rect 16221 11033 16255 11067
rect 21649 11033 21683 11067
rect 13645 10965 13679 10999
rect 25697 10965 25731 10999
rect 6745 10761 6779 10795
rect 8309 10761 8343 10795
rect 9505 10761 9539 10795
rect 10977 10761 11011 10795
rect 12817 10761 12851 10795
rect 16865 10761 16899 10795
rect 17509 10761 17543 10795
rect 21373 10761 21407 10795
rect 28273 10761 28307 10795
rect 13737 10693 13771 10727
rect 14841 10693 14875 10727
rect 15577 10693 15611 10727
rect 20269 10693 20303 10727
rect 22385 10693 22419 10727
rect 6929 10625 6963 10659
rect 9689 10625 9723 10659
rect 11161 10625 11195 10659
rect 12357 10625 12391 10659
rect 13001 10625 13035 10659
rect 14749 10625 14783 10659
rect 17049 10609 17083 10643
rect 17693 10629 17727 10663
rect 21289 10623 21323 10657
rect 22109 10625 22143 10659
rect 24777 10625 24811 10659
rect 28089 10625 28123 10659
rect 13645 10557 13679 10591
rect 15485 10557 15519 10591
rect 18245 10557 18279 10591
rect 18521 10557 18555 10591
rect 24133 10557 24167 10591
rect 24501 10557 24535 10591
rect 25053 10557 25087 10591
rect 12173 10489 12207 10523
rect 14197 10489 14231 10523
rect 16037 10489 16071 10523
rect 26525 10421 26559 10455
rect 24041 10217 24075 10251
rect 26893 10217 26927 10251
rect 10609 10149 10643 10183
rect 17141 10149 17175 10183
rect 28181 10149 28215 10183
rect 12725 10081 12759 10115
rect 13185 10081 13219 10115
rect 16589 10081 16623 10115
rect 17785 10081 17819 10115
rect 19809 10081 19843 10115
rect 25145 10081 25179 10115
rect 1593 10013 1627 10047
rect 4813 10013 4847 10047
rect 9689 10013 9723 10047
rect 10793 10013 10827 10047
rect 11253 10013 11287 10047
rect 11437 10013 11471 10047
rect 12541 10013 12575 10047
rect 22293 10013 22327 10047
rect 28365 10013 28399 10047
rect 14473 9945 14507 9979
rect 15209 9945 15243 9979
rect 15301 9945 15335 9979
rect 15853 9945 15887 9979
rect 16681 9945 16715 9979
rect 17877 9945 17911 9979
rect 18429 9945 18463 9979
rect 20085 9945 20119 9979
rect 21833 9945 21867 9979
rect 22569 9945 22603 9979
rect 25408 9945 25442 9979
rect 1777 9877 1811 9911
rect 4905 9877 4939 9911
rect 9505 9877 9539 9911
rect 11897 9877 11931 9911
rect 3617 9673 3651 9707
rect 10977 9673 11011 9707
rect 12173 9673 12207 9707
rect 14933 9673 14967 9707
rect 17509 9605 17543 9639
rect 18245 9605 18279 9639
rect 22845 9605 22879 9639
rect 3801 9537 3835 9571
rect 6653 9537 6687 9571
rect 8401 9537 8435 9571
rect 9229 9537 9263 9571
rect 9873 9537 9907 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 11161 9537 11195 9571
rect 12357 9537 12391 9571
rect 13001 9537 13035 9571
rect 13829 9537 13863 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15577 9537 15611 9571
rect 16865 9537 16899 9571
rect 17049 9537 17083 9571
rect 17969 9537 18003 9571
rect 22569 9537 22603 9571
rect 24869 9537 24903 9571
rect 28365 9537 28399 9571
rect 19717 9469 19751 9503
rect 25145 9469 25179 9503
rect 26617 9469 26651 9503
rect 9045 9401 9079 9435
rect 9689 9401 9723 9435
rect 13645 9401 13679 9435
rect 15669 9401 15703 9435
rect 28181 9401 28215 9435
rect 6745 9333 6779 9367
rect 8493 9333 8527 9367
rect 13093 9333 13127 9367
rect 14289 9333 14323 9367
rect 24317 9333 24351 9367
rect 8493 9129 8527 9163
rect 11345 9129 11379 9163
rect 12541 9129 12575 9163
rect 24685 9129 24719 9163
rect 14657 9061 14691 9095
rect 7849 8993 7883 9027
rect 9965 8993 9999 9027
rect 12081 8993 12115 9027
rect 14473 8993 14507 9027
rect 16037 8993 16071 9027
rect 17141 8993 17175 9027
rect 21005 8993 21039 9027
rect 22753 8993 22787 9027
rect 26065 8993 26099 9027
rect 26341 8993 26375 9027
rect 28089 8993 28123 9027
rect 1593 8925 1627 8959
rect 5917 8925 5951 8959
rect 7757 8925 7791 8959
rect 8401 8925 8435 8959
rect 9321 8925 9355 8959
rect 10149 8925 10183 8959
rect 11253 8925 11287 8959
rect 11897 8925 11931 8959
rect 13553 8925 13587 8959
rect 14289 8925 14323 8959
rect 23305 8925 23339 8959
rect 24593 8925 24627 8959
rect 25237 8925 25271 8959
rect 13645 8857 13679 8891
rect 16129 8857 16163 8891
rect 16681 8857 16715 8891
rect 17417 8857 17451 8891
rect 21281 8857 21315 8891
rect 23397 8857 23431 8891
rect 1685 8789 1719 8823
rect 5733 8789 5767 8823
rect 9413 8789 9447 8823
rect 10609 8789 10643 8823
rect 18889 8789 18923 8823
rect 25329 8789 25363 8823
rect 8217 8585 8251 8619
rect 9413 8585 9447 8619
rect 15945 8585 15979 8619
rect 16957 8585 16991 8619
rect 20085 8585 20119 8619
rect 28089 8585 28123 8619
rect 12449 8517 12483 8551
rect 14565 8517 14599 8551
rect 26617 8517 26651 8551
rect 1777 8449 1811 8483
rect 7481 8449 7515 8483
rect 8125 8449 8159 8483
rect 8767 8449 8801 8483
rect 9873 8449 9907 8483
rect 10701 8449 10735 8483
rect 11161 8449 11195 8483
rect 13277 8449 13311 8483
rect 13921 8449 13955 8483
rect 15853 8449 15887 8483
rect 17141 8449 17175 8483
rect 17785 8449 17819 8483
rect 19993 8449 20027 8483
rect 20637 8449 20671 8483
rect 21281 8449 21315 8483
rect 22017 8449 22051 8483
rect 28273 8449 28307 8483
rect 8953 8381 8987 8415
rect 10517 8381 10551 8415
rect 11805 8381 11839 8415
rect 11989 8381 12023 8415
rect 14473 8381 14507 8415
rect 14749 8381 14783 8415
rect 18061 8381 18095 8415
rect 19533 8381 19567 8415
rect 22293 8381 22327 8415
rect 24593 8381 24627 8415
rect 24869 8381 24903 8415
rect 9965 8313 9999 8347
rect 13093 8313 13127 8347
rect 13737 8313 13771 8347
rect 20729 8313 20763 8347
rect 21373 8313 21407 8347
rect 23765 8313 23799 8347
rect 1593 8245 1627 8279
rect 7573 8245 7607 8279
rect 7849 8041 7883 8075
rect 12449 8041 12483 8075
rect 23397 8041 23431 8075
rect 28273 8041 28307 8075
rect 1593 7973 1627 8007
rect 9965 7973 9999 8007
rect 21189 7973 21223 8007
rect 11253 7905 11287 7939
rect 13553 7905 13587 7939
rect 16313 7905 16347 7939
rect 18153 7905 18187 7939
rect 19441 7905 19475 7939
rect 21649 7905 21683 7939
rect 21925 7905 21959 7939
rect 26525 7905 26559 7939
rect 1777 7837 1811 7871
rect 6653 7837 6687 7871
rect 7113 7837 7147 7871
rect 7757 7837 7791 7871
rect 8585 7837 8619 7871
rect 9505 7837 9539 7871
rect 10149 7837 10183 7871
rect 10609 7837 10643 7871
rect 10793 7837 10827 7871
rect 11805 7837 11839 7871
rect 12633 7837 12667 7871
rect 23857 7837 23891 7871
rect 24777 7837 24811 7871
rect 14841 7769 14875 7803
rect 14933 7769 14967 7803
rect 15485 7769 15519 7803
rect 16405 7769 16439 7803
rect 16957 7769 16991 7803
rect 17877 7769 17911 7803
rect 17969 7769 18003 7803
rect 19717 7769 19751 7803
rect 26801 7769 26835 7803
rect 6469 7701 6503 7735
rect 7205 7701 7239 7735
rect 8401 7701 8435 7735
rect 9321 7701 9355 7735
rect 11897 7701 11931 7735
rect 23949 7701 23983 7735
rect 24593 7701 24627 7735
rect 12357 7497 12391 7531
rect 18429 7497 18463 7531
rect 20913 7497 20947 7531
rect 23305 7497 23339 7531
rect 25881 7497 25915 7531
rect 27629 7497 27663 7531
rect 8493 7429 8527 7463
rect 10425 7429 10459 7463
rect 15669 7429 15703 7463
rect 15761 7429 15795 7463
rect 16313 7429 16347 7463
rect 1593 7361 1627 7395
rect 9781 7361 9815 7395
rect 11897 7361 11931 7395
rect 14473 7361 14507 7395
rect 17969 7361 18003 7395
rect 19165 7361 19199 7395
rect 23213 7361 23247 7395
rect 24133 7361 24167 7395
rect 27537 7361 27571 7395
rect 28181 7361 28215 7395
rect 7665 7293 7699 7327
rect 8401 7293 8435 7327
rect 8677 7293 8711 7327
rect 10333 7293 10367 7327
rect 11713 7293 11747 7327
rect 13001 7293 13035 7327
rect 13185 7293 13219 7327
rect 14289 7293 14323 7327
rect 17325 7293 17359 7327
rect 17509 7293 17543 7327
rect 19441 7293 19475 7327
rect 22109 7293 22143 7327
rect 22293 7293 22327 7327
rect 24409 7293 24443 7327
rect 10885 7225 10919 7259
rect 1777 7157 1811 7191
rect 9597 7157 9631 7191
rect 13645 7157 13679 7191
rect 14749 7157 14783 7191
rect 22477 7157 22511 7191
rect 28273 7157 28307 7191
rect 8401 6953 8435 6987
rect 11437 6953 11471 6987
rect 18429 6953 18463 6987
rect 12357 6885 12391 6919
rect 9413 6817 9447 6851
rect 10057 6817 10091 6851
rect 16681 6817 16715 6851
rect 19533 6817 19567 6851
rect 21281 6817 21315 6851
rect 22201 6817 22235 6851
rect 23765 6817 23799 6851
rect 27169 6817 27203 6851
rect 7941 6749 7975 6783
rect 8585 6749 8619 6783
rect 9597 6749 9631 6783
rect 10793 6749 10827 6783
rect 11437 6749 11471 6783
rect 12541 6749 12575 6783
rect 13001 6749 13035 6783
rect 14933 6749 14967 6783
rect 15577 6749 15611 6783
rect 16037 6749 16071 6783
rect 16221 6749 16255 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 17785 6749 17819 6783
rect 18613 6749 18647 6783
rect 19441 6749 19475 6783
rect 24869 6749 24903 6783
rect 27077 6749 27111 6783
rect 28365 6749 28399 6783
rect 13093 6681 13127 6715
rect 17877 6681 17911 6715
rect 20637 6681 20671 6715
rect 20729 6681 20763 6715
rect 21833 6681 21867 6715
rect 21925 6681 21959 6715
rect 23121 6681 23155 6715
rect 23213 6681 23247 6715
rect 25145 6681 25179 6715
rect 7757 6613 7791 6647
rect 10609 6613 10643 6647
rect 14749 6613 14783 6647
rect 15393 6613 15427 6647
rect 26617 6613 26651 6647
rect 28181 6613 28215 6647
rect 8033 6409 8067 6443
rect 10425 6409 10459 6443
rect 15393 6409 15427 6443
rect 16221 6409 16255 6443
rect 19165 6409 19199 6443
rect 20821 6409 20855 6443
rect 27169 6409 27203 6443
rect 7481 6341 7515 6375
rect 17509 6341 17543 6375
rect 20269 6341 20303 6375
rect 22109 6341 22143 6375
rect 22845 6341 22879 6375
rect 23397 6341 23431 6375
rect 25421 6341 25455 6375
rect 1593 6273 1627 6307
rect 4353 6273 4387 6307
rect 7389 6273 7423 6307
rect 8217 6273 8251 6307
rect 9045 6273 9079 6307
rect 9873 6273 9907 6307
rect 10333 6273 10367 6307
rect 11161 6273 11195 6307
rect 11897 6273 11931 6307
rect 12725 6273 12759 6307
rect 13645 6273 13679 6307
rect 14933 6273 14967 6307
rect 16129 6273 16163 6307
rect 19809 6273 19843 6307
rect 20729 6273 20763 6307
rect 22017 6273 22051 6307
rect 24133 6273 24167 6307
rect 26617 6273 26651 6307
rect 27353 6273 27387 6307
rect 28089 6273 28123 6307
rect 9137 6205 9171 6239
rect 12541 6205 12575 6239
rect 13185 6205 13219 6239
rect 13829 6205 13863 6239
rect 14749 6205 14783 6239
rect 17417 6205 17451 6239
rect 18521 6205 18555 6239
rect 18705 6205 18739 6239
rect 19625 6205 19659 6239
rect 22753 6205 22787 6239
rect 24225 6205 24259 6239
rect 25329 6205 25363 6239
rect 25697 6205 25731 6239
rect 1777 6137 1811 6171
rect 10977 6137 11011 6171
rect 14013 6137 14047 6171
rect 17969 6137 18003 6171
rect 28273 6137 28307 6171
rect 4169 6069 4203 6103
rect 9689 6069 9723 6103
rect 11989 6069 12023 6103
rect 26433 6069 26467 6103
rect 5273 5865 5307 5899
rect 10701 5865 10735 5899
rect 14381 5865 14415 5899
rect 23029 5865 23063 5899
rect 25329 5865 25363 5899
rect 26617 5865 26651 5899
rect 27261 5865 27295 5899
rect 9965 5797 9999 5831
rect 13093 5797 13127 5831
rect 15577 5797 15611 5831
rect 22385 5797 22419 5831
rect 24685 5797 24719 5831
rect 9413 5729 9447 5763
rect 11253 5729 11287 5763
rect 15025 5729 15059 5763
rect 17509 5729 17543 5763
rect 4721 5661 4755 5695
rect 5181 5661 5215 5695
rect 7849 5661 7883 5695
rect 9321 5661 9355 5695
rect 10149 5661 10183 5695
rect 10609 5661 10643 5695
rect 11437 5661 11471 5695
rect 11897 5661 11931 5695
rect 12725 5661 12759 5695
rect 12909 5661 12943 5695
rect 14289 5661 14323 5695
rect 16405 5661 16439 5695
rect 16497 5661 16531 5695
rect 18705 5661 18739 5695
rect 19993 5661 20027 5695
rect 20177 5661 20211 5695
rect 20637 5661 20671 5695
rect 22293 5661 22327 5695
rect 22937 5661 22971 5695
rect 23581 5661 23615 5695
rect 24593 5661 24627 5695
rect 25237 5661 25271 5695
rect 26065 5661 26099 5695
rect 26525 5661 26559 5695
rect 27169 5661 27203 5695
rect 27813 5661 27847 5695
rect 15117 5593 15151 5627
rect 17601 5593 17635 5627
rect 18153 5593 18187 5627
rect 4537 5525 4571 5559
rect 7941 5525 7975 5559
rect 18797 5525 18831 5559
rect 23673 5525 23707 5559
rect 25881 5525 25915 5559
rect 27905 5525 27939 5559
rect 9321 5321 9355 5355
rect 10057 5321 10091 5355
rect 12357 5321 12391 5355
rect 14197 5321 14231 5355
rect 14841 5321 14875 5355
rect 15485 5321 15519 5355
rect 17877 5321 17911 5355
rect 16221 5253 16255 5287
rect 17233 5253 17267 5287
rect 19349 5253 19383 5287
rect 20913 5253 20947 5287
rect 26065 5253 26099 5287
rect 26617 5253 26651 5287
rect 1593 5185 1627 5219
rect 4169 5185 4203 5219
rect 8861 5185 8895 5219
rect 9505 5185 9539 5219
rect 9965 5185 9999 5219
rect 11161 5185 11195 5219
rect 12265 5185 12299 5219
rect 13093 5185 13127 5219
rect 13737 5185 13771 5219
rect 14381 5185 14415 5219
rect 15669 5185 15703 5219
rect 16129 5185 16163 5219
rect 17141 5185 17175 5219
rect 17785 5185 17819 5219
rect 18521 5185 18555 5219
rect 22569 5185 22603 5219
rect 24041 5185 24075 5219
rect 24961 5185 24995 5219
rect 28089 5185 28123 5219
rect 19257 5117 19291 5151
rect 19533 5117 19567 5151
rect 20821 5117 20855 5151
rect 21097 5117 21131 5151
rect 22753 5117 22787 5151
rect 23857 5117 23891 5151
rect 25973 5117 26007 5151
rect 12909 5049 12943 5083
rect 22937 5049 22971 5083
rect 24225 5049 24259 5083
rect 1777 4981 1811 5015
rect 3985 4981 4019 5015
rect 8677 4981 8711 5015
rect 10977 4981 11011 5015
rect 13553 4981 13587 5015
rect 18613 4981 18647 5015
rect 25053 4981 25087 5015
rect 28273 4981 28307 5015
rect 9137 4777 9171 4811
rect 12173 4777 12207 4811
rect 12909 4777 12943 4811
rect 14289 4777 14323 4811
rect 20729 4777 20763 4811
rect 21373 4777 21407 4811
rect 22385 4777 22419 4811
rect 23029 4777 23063 4811
rect 23673 4777 23707 4811
rect 25237 4777 25271 4811
rect 27629 4777 27663 4811
rect 13553 4709 13587 4743
rect 17601 4709 17635 4743
rect 19809 4709 19843 4743
rect 28273 4709 28307 4743
rect 11805 4641 11839 4675
rect 18521 4641 18555 4675
rect 19441 4641 19475 4675
rect 6193 4573 6227 4607
rect 9321 4573 9355 4607
rect 10977 4573 11011 4607
rect 11621 4573 11655 4607
rect 13093 4573 13127 4607
rect 13737 4573 13771 4607
rect 14473 4573 14507 4607
rect 15209 4573 15243 4607
rect 17233 4573 17267 4607
rect 17417 4573 17451 4607
rect 19625 4573 19659 4607
rect 20637 4573 20671 4607
rect 21281 4573 21315 4607
rect 22293 4573 22327 4607
rect 22937 4573 22971 4607
rect 23581 4573 23615 4607
rect 24593 4573 24627 4607
rect 24777 4573 24811 4607
rect 25881 4573 25915 4607
rect 27537 4573 27571 4607
rect 28181 4573 28215 4607
rect 15301 4505 15335 4539
rect 6009 4437 6043 4471
rect 10333 4437 10367 4471
rect 15853 4437 15887 4471
rect 25697 4437 25731 4471
rect 22201 4233 22235 4267
rect 23949 4233 23983 4267
rect 24685 4233 24719 4267
rect 13553 4165 13587 4199
rect 7573 4097 7607 4131
rect 8401 4097 8435 4131
rect 9045 4097 9079 4131
rect 10517 4097 10551 4131
rect 11161 4097 11195 4131
rect 11713 4097 11747 4131
rect 14105 4097 14139 4131
rect 14749 4097 14783 4131
rect 15485 4097 15519 4131
rect 17049 4097 17083 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 19441 4097 19475 4131
rect 19533 4097 19567 4131
rect 20085 4097 20119 4131
rect 20177 4097 20211 4131
rect 20913 4097 20947 4131
rect 22385 4097 22419 4131
rect 23305 4097 23339 4131
rect 23397 4097 23431 4131
rect 24593 4097 24627 4131
rect 27169 4097 27203 4131
rect 27813 4097 27847 4131
rect 11897 4029 11931 4063
rect 13461 4029 13495 4063
rect 15669 4029 15703 4063
rect 27905 4029 27939 4063
rect 8217 3961 8251 3995
rect 8861 3961 8895 3995
rect 10333 3961 10367 3995
rect 15853 3961 15887 3995
rect 17693 3961 17727 3995
rect 18337 3961 18371 3995
rect 7665 3893 7699 3927
rect 10977 3893 11011 3927
rect 12173 3893 12207 3927
rect 14565 3893 14599 3927
rect 17141 3893 17175 3927
rect 20729 3893 20763 3927
rect 27261 3893 27295 3927
rect 12449 3689 12483 3723
rect 13461 3689 13495 3723
rect 14749 3689 14783 3723
rect 15577 3689 15611 3723
rect 18705 3689 18739 3723
rect 22385 3689 22419 3723
rect 23765 3689 23799 3723
rect 25237 3689 25271 3723
rect 26249 3689 26283 3723
rect 26801 3689 26835 3723
rect 11805 3621 11839 3655
rect 18153 3621 18187 3655
rect 19441 3621 19475 3655
rect 21189 3621 21223 3655
rect 14473 3553 14507 3587
rect 20637 3553 20671 3587
rect 21741 3553 21775 3587
rect 25605 3553 25639 3587
rect 25789 3553 25823 3587
rect 1593 3485 1627 3519
rect 11989 3485 12023 3519
rect 12633 3485 12667 3519
rect 13645 3485 13679 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 17049 3485 17083 3519
rect 18061 3485 18095 3519
rect 18889 3485 18923 3519
rect 19625 3485 19659 3519
rect 22569 3485 22603 3519
rect 23673 3485 23707 3519
rect 26985 3485 27019 3519
rect 27629 3485 27663 3519
rect 28089 3485 28123 3519
rect 20706 3417 20740 3451
rect 1777 3349 1811 3383
rect 16865 3349 16899 3383
rect 27445 3349 27479 3383
rect 28273 3349 28307 3383
rect 2329 3145 2363 3179
rect 9413 3145 9447 3179
rect 13645 3145 13679 3179
rect 18245 3145 18279 3179
rect 20637 3145 20671 3179
rect 22017 3145 22051 3179
rect 23397 3145 23431 3179
rect 25513 3145 25547 3179
rect 27445 3145 27479 3179
rect 12725 3077 12759 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3157 3009 3191 3043
rect 5733 3009 5767 3043
rect 8861 3009 8895 3043
rect 8953 3009 8987 3043
rect 9597 3009 9631 3043
rect 10425 3009 10459 3043
rect 11161 3009 11195 3043
rect 11989 3009 12023 3043
rect 12633 3009 12667 3043
rect 13829 3009 13863 3043
rect 14841 3009 14875 3043
rect 15761 3009 15795 3043
rect 17049 3009 17083 3043
rect 17509 3009 17543 3043
rect 17601 3009 17635 3043
rect 18153 3009 18187 3043
rect 18981 3009 19015 3043
rect 20821 3009 20855 3043
rect 21281 3009 21315 3043
rect 22201 3009 22235 3043
rect 22661 3009 22695 3043
rect 23305 3009 23339 3043
rect 24225 3009 24259 3043
rect 24317 3009 24351 3043
rect 25053 3009 25087 3043
rect 25697 3009 25731 3043
rect 26433 3009 26467 3043
rect 27629 3009 27663 3043
rect 28089 3009 28123 3043
rect 12081 2941 12115 2975
rect 15853 2941 15887 2975
rect 19533 2941 19567 2975
rect 19717 2941 19751 2975
rect 21373 2941 21407 2975
rect 2973 2873 3007 2907
rect 10977 2873 11011 2907
rect 26249 2873 26283 2907
rect 1777 2805 1811 2839
rect 5549 2805 5583 2839
rect 10241 2805 10275 2839
rect 14657 2805 14691 2839
rect 16865 2805 16899 2839
rect 18797 2805 18831 2839
rect 19901 2805 19935 2839
rect 22753 2805 22787 2839
rect 24869 2805 24903 2839
rect 28273 2805 28307 2839
rect 7849 2601 7883 2635
rect 9137 2601 9171 2635
rect 11713 2601 11747 2635
rect 16865 2601 16899 2635
rect 18245 2601 18279 2635
rect 19717 2601 19751 2635
rect 20545 2601 20579 2635
rect 22661 2601 22695 2635
rect 24593 2601 24627 2635
rect 25881 2601 25915 2635
rect 27169 2601 27203 2635
rect 21097 2533 21131 2567
rect 23305 2533 23339 2567
rect 25237 2533 25271 2567
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 3157 2397 3191 2431
rect 4629 2397 4663 2431
rect 5733 2397 5767 2431
rect 6561 2397 6595 2431
rect 8033 2397 8067 2431
rect 9321 2397 9355 2431
rect 10425 2397 10459 2431
rect 11897 2397 11931 2431
rect 12725 2397 12759 2431
rect 13461 2397 13495 2431
rect 14933 2397 14967 2431
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 19901 2397 19935 2431
rect 20453 2397 20487 2431
rect 21281 2397 21315 2431
rect 22201 2397 22235 2431
rect 22845 2397 22879 2431
rect 23489 2397 23523 2431
rect 24777 2397 24811 2431
rect 25421 2397 25455 2431
rect 26065 2397 26099 2431
rect 27353 2397 27387 2431
rect 27813 2397 27847 2431
rect 1777 2261 1811 2295
rect 2329 2261 2363 2295
rect 3341 2261 3375 2295
rect 4813 2261 4847 2295
rect 5917 2261 5951 2295
rect 6745 2261 6779 2295
rect 10609 2261 10643 2295
rect 12909 2261 12943 2295
rect 13645 2261 13679 2295
rect 15117 2261 15151 2295
rect 17693 2261 17727 2295
rect 22017 2261 22051 2295
rect 27997 2261 28031 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 24504 27628 24716 27656
rect 1026 27548 1032 27600
rect 1084 27588 1090 27600
rect 2501 27591 2559 27597
rect 2501 27588 2513 27591
rect 1084 27560 2513 27588
rect 1084 27548 1090 27560
rect 2501 27557 2513 27560
rect 2547 27557 2559 27591
rect 2501 27551 2559 27557
rect 3237 27591 3295 27597
rect 3237 27557 3249 27591
rect 3283 27557 3295 27591
rect 3237 27551 3295 27557
rect 3973 27591 4031 27597
rect 3973 27557 3985 27591
rect 4019 27588 4031 27591
rect 6086 27588 6092 27600
rect 4019 27560 6092 27588
rect 4019 27557 4031 27560
rect 3973 27551 4031 27557
rect 3252 27520 3280 27551
rect 6086 27548 6092 27560
rect 6144 27548 6150 27600
rect 7837 27591 7895 27597
rect 7837 27557 7849 27591
rect 7883 27557 7895 27591
rect 7837 27551 7895 27557
rect 7282 27520 7288 27532
rect 3252 27492 7288 27520
rect 7282 27480 7288 27492
rect 7340 27480 7346 27532
rect 7852 27520 7880 27551
rect 10318 27548 10324 27600
rect 10376 27588 10382 27600
rect 10597 27591 10655 27597
rect 10597 27588 10609 27591
rect 10376 27560 10609 27588
rect 10376 27548 10382 27560
rect 10597 27557 10609 27560
rect 10643 27557 10655 27591
rect 10597 27551 10655 27557
rect 13538 27548 13544 27600
rect 13596 27588 13602 27600
rect 13633 27591 13691 27597
rect 13633 27588 13645 27591
rect 13596 27560 13645 27588
rect 13596 27548 13602 27560
rect 13633 27557 13645 27560
rect 13679 27557 13691 27591
rect 15102 27588 15108 27600
rect 15063 27560 15108 27588
rect 13633 27551 13691 27557
rect 15102 27548 15108 27560
rect 15160 27548 15166 27600
rect 16114 27548 16120 27600
rect 16172 27588 16178 27600
rect 17037 27591 17095 27597
rect 17037 27588 17049 27591
rect 16172 27560 17049 27588
rect 16172 27548 16178 27560
rect 17037 27557 17049 27560
rect 17083 27557 17095 27591
rect 17037 27551 17095 27557
rect 18046 27548 18052 27600
rect 18104 27588 18110 27600
rect 18325 27591 18383 27597
rect 18325 27588 18337 27591
rect 18104 27560 18337 27588
rect 18104 27548 18110 27560
rect 18325 27557 18337 27560
rect 18371 27557 18383 27591
rect 18325 27551 18383 27557
rect 19429 27591 19487 27597
rect 19429 27557 19441 27591
rect 19475 27557 19487 27591
rect 19429 27551 19487 27557
rect 7852 27492 14320 27520
rect 2317 27455 2375 27461
rect 2317 27421 2329 27455
rect 2363 27452 2375 27455
rect 3234 27452 3240 27464
rect 2363 27424 3240 27452
rect 2363 27421 2375 27424
rect 2317 27415 2375 27421
rect 3234 27412 3240 27424
rect 3292 27412 3298 27464
rect 3418 27452 3424 27464
rect 3379 27424 3424 27452
rect 3418 27412 3424 27424
rect 3476 27412 3482 27464
rect 4154 27452 4160 27464
rect 4115 27424 4160 27452
rect 4154 27412 4160 27424
rect 4212 27412 4218 27464
rect 5442 27452 5448 27464
rect 5403 27424 5448 27452
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 6730 27452 6736 27464
rect 6691 27424 6736 27452
rect 6730 27412 6736 27424
rect 6788 27412 6794 27464
rect 8018 27452 8024 27464
rect 7979 27424 8024 27452
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 9030 27412 9036 27464
rect 9088 27452 9094 27464
rect 9309 27455 9367 27461
rect 9309 27452 9321 27455
rect 9088 27424 9321 27452
rect 9088 27412 9094 27424
rect 9309 27421 9321 27424
rect 9355 27421 9367 27455
rect 10410 27452 10416 27464
rect 10371 27424 10416 27452
rect 9309 27415 9367 27421
rect 10410 27412 10416 27424
rect 10468 27412 10474 27464
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 11885 27455 11943 27461
rect 11885 27452 11897 27455
rect 11112 27424 11897 27452
rect 11112 27412 11118 27424
rect 11885 27421 11897 27424
rect 11931 27421 11943 27455
rect 11885 27415 11943 27421
rect 12434 27412 12440 27464
rect 12492 27452 12498 27464
rect 12529 27455 12587 27461
rect 12529 27452 12541 27455
rect 12492 27424 12541 27452
rect 12492 27412 12498 27424
rect 12529 27421 12541 27424
rect 12575 27421 12587 27455
rect 12529 27415 12587 27421
rect 13170 27412 13176 27464
rect 13228 27452 13234 27464
rect 14292 27461 14320 27492
rect 13449 27455 13507 27461
rect 13449 27452 13461 27455
rect 13228 27424 13461 27452
rect 13228 27412 13234 27424
rect 13449 27421 13461 27424
rect 13495 27421 13507 27455
rect 13449 27415 13507 27421
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14366 27412 14372 27464
rect 14424 27452 14430 27464
rect 14921 27455 14979 27461
rect 14921 27452 14933 27455
rect 14424 27424 14933 27452
rect 14424 27412 14430 27424
rect 14921 27421 14933 27424
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 15841 27455 15899 27461
rect 15841 27421 15853 27455
rect 15887 27421 15899 27455
rect 16850 27452 16856 27464
rect 16811 27424 16856 27452
rect 15841 27415 15899 27421
rect 1670 27384 1676 27396
rect 1631 27356 1676 27384
rect 1670 27344 1676 27356
rect 1728 27344 1734 27396
rect 1854 27384 1860 27396
rect 1815 27356 1860 27384
rect 1854 27344 1860 27356
rect 1912 27344 1918 27396
rect 11974 27384 11980 27396
rect 6564 27356 11980 27384
rect 5261 27319 5319 27325
rect 5261 27285 5273 27319
rect 5307 27316 5319 27319
rect 6454 27316 6460 27328
rect 5307 27288 6460 27316
rect 5307 27285 5319 27288
rect 5261 27279 5319 27285
rect 6454 27276 6460 27288
rect 6512 27276 6518 27328
rect 6564 27325 6592 27356
rect 11974 27344 11980 27356
rect 12032 27344 12038 27396
rect 15856 27384 15884 27415
rect 16850 27412 16856 27424
rect 16908 27412 16914 27464
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 19444 27452 19472 27551
rect 20714 27548 20720 27600
rect 20772 27588 20778 27600
rect 20901 27591 20959 27597
rect 20901 27588 20913 27591
rect 20772 27560 20913 27588
rect 20772 27548 20778 27560
rect 20901 27557 20913 27560
rect 20947 27557 20959 27591
rect 20901 27551 20959 27557
rect 23474 27548 23480 27600
rect 23532 27588 23538 27600
rect 24504 27588 24532 27628
rect 23532 27560 24532 27588
rect 24581 27591 24639 27597
rect 23532 27548 23538 27560
rect 24581 27557 24593 27591
rect 24627 27557 24639 27591
rect 24581 27551 24639 27557
rect 19610 27452 19616 27464
rect 18187 27424 19472 27452
rect 19571 27424 19616 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 20073 27455 20131 27461
rect 20073 27421 20085 27455
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27452 20775 27455
rect 21358 27452 21364 27464
rect 20763 27424 21364 27452
rect 20763 27421 20775 27424
rect 20717 27415 20775 27421
rect 17770 27384 17776 27396
rect 15856 27356 17776 27384
rect 17770 27344 17776 27356
rect 17828 27344 17834 27396
rect 6549 27319 6607 27325
rect 6549 27285 6561 27319
rect 6595 27285 6607 27319
rect 6549 27279 6607 27285
rect 9125 27319 9183 27325
rect 9125 27285 9137 27319
rect 9171 27316 9183 27319
rect 9582 27316 9588 27328
rect 9171 27288 9588 27316
rect 9171 27285 9183 27288
rect 9125 27279 9183 27285
rect 9582 27276 9588 27288
rect 9640 27276 9646 27328
rect 11698 27316 11704 27328
rect 11659 27288 11704 27316
rect 11698 27276 11704 27288
rect 11756 27276 11762 27328
rect 12345 27319 12403 27325
rect 12345 27285 12357 27319
rect 12391 27316 12403 27319
rect 12710 27316 12716 27328
rect 12391 27288 12716 27316
rect 12391 27285 12403 27288
rect 12345 27279 12403 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 14369 27319 14427 27325
rect 14369 27285 14381 27319
rect 14415 27316 14427 27319
rect 14734 27316 14740 27328
rect 14415 27288 14740 27316
rect 14415 27285 14427 27288
rect 14369 27279 14427 27285
rect 14734 27276 14740 27288
rect 14792 27276 14798 27328
rect 15654 27316 15660 27328
rect 15615 27288 15660 27316
rect 15654 27276 15660 27288
rect 15712 27276 15718 27328
rect 15930 27276 15936 27328
rect 15988 27316 15994 27328
rect 20088 27316 20116 27415
rect 21358 27412 21364 27424
rect 21416 27412 21422 27464
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 22833 27455 22891 27461
rect 22833 27452 22845 27455
rect 22152 27424 22845 27452
rect 22152 27412 22158 27424
rect 22833 27421 22845 27424
rect 22879 27421 22891 27455
rect 22833 27415 22891 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27452 23351 27455
rect 24596 27452 24624 27551
rect 23339 27424 24624 27452
rect 24688 27452 24716 27628
rect 27522 27616 27528 27668
rect 27580 27656 27586 27668
rect 29270 27656 29276 27668
rect 27580 27628 29276 27656
rect 27580 27616 27586 27628
rect 29270 27616 29276 27628
rect 29328 27616 29334 27668
rect 27706 27548 27712 27600
rect 27764 27588 27770 27600
rect 27985 27591 28043 27597
rect 27985 27588 27997 27591
rect 27764 27560 27997 27588
rect 27764 27548 27770 27560
rect 27985 27557 27997 27560
rect 28031 27557 28043 27591
rect 27985 27551 28043 27557
rect 25130 27480 25136 27532
rect 25188 27520 25194 27532
rect 25188 27492 26096 27520
rect 25188 27480 25194 27492
rect 26068 27461 26096 27492
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 24688 27424 24777 27452
rect 23339 27421 23351 27424
rect 23293 27415 23351 27421
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 24210 27344 24216 27396
rect 24268 27384 24274 27396
rect 25424 27384 25452 27415
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 27341 27455 27399 27461
rect 27341 27452 27353 27455
rect 26476 27424 27353 27452
rect 26476 27412 26482 27424
rect 27341 27421 27353 27424
rect 27387 27421 27399 27455
rect 27341 27415 27399 27421
rect 27430 27412 27436 27464
rect 27488 27452 27494 27464
rect 27801 27455 27859 27461
rect 27801 27452 27813 27455
rect 27488 27424 27813 27452
rect 27488 27412 27494 27424
rect 27801 27421 27813 27424
rect 27847 27421 27859 27455
rect 27801 27415 27859 27421
rect 24268 27356 25452 27384
rect 24268 27344 24274 27356
rect 15988 27288 20116 27316
rect 20165 27319 20223 27325
rect 15988 27276 15994 27288
rect 20165 27285 20177 27319
rect 20211 27316 20223 27319
rect 21542 27316 21548 27328
rect 20211 27288 21548 27316
rect 20211 27285 20223 27288
rect 20165 27279 20223 27285
rect 21542 27276 21548 27288
rect 21600 27276 21606 27328
rect 21634 27276 21640 27328
rect 21692 27316 21698 27328
rect 22005 27319 22063 27325
rect 22005 27316 22017 27319
rect 21692 27288 22017 27316
rect 21692 27276 21698 27288
rect 22005 27285 22017 27288
rect 22051 27285 22063 27319
rect 22646 27316 22652 27328
rect 22607 27288 22652 27316
rect 22005 27279 22063 27285
rect 22646 27276 22652 27288
rect 22704 27276 22710 27328
rect 23382 27316 23388 27328
rect 23343 27288 23388 27316
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 25038 27276 25044 27328
rect 25096 27316 25102 27328
rect 25225 27319 25283 27325
rect 25225 27316 25237 27319
rect 25096 27288 25237 27316
rect 25096 27276 25102 27288
rect 25225 27285 25237 27288
rect 25271 27285 25283 27319
rect 25225 27279 25283 27285
rect 25590 27276 25596 27328
rect 25648 27316 25654 27328
rect 25869 27319 25927 27325
rect 25869 27316 25881 27319
rect 25648 27288 25881 27316
rect 25648 27276 25654 27288
rect 25869 27285 25881 27288
rect 25915 27285 25927 27319
rect 27154 27316 27160 27328
rect 27115 27288 27160 27316
rect 25869 27279 25927 27285
rect 27154 27276 27160 27288
rect 27212 27276 27218 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 1765 27115 1823 27121
rect 1765 27081 1777 27115
rect 1811 27112 1823 27115
rect 2774 27112 2780 27124
rect 1811 27084 2780 27112
rect 1811 27081 1823 27084
rect 1765 27075 1823 27081
rect 2774 27072 2780 27084
rect 2832 27072 2838 27124
rect 3234 27072 3240 27124
rect 3292 27112 3298 27124
rect 3881 27115 3939 27121
rect 3881 27112 3893 27115
rect 3292 27084 3893 27112
rect 3292 27072 3298 27084
rect 3881 27081 3893 27084
rect 3927 27081 3939 27115
rect 13170 27112 13176 27124
rect 13131 27084 13176 27112
rect 3881 27075 3939 27081
rect 13170 27072 13176 27084
rect 13228 27072 13234 27124
rect 19334 27112 19340 27124
rect 16684 27084 19340 27112
rect 15654 27044 15660 27056
rect 14016 27016 15660 27044
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26945 1639 26979
rect 1581 26939 1639 26945
rect 1596 26908 1624 26939
rect 1946 26936 1952 26988
rect 2004 26976 2010 26988
rect 2501 26979 2559 26985
rect 2501 26976 2513 26979
rect 2004 26948 2513 26976
rect 2004 26936 2010 26948
rect 2501 26945 2513 26948
rect 2547 26945 2559 26979
rect 3142 26976 3148 26988
rect 3103 26948 3148 26976
rect 2501 26939 2559 26945
rect 3142 26936 3148 26948
rect 3200 26936 3206 26988
rect 4065 26979 4123 26985
rect 4065 26945 4077 26979
rect 4111 26976 4123 26979
rect 4246 26976 4252 26988
rect 4111 26948 4252 26976
rect 4111 26945 4123 26948
rect 4065 26939 4123 26945
rect 4246 26936 4252 26948
rect 4304 26936 4310 26988
rect 13357 26979 13415 26985
rect 13357 26945 13369 26979
rect 13403 26976 13415 26979
rect 13906 26976 13912 26988
rect 13403 26948 13912 26976
rect 13403 26945 13415 26948
rect 13357 26939 13415 26945
rect 13906 26936 13912 26948
rect 13964 26936 13970 26988
rect 14016 26985 14044 27016
rect 15654 27004 15660 27016
rect 15712 27004 15718 27056
rect 14001 26979 14059 26985
rect 14001 26945 14013 26979
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14461 26979 14519 26985
rect 14461 26945 14473 26979
rect 14507 26945 14519 26979
rect 14461 26939 14519 26945
rect 4890 26908 4896 26920
rect 1596 26880 4896 26908
rect 4890 26868 4896 26880
rect 4948 26868 4954 26920
rect 11701 26911 11759 26917
rect 11701 26877 11713 26911
rect 11747 26908 11759 26911
rect 11790 26908 11796 26920
rect 11747 26880 11796 26908
rect 11747 26877 11759 26880
rect 11701 26871 11759 26877
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 14476 26908 14504 26939
rect 14734 26936 14740 26988
rect 14792 26976 14798 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14792 26948 15117 26976
rect 14792 26936 14798 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 16684 26976 16712 27084
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 27522 27112 27528 27124
rect 27483 27084 27528 27112
rect 27522 27072 27528 27084
rect 27580 27072 27586 27124
rect 28261 27115 28319 27121
rect 28261 27081 28273 27115
rect 28307 27112 28319 27115
rect 29914 27112 29920 27124
rect 28307 27084 29920 27112
rect 28307 27081 28319 27084
rect 28261 27075 28319 27081
rect 29914 27072 29920 27084
rect 29972 27072 29978 27124
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 16816 27016 18644 27044
rect 16816 27004 16822 27016
rect 15105 26939 15163 26945
rect 15212 26948 16712 26976
rect 16853 26979 16911 26985
rect 15212 26908 15240 26948
rect 16853 26945 16865 26979
rect 16899 26976 16911 26979
rect 17126 26976 17132 26988
rect 16899 26948 17132 26976
rect 16899 26945 16911 26948
rect 16853 26939 16911 26945
rect 17126 26936 17132 26948
rect 17184 26936 17190 26988
rect 17770 26976 17776 26988
rect 17683 26948 17776 26976
rect 17770 26936 17776 26948
rect 17828 26936 17834 26988
rect 18616 26985 18644 27016
rect 18782 27004 18788 27056
rect 18840 27044 18846 27056
rect 20717 27047 20775 27053
rect 20717 27044 20729 27047
rect 18840 27016 20729 27044
rect 18840 27004 18846 27016
rect 20717 27013 20729 27016
rect 20763 27013 20775 27047
rect 20717 27007 20775 27013
rect 22646 27004 22652 27056
rect 22704 27044 22710 27056
rect 27154 27044 27160 27056
rect 22704 27016 23796 27044
rect 22704 27004 22710 27016
rect 18601 26979 18659 26985
rect 18601 26945 18613 26979
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 19245 26979 19303 26985
rect 19245 26945 19257 26979
rect 19291 26976 19303 26979
rect 19426 26976 19432 26988
rect 19291 26948 19432 26976
rect 19291 26945 19303 26948
rect 19245 26939 19303 26945
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19702 26936 19708 26988
rect 19760 26976 19766 26988
rect 21361 26979 21419 26985
rect 21361 26976 21373 26979
rect 19760 26948 21373 26976
rect 19760 26936 19766 26948
rect 21361 26945 21373 26948
rect 21407 26945 21419 26979
rect 21361 26939 21419 26945
rect 21634 26936 21640 26988
rect 21692 26976 21698 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21692 26948 22017 26976
rect 21692 26936 21698 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 23014 26936 23020 26988
rect 23072 26976 23078 26988
rect 23768 26985 23796 27016
rect 24412 27016 27160 27044
rect 24412 26985 24440 27016
rect 27154 27004 27160 27016
rect 27212 27004 27218 27056
rect 23293 26979 23351 26985
rect 23293 26976 23305 26979
rect 23072 26948 23305 26976
rect 23072 26936 23078 26948
rect 23293 26945 23305 26948
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 23753 26979 23811 26985
rect 23753 26945 23765 26979
rect 23799 26945 23811 26979
rect 23753 26939 23811 26945
rect 24397 26979 24455 26985
rect 24397 26945 24409 26979
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 25501 26979 25559 26985
rect 25501 26945 25513 26979
rect 25547 26945 25559 26979
rect 25501 26939 25559 26945
rect 25961 26979 26019 26985
rect 25961 26945 25973 26979
rect 26007 26976 26019 26979
rect 26510 26976 26516 26988
rect 26007 26948 26516 26976
rect 26007 26945 26019 26948
rect 25961 26939 26019 26945
rect 14476 26880 15240 26908
rect 15289 26911 15347 26917
rect 15289 26877 15301 26911
rect 15335 26908 15347 26911
rect 16942 26908 16948 26920
rect 15335 26880 16948 26908
rect 15335 26877 15347 26880
rect 15289 26871 15347 26877
rect 16942 26868 16948 26880
rect 17000 26868 17006 26920
rect 17037 26911 17095 26917
rect 17037 26877 17049 26911
rect 17083 26908 17095 26911
rect 17678 26908 17684 26920
rect 17083 26880 17684 26908
rect 17083 26877 17095 26880
rect 17037 26871 17095 26877
rect 17678 26868 17684 26880
rect 17736 26868 17742 26920
rect 17788 26908 17816 26936
rect 20073 26911 20131 26917
rect 17788 26880 19196 26908
rect 2317 26843 2375 26849
rect 2317 26809 2329 26843
rect 2363 26840 2375 26843
rect 8294 26840 8300 26852
rect 2363 26812 8300 26840
rect 2363 26809 2375 26812
rect 2317 26803 2375 26809
rect 8294 26800 8300 26812
rect 8352 26800 8358 26852
rect 10410 26800 10416 26852
rect 10468 26840 10474 26852
rect 14274 26840 14280 26852
rect 10468 26812 14280 26840
rect 10468 26800 10474 26812
rect 14274 26800 14280 26812
rect 14332 26800 14338 26852
rect 16114 26800 16120 26852
rect 16172 26840 16178 26852
rect 18417 26843 18475 26849
rect 18417 26840 18429 26843
rect 16172 26812 18429 26840
rect 16172 26800 16178 26812
rect 18417 26809 18429 26812
rect 18463 26809 18475 26843
rect 18417 26803 18475 26809
rect 2961 26775 3019 26781
rect 2961 26741 2973 26775
rect 3007 26772 3019 26775
rect 10226 26772 10232 26784
rect 3007 26744 10232 26772
rect 3007 26741 3019 26744
rect 2961 26735 3019 26741
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 13814 26772 13820 26784
rect 13775 26744 13820 26772
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 14550 26772 14556 26784
rect 14511 26744 14556 26772
rect 14550 26732 14556 26744
rect 14608 26732 14614 26784
rect 15746 26772 15752 26784
rect 15707 26744 15752 26772
rect 15746 26732 15752 26744
rect 15804 26732 15810 26784
rect 16666 26732 16672 26784
rect 16724 26772 16730 26784
rect 17865 26775 17923 26781
rect 17865 26772 17877 26775
rect 16724 26744 17877 26772
rect 16724 26732 16730 26744
rect 17865 26741 17877 26744
rect 17911 26741 17923 26775
rect 17865 26735 17923 26741
rect 18690 26732 18696 26784
rect 18748 26772 18754 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 18748 26744 19073 26772
rect 18748 26732 18754 26744
rect 19061 26741 19073 26744
rect 19107 26741 19119 26775
rect 19168 26772 19196 26880
rect 20073 26877 20085 26911
rect 20119 26877 20131 26911
rect 20073 26871 20131 26877
rect 20257 26911 20315 26917
rect 20257 26877 20269 26911
rect 20303 26908 20315 26911
rect 20714 26908 20720 26920
rect 20303 26880 20720 26908
rect 20303 26877 20315 26880
rect 20257 26871 20315 26877
rect 19702 26800 19708 26852
rect 19760 26840 19766 26852
rect 20088 26840 20116 26871
rect 20714 26868 20720 26880
rect 20772 26868 20778 26920
rect 22189 26911 22247 26917
rect 22189 26877 22201 26911
rect 22235 26908 22247 26911
rect 22646 26908 22652 26920
rect 22235 26880 22652 26908
rect 22235 26877 22247 26880
rect 22189 26871 22247 26877
rect 22646 26868 22652 26880
rect 22704 26868 22710 26920
rect 25516 26908 25544 26939
rect 26510 26936 26516 26948
rect 26568 26936 26574 26988
rect 27338 26976 27344 26988
rect 27299 26948 27344 26976
rect 27338 26936 27344 26948
rect 27396 26936 27402 26988
rect 27522 26936 27528 26988
rect 27580 26976 27586 26988
rect 28077 26979 28135 26985
rect 28077 26976 28089 26979
rect 27580 26948 28089 26976
rect 27580 26936 27586 26948
rect 28077 26945 28089 26948
rect 28123 26945 28135 26979
rect 28077 26939 28135 26945
rect 27890 26908 27896 26920
rect 25516 26880 27896 26908
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 23382 26840 23388 26852
rect 19760 26812 23388 26840
rect 19760 26800 19766 26812
rect 23382 26800 23388 26812
rect 23440 26800 23446 26852
rect 19886 26772 19892 26784
rect 19168 26744 19892 26772
rect 19061 26735 19119 26741
rect 19886 26732 19892 26744
rect 19944 26732 19950 26784
rect 21174 26772 21180 26784
rect 21135 26744 21180 26772
rect 21174 26732 21180 26744
rect 21232 26732 21238 26784
rect 22554 26772 22560 26784
rect 22515 26744 22560 26772
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 23109 26775 23167 26781
rect 23109 26772 23121 26775
rect 22796 26744 23121 26772
rect 22796 26732 22802 26744
rect 23109 26741 23121 26744
rect 23155 26741 23167 26775
rect 23842 26772 23848 26784
rect 23803 26744 23848 26772
rect 23109 26735 23167 26741
rect 23842 26732 23848 26744
rect 23900 26732 23906 26784
rect 24486 26772 24492 26784
rect 24447 26744 24492 26772
rect 24486 26732 24492 26744
rect 24544 26732 24550 26784
rect 25317 26775 25375 26781
rect 25317 26741 25329 26775
rect 25363 26772 25375 26775
rect 25958 26772 25964 26784
rect 25363 26744 25964 26772
rect 25363 26741 25375 26744
rect 25317 26735 25375 26741
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 26050 26732 26056 26784
rect 26108 26772 26114 26784
rect 26108 26744 26153 26772
rect 26108 26732 26114 26744
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 1581 26571 1639 26577
rect 1581 26537 1593 26571
rect 1627 26568 1639 26571
rect 4246 26568 4252 26580
rect 1627 26540 2774 26568
rect 4207 26540 4252 26568
rect 1627 26537 1639 26540
rect 1581 26531 1639 26537
rect 2746 26500 2774 26540
rect 4246 26528 4252 26540
rect 4304 26528 4310 26580
rect 4890 26568 4896 26580
rect 4851 26540 4896 26568
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 10689 26571 10747 26577
rect 10689 26537 10701 26571
rect 10735 26568 10747 26571
rect 11882 26568 11888 26580
rect 10735 26540 11888 26568
rect 10735 26537 10747 26540
rect 10689 26531 10747 26537
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 18785 26571 18843 26577
rect 18785 26568 18797 26571
rect 17000 26540 18797 26568
rect 17000 26528 17006 26540
rect 18785 26537 18797 26540
rect 18831 26537 18843 26571
rect 19426 26568 19432 26580
rect 19387 26540 19432 26568
rect 18785 26531 18843 26537
rect 19426 26528 19432 26540
rect 19484 26528 19490 26580
rect 19610 26528 19616 26580
rect 19668 26568 19674 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 19668 26540 20177 26568
rect 19668 26528 19674 26540
rect 20165 26537 20177 26540
rect 20211 26537 20223 26571
rect 20714 26568 20720 26580
rect 20675 26540 20720 26568
rect 20165 26531 20223 26537
rect 20714 26528 20720 26540
rect 20772 26528 20778 26580
rect 21358 26568 21364 26580
rect 21319 26540 21364 26568
rect 21358 26528 21364 26540
rect 21416 26528 21422 26580
rect 22646 26568 22652 26580
rect 22607 26540 22652 26568
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 27338 26568 27344 26580
rect 27299 26540 27344 26568
rect 27338 26528 27344 26540
rect 27396 26528 27402 26580
rect 28261 26571 28319 26577
rect 28261 26537 28273 26571
rect 28307 26568 28319 26571
rect 28626 26568 28632 26580
rect 28307 26540 28632 26568
rect 28307 26537 28319 26540
rect 28261 26531 28319 26537
rect 28626 26528 28632 26540
rect 28684 26528 28690 26580
rect 9306 26500 9312 26512
rect 2746 26472 9312 26500
rect 9306 26460 9312 26472
rect 9364 26460 9370 26512
rect 11333 26503 11391 26509
rect 11333 26469 11345 26503
rect 11379 26469 11391 26503
rect 11333 26463 11391 26469
rect 1762 26364 1768 26376
rect 1723 26336 1768 26364
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 4157 26367 4215 26373
rect 4157 26333 4169 26367
rect 4203 26333 4215 26367
rect 5074 26364 5080 26376
rect 5035 26336 5080 26364
rect 4157 26327 4215 26333
rect 4172 26296 4200 26327
rect 5074 26324 5080 26336
rect 5132 26324 5138 26376
rect 10873 26367 10931 26373
rect 10873 26333 10885 26367
rect 10919 26364 10931 26367
rect 11348 26364 11376 26463
rect 15286 26460 15292 26512
rect 15344 26500 15350 26512
rect 15657 26503 15715 26509
rect 15657 26500 15669 26503
rect 15344 26472 15669 26500
rect 15344 26460 15350 26472
rect 15657 26469 15669 26472
rect 15703 26500 15715 26503
rect 16853 26503 16911 26509
rect 16853 26500 16865 26503
rect 15703 26472 16865 26500
rect 15703 26469 15715 26472
rect 15657 26463 15715 26469
rect 16853 26469 16865 26472
rect 16899 26469 16911 26503
rect 16853 26463 16911 26469
rect 18874 26460 18880 26512
rect 18932 26500 18938 26512
rect 23293 26503 23351 26509
rect 18932 26472 20116 26500
rect 18932 26460 18938 26472
rect 11532 26404 13400 26432
rect 11532 26373 11560 26404
rect 10919 26336 11376 26364
rect 11517 26367 11575 26373
rect 10919 26333 10931 26336
rect 10873 26327 10931 26333
rect 11517 26333 11529 26367
rect 11563 26333 11575 26367
rect 11974 26364 11980 26376
rect 11935 26336 11980 26364
rect 11517 26327 11575 26333
rect 11974 26324 11980 26336
rect 12032 26324 12038 26376
rect 12710 26364 12716 26376
rect 12671 26336 12716 26364
rect 12710 26324 12716 26336
rect 12768 26324 12774 26376
rect 13372 26373 13400 26404
rect 13814 26392 13820 26444
rect 13872 26432 13878 26444
rect 15197 26435 15255 26441
rect 15197 26432 15209 26435
rect 13872 26404 15209 26432
rect 13872 26392 13878 26404
rect 15197 26401 15209 26404
rect 15243 26401 15255 26435
rect 16666 26432 16672 26444
rect 16627 26404 16672 26432
rect 15197 26395 15255 26401
rect 16666 26392 16672 26404
rect 16724 26392 16730 26444
rect 18782 26432 18788 26444
rect 17696 26404 18788 26432
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26364 13415 26367
rect 14182 26364 14188 26376
rect 13403 26336 14188 26364
rect 13403 26333 13415 26336
rect 13357 26327 13415 26333
rect 14182 26324 14188 26336
rect 14240 26324 14246 26376
rect 14369 26367 14427 26373
rect 14369 26333 14381 26367
rect 14415 26364 14427 26367
rect 15013 26367 15071 26373
rect 15013 26364 15025 26367
rect 14415 26336 15025 26364
rect 14415 26333 14427 26336
rect 14369 26327 14427 26333
rect 15013 26333 15025 26336
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 15746 26324 15752 26376
rect 15804 26364 15810 26376
rect 16485 26367 16543 26373
rect 16485 26364 16497 26367
rect 15804 26336 16497 26364
rect 15804 26324 15810 26336
rect 16485 26333 16497 26336
rect 16531 26364 16543 26367
rect 17696 26364 17724 26404
rect 18782 26392 18788 26404
rect 18840 26392 18846 26444
rect 16531 26336 17724 26364
rect 18049 26367 18107 26373
rect 16531 26333 16543 26336
rect 16485 26327 16543 26333
rect 18049 26333 18061 26367
rect 18095 26333 18107 26367
rect 18049 26327 18107 26333
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26364 18751 26367
rect 18966 26364 18972 26376
rect 18739 26336 18972 26364
rect 18739 26333 18751 26336
rect 18693 26327 18751 26333
rect 4172 26268 12020 26296
rect 11992 26240 12020 26268
rect 12250 26256 12256 26308
rect 12308 26296 12314 26308
rect 12805 26299 12863 26305
rect 12805 26296 12817 26299
rect 12308 26268 12817 26296
rect 12308 26256 12314 26268
rect 12805 26265 12817 26268
rect 12851 26265 12863 26299
rect 18064 26296 18092 26327
rect 18966 26324 18972 26336
rect 19024 26324 19030 26376
rect 19426 26324 19432 26376
rect 19484 26364 19490 26376
rect 20088 26373 20116 26472
rect 23293 26469 23305 26503
rect 23339 26469 23351 26503
rect 23293 26463 23351 26469
rect 19613 26367 19671 26373
rect 19613 26364 19625 26367
rect 19484 26336 19625 26364
rect 19484 26324 19490 26336
rect 19613 26333 19625 26336
rect 19659 26364 19671 26367
rect 20073 26367 20131 26373
rect 19659 26336 19840 26364
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 19058 26296 19064 26308
rect 18064 26268 19064 26296
rect 12805 26259 12863 26265
rect 19058 26256 19064 26268
rect 19116 26256 19122 26308
rect 19812 26296 19840 26336
rect 20073 26333 20085 26367
rect 20119 26333 20131 26367
rect 20073 26327 20131 26333
rect 20162 26324 20168 26376
rect 20220 26364 20226 26376
rect 20901 26367 20959 26373
rect 20901 26364 20913 26367
rect 20220 26336 20913 26364
rect 20220 26324 20226 26336
rect 20901 26333 20913 26336
rect 20947 26333 20959 26367
rect 21542 26364 21548 26376
rect 21503 26336 21548 26364
rect 20901 26327 20959 26333
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 22189 26367 22247 26373
rect 22189 26333 22201 26367
rect 22235 26364 22247 26367
rect 22738 26364 22744 26376
rect 22235 26336 22744 26364
rect 22235 26333 22247 26336
rect 22189 26327 22247 26333
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26364 22891 26367
rect 23308 26364 23336 26463
rect 25866 26460 25872 26512
rect 25924 26500 25930 26512
rect 26053 26503 26111 26509
rect 26053 26500 26065 26503
rect 25924 26472 26065 26500
rect 25924 26460 25930 26472
rect 26053 26469 26065 26472
rect 26099 26469 26111 26503
rect 26053 26463 26111 26469
rect 25958 26392 25964 26444
rect 26016 26432 26022 26444
rect 26016 26404 28120 26432
rect 26016 26392 26022 26404
rect 22879 26336 23336 26364
rect 23477 26367 23535 26373
rect 22879 26333 22891 26336
rect 22833 26327 22891 26333
rect 23477 26333 23489 26367
rect 23523 26333 23535 26367
rect 23477 26327 23535 26333
rect 21450 26296 21456 26308
rect 19812 26268 21456 26296
rect 21450 26256 21456 26268
rect 21508 26256 21514 26308
rect 23492 26296 23520 26327
rect 23566 26324 23572 26376
rect 23624 26364 23630 26376
rect 25133 26367 25191 26373
rect 25133 26364 25145 26367
rect 23624 26336 25145 26364
rect 23624 26324 23630 26336
rect 25133 26333 25145 26336
rect 25179 26333 25191 26367
rect 26234 26364 26240 26376
rect 26195 26336 26240 26364
rect 25133 26327 25191 26333
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 26878 26364 26884 26376
rect 26839 26336 26884 26364
rect 26878 26324 26884 26336
rect 26936 26324 26942 26376
rect 27246 26324 27252 26376
rect 27304 26364 27310 26376
rect 28092 26373 28120 26404
rect 27525 26367 27583 26373
rect 27525 26364 27537 26367
rect 27304 26336 27537 26364
rect 27304 26324 27310 26336
rect 27525 26333 27537 26336
rect 27571 26333 27583 26367
rect 27525 26327 27583 26333
rect 28077 26367 28135 26373
rect 28077 26333 28089 26367
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 26510 26296 26516 26308
rect 23492 26268 26516 26296
rect 26510 26256 26516 26268
rect 26568 26256 26574 26308
rect 11974 26188 11980 26240
rect 12032 26188 12038 26240
rect 12069 26231 12127 26237
rect 12069 26197 12081 26231
rect 12115 26228 12127 26231
rect 12434 26228 12440 26240
rect 12115 26200 12440 26228
rect 12115 26197 12127 26200
rect 12069 26191 12127 26197
rect 12434 26188 12440 26200
rect 12492 26188 12498 26240
rect 13354 26188 13360 26240
rect 13412 26228 13418 26240
rect 13449 26231 13507 26237
rect 13449 26228 13461 26231
rect 13412 26200 13461 26228
rect 13412 26188 13418 26200
rect 13449 26197 13461 26200
rect 13495 26197 13507 26231
rect 18138 26228 18144 26240
rect 18099 26200 18144 26228
rect 13449 26191 13507 26197
rect 18138 26188 18144 26200
rect 18196 26188 18202 26240
rect 22005 26231 22063 26237
rect 22005 26197 22017 26231
rect 22051 26228 22063 26231
rect 22830 26228 22836 26240
rect 22051 26200 22836 26228
rect 22051 26197 22063 26200
rect 22005 26191 22063 26197
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 24946 26228 24952 26240
rect 24907 26200 24952 26228
rect 24946 26188 24952 26200
rect 25004 26188 25010 26240
rect 26694 26228 26700 26240
rect 26655 26200 26700 26228
rect 26694 26188 26700 26200
rect 26752 26188 26758 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 4985 26027 5043 26033
rect 4985 25993 4997 26027
rect 5031 26024 5043 26027
rect 5074 26024 5080 26036
rect 5031 25996 5080 26024
rect 5031 25993 5043 25996
rect 4985 25987 5043 25993
rect 5074 25984 5080 25996
rect 5132 25984 5138 26036
rect 13906 25984 13912 26036
rect 13964 26024 13970 26036
rect 15105 26027 15163 26033
rect 15105 26024 15117 26027
rect 13964 25996 15117 26024
rect 13964 25984 13970 25996
rect 15105 25993 15117 25996
rect 15151 25993 15163 26027
rect 27522 26024 27528 26036
rect 27483 25996 27528 26024
rect 15105 25987 15163 25993
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 11790 25956 11796 25968
rect 11751 25928 11796 25956
rect 11790 25916 11796 25928
rect 11848 25916 11854 25968
rect 11882 25916 11888 25968
rect 11940 25956 11946 25968
rect 13354 25956 13360 25968
rect 11940 25928 11985 25956
rect 13315 25928 13360 25956
rect 11940 25916 11946 25928
rect 13354 25916 13360 25928
rect 13412 25916 13418 25968
rect 19426 25956 19432 25968
rect 17880 25928 19432 25956
rect 4893 25891 4951 25897
rect 4893 25857 4905 25891
rect 4939 25857 4951 25891
rect 4893 25851 4951 25857
rect 4908 25820 4936 25851
rect 6454 25848 6460 25900
rect 6512 25888 6518 25900
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 6512 25860 8125 25888
rect 6512 25848 6518 25860
rect 8113 25857 8125 25860
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 9766 25848 9772 25900
rect 9824 25888 9830 25900
rect 10597 25891 10655 25897
rect 10597 25888 10609 25891
rect 9824 25860 10609 25888
rect 9824 25848 9830 25860
rect 10597 25857 10609 25860
rect 10643 25857 10655 25891
rect 14550 25888 14556 25900
rect 14511 25860 14556 25888
rect 10597 25851 10655 25857
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 15013 25891 15071 25897
rect 15013 25857 15025 25891
rect 15059 25888 15071 25891
rect 15286 25888 15292 25900
rect 15059 25860 15292 25888
rect 15059 25857 15071 25860
rect 15013 25851 15071 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25888 17095 25891
rect 17218 25888 17224 25900
rect 17083 25860 17224 25888
rect 17083 25857 17095 25860
rect 17037 25851 17095 25857
rect 17218 25848 17224 25860
rect 17276 25848 17282 25900
rect 17880 25897 17908 25928
rect 19426 25916 19432 25928
rect 19484 25916 19490 25968
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25857 17923 25891
rect 17865 25851 17923 25857
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25888 18567 25891
rect 19613 25891 19671 25897
rect 19613 25888 19625 25891
rect 18555 25860 19625 25888
rect 18555 25857 18567 25860
rect 18509 25851 18567 25857
rect 19613 25857 19625 25860
rect 19659 25857 19671 25891
rect 20990 25888 20996 25900
rect 20951 25860 20996 25888
rect 19613 25851 19671 25857
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 21082 25848 21088 25900
rect 21140 25888 21146 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21140 25860 22017 25888
rect 21140 25848 21146 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 24397 25891 24455 25897
rect 24397 25857 24409 25891
rect 24443 25888 24455 25891
rect 24946 25888 24952 25900
rect 24443 25860 24952 25888
rect 24443 25857 24455 25860
rect 24397 25851 24455 25857
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25888 25651 25891
rect 26694 25888 26700 25900
rect 25639 25860 26700 25888
rect 25639 25857 25651 25860
rect 25593 25851 25651 25857
rect 26694 25848 26700 25860
rect 26752 25848 26758 25900
rect 27706 25888 27712 25900
rect 27667 25860 27712 25888
rect 27706 25848 27712 25860
rect 27764 25848 27770 25900
rect 28353 25891 28411 25897
rect 28353 25857 28365 25891
rect 28399 25857 28411 25891
rect 28353 25851 28411 25857
rect 12069 25823 12127 25829
rect 12069 25820 12081 25823
rect 4908 25792 12081 25820
rect 12069 25789 12081 25792
rect 12115 25820 12127 25823
rect 13262 25820 13268 25832
rect 12115 25792 12434 25820
rect 13223 25792 13268 25820
rect 12115 25789 12127 25792
rect 12069 25783 12127 25789
rect 8205 25755 8263 25761
rect 8205 25721 8217 25755
rect 8251 25752 8263 25755
rect 12406 25752 12434 25792
rect 13262 25780 13268 25792
rect 13320 25780 13326 25832
rect 13541 25823 13599 25829
rect 13541 25789 13553 25823
rect 13587 25789 13599 25823
rect 13541 25783 13599 25789
rect 15657 25823 15715 25829
rect 15657 25789 15669 25823
rect 15703 25789 15715 25823
rect 15657 25783 15715 25789
rect 15841 25823 15899 25829
rect 15841 25789 15853 25823
rect 15887 25820 15899 25823
rect 18230 25820 18236 25832
rect 15887 25792 18236 25820
rect 15887 25789 15899 25792
rect 15841 25783 15899 25789
rect 13556 25752 13584 25783
rect 15672 25752 15700 25783
rect 18230 25780 18236 25792
rect 18288 25780 18294 25832
rect 18690 25820 18696 25832
rect 18651 25792 18696 25820
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 22646 25820 22652 25832
rect 22607 25792 22652 25820
rect 22646 25780 22652 25792
rect 22704 25780 22710 25832
rect 22833 25823 22891 25829
rect 22833 25789 22845 25823
rect 22879 25820 22891 25823
rect 24118 25820 24124 25832
rect 22879 25792 24124 25820
rect 22879 25789 22891 25792
rect 22833 25783 22891 25789
rect 24118 25780 24124 25792
rect 24176 25780 24182 25832
rect 27522 25780 27528 25832
rect 27580 25820 27586 25832
rect 28368 25820 28396 25851
rect 27580 25792 28396 25820
rect 27580 25780 27586 25792
rect 8251 25724 11376 25752
rect 12406 25724 13584 25752
rect 14016 25724 15700 25752
rect 16301 25755 16359 25761
rect 8251 25721 8263 25724
rect 8205 25715 8263 25721
rect 10413 25687 10471 25693
rect 10413 25653 10425 25687
rect 10459 25684 10471 25687
rect 11238 25684 11244 25696
rect 10459 25656 11244 25684
rect 10459 25653 10471 25656
rect 10413 25647 10471 25653
rect 11238 25644 11244 25656
rect 11296 25644 11302 25696
rect 11348 25684 11376 25724
rect 11882 25684 11888 25696
rect 11348 25656 11888 25684
rect 11882 25644 11888 25656
rect 11940 25684 11946 25696
rect 14016 25684 14044 25724
rect 16301 25721 16313 25755
rect 16347 25752 16359 25755
rect 21542 25752 21548 25764
rect 16347 25724 21548 25752
rect 16347 25721 16359 25724
rect 16301 25715 16359 25721
rect 11940 25656 14044 25684
rect 11940 25644 11946 25656
rect 14274 25644 14280 25696
rect 14332 25684 14338 25696
rect 14369 25687 14427 25693
rect 14369 25684 14381 25687
rect 14332 25656 14381 25684
rect 14332 25644 14338 25656
rect 14369 25653 14381 25656
rect 14415 25653 14427 25687
rect 14369 25647 14427 25653
rect 15102 25644 15108 25696
rect 15160 25684 15166 25696
rect 16316 25684 16344 25715
rect 21542 25712 21548 25724
rect 21600 25712 21606 25764
rect 23293 25755 23351 25761
rect 23293 25721 23305 25755
rect 23339 25752 23351 25755
rect 24762 25752 24768 25764
rect 23339 25724 24768 25752
rect 23339 25721 23351 25724
rect 23293 25715 23351 25721
rect 24762 25712 24768 25724
rect 24820 25712 24826 25764
rect 17126 25684 17132 25696
rect 15160 25656 16344 25684
rect 17087 25656 17132 25684
rect 15160 25644 15166 25656
rect 17126 25644 17132 25656
rect 17184 25644 17190 25696
rect 17954 25684 17960 25696
rect 17915 25656 17960 25684
rect 17954 25644 17960 25656
rect 18012 25644 18018 25696
rect 18874 25684 18880 25696
rect 18835 25656 18880 25684
rect 18874 25644 18880 25656
rect 18932 25644 18938 25696
rect 20809 25687 20867 25693
rect 20809 25653 20821 25687
rect 20855 25684 20867 25687
rect 21358 25684 21364 25696
rect 20855 25656 21364 25684
rect 20855 25653 20867 25656
rect 20809 25647 20867 25653
rect 21358 25644 21364 25656
rect 21416 25644 21422 25696
rect 22094 25644 22100 25696
rect 22152 25684 22158 25696
rect 22152 25656 22197 25684
rect 22152 25644 22158 25656
rect 23382 25644 23388 25696
rect 23440 25684 23446 25696
rect 24213 25687 24271 25693
rect 24213 25684 24225 25687
rect 23440 25656 24225 25684
rect 23440 25644 23446 25656
rect 24213 25653 24225 25656
rect 24259 25653 24271 25687
rect 25682 25684 25688 25696
rect 25643 25656 25688 25684
rect 24213 25647 24271 25653
rect 25682 25644 25688 25656
rect 25740 25644 25746 25696
rect 27338 25644 27344 25696
rect 27396 25684 27402 25696
rect 28169 25687 28227 25693
rect 28169 25684 28181 25687
rect 27396 25656 28181 25684
rect 27396 25644 27402 25656
rect 28169 25653 28181 25656
rect 28215 25653 28227 25687
rect 28169 25647 28227 25653
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 12253 25483 12311 25489
rect 12253 25449 12265 25483
rect 12299 25480 12311 25483
rect 13906 25480 13912 25492
rect 12299 25452 13912 25480
rect 12299 25449 12311 25452
rect 12253 25443 12311 25449
rect 13906 25440 13912 25452
rect 13964 25440 13970 25492
rect 14366 25480 14372 25492
rect 14327 25452 14372 25480
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 16850 25440 16856 25492
rect 16908 25480 16914 25492
rect 17589 25483 17647 25489
rect 17589 25480 17601 25483
rect 16908 25452 17601 25480
rect 16908 25440 16914 25452
rect 17589 25449 17601 25452
rect 17635 25449 17647 25483
rect 17589 25443 17647 25449
rect 18230 25440 18236 25492
rect 18288 25480 18294 25492
rect 19889 25483 19947 25489
rect 19889 25480 19901 25483
rect 18288 25452 19901 25480
rect 18288 25440 18294 25452
rect 19889 25449 19901 25452
rect 19935 25449 19947 25483
rect 21542 25480 21548 25492
rect 21503 25452 21548 25480
rect 19889 25443 19947 25449
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 25225 25483 25283 25489
rect 25225 25449 25237 25483
rect 25271 25480 25283 25483
rect 27430 25480 27436 25492
rect 25271 25452 27436 25480
rect 25271 25449 25283 25452
rect 25225 25443 25283 25449
rect 27430 25440 27436 25452
rect 27488 25440 27494 25492
rect 27890 25480 27896 25492
rect 27851 25452 27896 25480
rect 27890 25440 27896 25452
rect 27948 25440 27954 25492
rect 11701 25415 11759 25421
rect 11701 25381 11713 25415
rect 11747 25412 11759 25415
rect 13170 25412 13176 25424
rect 11747 25384 13176 25412
rect 11747 25381 11759 25384
rect 11701 25375 11759 25381
rect 13170 25372 13176 25384
rect 13228 25372 13234 25424
rect 13262 25372 13268 25424
rect 13320 25412 13326 25424
rect 17037 25415 17095 25421
rect 17037 25412 17049 25415
rect 13320 25384 17049 25412
rect 13320 25372 13326 25384
rect 17037 25381 17049 25384
rect 17083 25412 17095 25415
rect 25682 25412 25688 25424
rect 17083 25384 20576 25412
rect 17083 25381 17095 25384
rect 17037 25375 17095 25381
rect 17126 25344 17132 25356
rect 14568 25316 17132 25344
rect 11146 25276 11152 25288
rect 11107 25248 11152 25276
rect 11146 25236 11152 25248
rect 11204 25236 11210 25288
rect 11609 25279 11667 25285
rect 11609 25245 11621 25279
rect 11655 25276 11667 25279
rect 11698 25276 11704 25288
rect 11655 25248 11704 25276
rect 11655 25245 11667 25248
rect 11609 25239 11667 25245
rect 11698 25236 11704 25248
rect 11756 25236 11762 25288
rect 12437 25279 12495 25285
rect 12437 25245 12449 25279
rect 12483 25245 12495 25279
rect 13078 25276 13084 25288
rect 13039 25248 13084 25276
rect 12437 25239 12495 25245
rect 11054 25168 11060 25220
rect 11112 25208 11118 25220
rect 12452 25208 12480 25239
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25276 13599 25279
rect 13722 25276 13728 25288
rect 13587 25248 13728 25276
rect 13587 25245 13599 25248
rect 13541 25239 13599 25245
rect 13722 25236 13728 25248
rect 13780 25236 13786 25288
rect 14568 25285 14596 25316
rect 17126 25304 17132 25316
rect 17184 25304 17190 25356
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 16482 25276 16488 25288
rect 16443 25248 16488 25276
rect 14553 25239 14611 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 16669 25279 16727 25285
rect 16669 25245 16681 25279
rect 16715 25245 16727 25279
rect 16669 25239 16727 25245
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25276 17831 25279
rect 18138 25276 18144 25288
rect 17819 25248 18144 25276
rect 17819 25245 17831 25248
rect 17773 25239 17831 25245
rect 15102 25208 15108 25220
rect 11112 25180 12480 25208
rect 15063 25180 15108 25208
rect 11112 25168 11118 25180
rect 15102 25168 15108 25180
rect 15160 25168 15166 25220
rect 15197 25211 15255 25217
rect 15197 25177 15209 25211
rect 15243 25177 15255 25211
rect 15746 25208 15752 25220
rect 15707 25180 15752 25208
rect 15197 25171 15255 25177
rect 10318 25140 10324 25152
rect 10279 25112 10324 25140
rect 10318 25100 10324 25112
rect 10376 25100 10382 25152
rect 10965 25143 11023 25149
rect 10965 25109 10977 25143
rect 11011 25140 11023 25143
rect 11790 25140 11796 25152
rect 11011 25112 11796 25140
rect 11011 25109 11023 25112
rect 10965 25103 11023 25109
rect 11790 25100 11796 25112
rect 11848 25100 11854 25152
rect 12618 25100 12624 25152
rect 12676 25140 12682 25152
rect 12897 25143 12955 25149
rect 12897 25140 12909 25143
rect 12676 25112 12909 25140
rect 12676 25100 12682 25112
rect 12897 25109 12909 25112
rect 12943 25109 12955 25143
rect 12897 25103 12955 25109
rect 13633 25143 13691 25149
rect 13633 25109 13645 25143
rect 13679 25140 13691 25143
rect 14090 25140 14096 25152
rect 13679 25112 14096 25140
rect 13679 25109 13691 25112
rect 13633 25103 13691 25109
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 14366 25100 14372 25152
rect 14424 25140 14430 25152
rect 15212 25140 15240 25171
rect 15746 25168 15752 25180
rect 15804 25168 15810 25220
rect 16684 25208 16712 25239
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25276 18475 25279
rect 18966 25276 18972 25288
rect 18463 25248 18972 25276
rect 18463 25245 18475 25248
rect 18417 25239 18475 25245
rect 18966 25236 18972 25248
rect 19024 25236 19030 25288
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25276 19855 25279
rect 19978 25276 19984 25288
rect 19843 25248 19984 25276
rect 19843 25245 19855 25248
rect 19797 25239 19855 25245
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 20254 25236 20260 25288
rect 20312 25276 20318 25288
rect 20441 25279 20499 25285
rect 20441 25276 20453 25279
rect 20312 25248 20453 25276
rect 20312 25236 20318 25248
rect 20441 25245 20453 25248
rect 20487 25245 20499 25279
rect 20548 25276 20576 25384
rect 21192 25384 25688 25412
rect 21192 25353 21220 25384
rect 25682 25372 25688 25384
rect 25740 25372 25746 25424
rect 21177 25347 21235 25353
rect 21177 25313 21189 25347
rect 21223 25313 21235 25347
rect 21358 25344 21364 25356
rect 21319 25316 21364 25344
rect 21177 25307 21235 25313
rect 21358 25304 21364 25316
rect 21416 25304 21422 25356
rect 22833 25347 22891 25353
rect 22833 25313 22845 25347
rect 22879 25344 22891 25347
rect 23569 25347 23627 25353
rect 23569 25344 23581 25347
rect 22879 25316 23581 25344
rect 22879 25313 22891 25316
rect 22833 25307 22891 25313
rect 23569 25313 23581 25316
rect 23615 25313 23627 25347
rect 23569 25307 23627 25313
rect 23750 25304 23756 25356
rect 23808 25344 23814 25356
rect 26605 25347 26663 25353
rect 26605 25344 26617 25347
rect 23808 25316 26617 25344
rect 23808 25304 23814 25316
rect 26605 25313 26617 25316
rect 26651 25313 26663 25347
rect 26605 25307 26663 25313
rect 22738 25276 22744 25288
rect 20548 25248 22094 25276
rect 22699 25248 22744 25276
rect 20441 25239 20499 25245
rect 19242 25208 19248 25220
rect 16684 25180 19248 25208
rect 19242 25168 19248 25180
rect 19300 25168 19306 25220
rect 20533 25211 20591 25217
rect 20533 25177 20545 25211
rect 20579 25208 20591 25211
rect 22066 25208 22094 25248
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25276 23443 25279
rect 24486 25276 24492 25288
rect 23431 25248 24492 25276
rect 23431 25245 23443 25248
rect 23385 25239 23443 25245
rect 24486 25236 24492 25248
rect 24544 25236 24550 25288
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 25038 25276 25044 25288
rect 24811 25248 25044 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 25406 25276 25412 25288
rect 25367 25248 25412 25276
rect 25406 25236 25412 25248
rect 25464 25236 25470 25288
rect 25498 25236 25504 25288
rect 25556 25276 25562 25288
rect 25869 25279 25927 25285
rect 25869 25276 25881 25279
rect 25556 25248 25881 25276
rect 25556 25236 25562 25248
rect 25869 25245 25881 25248
rect 25915 25245 25927 25279
rect 25869 25239 25927 25245
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25276 26571 25279
rect 26786 25276 26792 25288
rect 26559 25248 26792 25276
rect 26559 25245 26571 25248
rect 26513 25239 26571 25245
rect 26786 25236 26792 25248
rect 26844 25236 26850 25288
rect 27798 25276 27804 25288
rect 27759 25248 27804 25276
rect 27798 25236 27804 25248
rect 27856 25236 27862 25288
rect 24029 25211 24087 25217
rect 24029 25208 24041 25211
rect 20579 25180 21956 25208
rect 22066 25180 24041 25208
rect 20579 25177 20591 25180
rect 20533 25171 20591 25177
rect 14424 25112 15240 25140
rect 18233 25143 18291 25149
rect 14424 25100 14430 25112
rect 18233 25109 18245 25143
rect 18279 25140 18291 25143
rect 20162 25140 20168 25152
rect 18279 25112 20168 25140
rect 18279 25109 18291 25112
rect 18233 25103 18291 25109
rect 20162 25100 20168 25112
rect 20220 25100 20226 25152
rect 21928 25140 21956 25180
rect 24029 25177 24041 25180
rect 24075 25177 24087 25211
rect 24029 25171 24087 25177
rect 25961 25211 26019 25217
rect 25961 25177 25973 25211
rect 26007 25208 26019 25211
rect 28166 25208 28172 25220
rect 26007 25180 28172 25208
rect 26007 25177 26019 25180
rect 25961 25171 26019 25177
rect 28166 25168 28172 25180
rect 28224 25168 28230 25220
rect 23198 25140 23204 25152
rect 21928 25112 23204 25140
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 24581 25143 24639 25149
rect 24581 25109 24593 25143
rect 24627 25140 24639 25143
rect 25130 25140 25136 25152
rect 24627 25112 25136 25140
rect 24627 25109 24639 25112
rect 24581 25103 24639 25109
rect 25130 25100 25136 25112
rect 25188 25100 25194 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 11974 24896 11980 24948
rect 12032 24936 12038 24948
rect 15746 24936 15752 24948
rect 12032 24908 15752 24936
rect 12032 24896 12038 24908
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 18141 24939 18199 24945
rect 18141 24905 18153 24939
rect 18187 24905 18199 24939
rect 18141 24899 18199 24905
rect 17129 24871 17187 24877
rect 17129 24868 17141 24871
rect 16868 24840 17141 24868
rect 1762 24800 1768 24812
rect 1723 24772 1768 24800
rect 1762 24760 1768 24772
rect 1820 24760 1826 24812
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 9217 24803 9275 24809
rect 9217 24800 9229 24803
rect 8444 24772 9229 24800
rect 8444 24760 8450 24772
rect 9217 24769 9229 24772
rect 9263 24769 9275 24803
rect 9858 24800 9864 24812
rect 9819 24772 9864 24800
rect 9217 24763 9275 24769
rect 9858 24760 9864 24772
rect 9916 24760 9922 24812
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24769 10563 24803
rect 10505 24763 10563 24769
rect 10520 24732 10548 24763
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 10744 24772 11713 24800
rect 10744 24760 10750 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 11790 24760 11796 24812
rect 11848 24800 11854 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 11848 24772 13001 24800
rect 11848 24760 11854 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13170 24760 13176 24812
rect 13228 24800 13234 24812
rect 13909 24803 13967 24809
rect 13909 24800 13921 24803
rect 13228 24772 13921 24800
rect 13228 24760 13234 24772
rect 13909 24769 13921 24772
rect 13955 24769 13967 24803
rect 14090 24800 14096 24812
rect 14051 24772 14096 24800
rect 13909 24763 13967 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 14550 24760 14556 24812
rect 14608 24800 14614 24812
rect 16868 24800 16896 24840
rect 17129 24837 17141 24840
rect 17175 24837 17187 24871
rect 18156 24868 18184 24899
rect 20898 24896 20904 24948
rect 20956 24936 20962 24948
rect 20956 24908 25176 24936
rect 20956 24896 20962 24908
rect 22738 24868 22744 24880
rect 18156 24840 18460 24868
rect 17129 24831 17187 24837
rect 14608 24772 16896 24800
rect 18325 24803 18383 24809
rect 14608 24760 14614 24772
rect 18325 24769 18337 24803
rect 18371 24769 18383 24803
rect 18432 24800 18460 24840
rect 22066 24840 22744 24868
rect 18969 24803 19027 24809
rect 18969 24800 18981 24803
rect 18432 24772 18981 24800
rect 18325 24763 18383 24769
rect 18969 24769 18981 24772
rect 19015 24769 19027 24803
rect 18969 24763 19027 24769
rect 19429 24803 19487 24809
rect 19429 24769 19441 24803
rect 19475 24800 19487 24803
rect 20162 24800 20168 24812
rect 19475 24772 20168 24800
rect 19475 24769 19487 24772
rect 19429 24763 19487 24769
rect 10870 24732 10876 24744
rect 10520 24704 10876 24732
rect 10870 24692 10876 24704
rect 10928 24692 10934 24744
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 12805 24735 12863 24741
rect 12805 24732 12817 24735
rect 11011 24704 12817 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 12805 24701 12817 24704
rect 12851 24701 12863 24735
rect 12805 24695 12863 24701
rect 16482 24692 16488 24744
rect 16540 24732 16546 24744
rect 17037 24735 17095 24741
rect 17037 24732 17049 24735
rect 16540 24704 17049 24732
rect 16540 24692 16546 24704
rect 17037 24701 17049 24704
rect 17083 24701 17095 24735
rect 18340 24732 18368 24763
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 20257 24803 20315 24809
rect 20257 24769 20269 24803
rect 20303 24769 20315 24803
rect 20257 24763 20315 24769
rect 20717 24803 20775 24809
rect 20717 24769 20729 24803
rect 20763 24800 20775 24803
rect 21082 24800 21088 24812
rect 20763 24772 21088 24800
rect 20763 24769 20775 24772
rect 20717 24763 20775 24769
rect 18782 24732 18788 24744
rect 18340 24704 18788 24732
rect 17037 24695 17095 24701
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 19794 24732 19800 24744
rect 19300 24704 19800 24732
rect 19300 24692 19306 24704
rect 19794 24692 19800 24704
rect 19852 24692 19858 24744
rect 20272 24732 20300 24763
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 22066 24800 22094 24840
rect 22738 24828 22744 24840
rect 22796 24868 22802 24880
rect 23934 24868 23940 24880
rect 22796 24840 23940 24868
rect 22796 24828 22802 24840
rect 23934 24828 23940 24840
rect 23992 24828 23998 24880
rect 21192 24772 22094 24800
rect 23569 24803 23627 24809
rect 21192 24732 21220 24772
rect 23569 24769 23581 24803
rect 23615 24800 23627 24803
rect 23842 24800 23848 24812
rect 23615 24772 23848 24800
rect 23615 24769 23627 24772
rect 23569 24763 23627 24769
rect 23842 24760 23848 24772
rect 23900 24760 23906 24812
rect 25148 24809 25176 24908
rect 25406 24868 25412 24880
rect 25367 24840 25412 24868
rect 25406 24828 25412 24840
rect 25464 24828 25470 24880
rect 25133 24803 25191 24809
rect 25133 24769 25145 24803
rect 25179 24769 25191 24803
rect 25866 24800 25872 24812
rect 25827 24772 25872 24800
rect 25133 24763 25191 24769
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 27249 24803 27307 24809
rect 27249 24769 27261 24803
rect 27295 24800 27307 24803
rect 27338 24800 27344 24812
rect 27295 24772 27344 24800
rect 27295 24769 27307 24772
rect 27249 24763 27307 24769
rect 27338 24760 27344 24772
rect 27396 24760 27402 24812
rect 28166 24800 28172 24812
rect 28127 24772 28172 24800
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 20272 24704 21220 24732
rect 21266 24692 21272 24744
rect 21324 24732 21330 24744
rect 22005 24735 22063 24741
rect 22005 24732 22017 24735
rect 21324 24704 22017 24732
rect 21324 24692 21330 24704
rect 22005 24701 22017 24704
rect 22051 24701 22063 24735
rect 22186 24732 22192 24744
rect 22147 24704 22192 24732
rect 22005 24695 22063 24701
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 23290 24732 23296 24744
rect 22572 24704 23296 24732
rect 9033 24667 9091 24673
rect 9033 24633 9045 24667
rect 9079 24664 9091 24667
rect 9766 24664 9772 24676
rect 9079 24636 9772 24664
rect 9079 24633 9091 24636
rect 9033 24627 9091 24633
rect 9766 24624 9772 24636
rect 9824 24624 9830 24676
rect 10321 24667 10379 24673
rect 10321 24633 10333 24667
rect 10367 24664 10379 24667
rect 11146 24664 11152 24676
rect 10367 24636 11152 24664
rect 10367 24633 10379 24636
rect 10321 24627 10379 24633
rect 11146 24624 11152 24636
rect 11204 24624 11210 24676
rect 17589 24667 17647 24673
rect 17589 24633 17601 24667
rect 17635 24664 17647 24667
rect 22572 24664 22600 24704
rect 23290 24692 23296 24704
rect 23348 24692 23354 24744
rect 23753 24735 23811 24741
rect 23753 24701 23765 24735
rect 23799 24732 23811 24735
rect 26050 24732 26056 24744
rect 23799 24704 26056 24732
rect 23799 24701 23811 24704
rect 23753 24695 23811 24701
rect 26050 24692 26056 24704
rect 26108 24692 26114 24744
rect 17635 24636 22600 24664
rect 22649 24667 22707 24673
rect 17635 24633 17647 24636
rect 17589 24627 17647 24633
rect 22649 24633 22661 24667
rect 22695 24664 22707 24667
rect 22922 24664 22928 24676
rect 22695 24636 22928 24664
rect 22695 24633 22707 24636
rect 22649 24627 22707 24633
rect 22922 24624 22928 24636
rect 22980 24664 22986 24676
rect 25498 24664 25504 24676
rect 22980 24636 25504 24664
rect 22980 24624 22986 24636
rect 25498 24624 25504 24636
rect 25556 24624 25562 24676
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 4062 24596 4068 24608
rect 1627 24568 4068 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 4062 24556 4068 24568
rect 4120 24556 4126 24608
rect 9677 24599 9735 24605
rect 9677 24565 9689 24599
rect 9723 24596 9735 24599
rect 11054 24596 11060 24608
rect 9723 24568 11060 24596
rect 9723 24565 9735 24568
rect 9677 24559 9735 24565
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 11793 24599 11851 24605
rect 11793 24565 11805 24599
rect 11839 24596 11851 24599
rect 12986 24596 12992 24608
rect 11839 24568 12992 24596
rect 11839 24565 11851 24568
rect 11793 24559 11851 24565
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 13449 24599 13507 24605
rect 13449 24565 13461 24599
rect 13495 24596 13507 24599
rect 14277 24599 14335 24605
rect 14277 24596 14289 24599
rect 13495 24568 14289 24596
rect 13495 24565 13507 24568
rect 13449 24559 13507 24565
rect 14277 24565 14289 24568
rect 14323 24596 14335 24599
rect 14642 24596 14648 24608
rect 14323 24568 14648 24596
rect 14323 24565 14335 24568
rect 14277 24559 14335 24565
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 18785 24599 18843 24605
rect 18785 24565 18797 24599
rect 18831 24596 18843 24599
rect 19334 24596 19340 24608
rect 18831 24568 19340 24596
rect 18831 24565 18843 24568
rect 18785 24559 18843 24565
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 19518 24596 19524 24608
rect 19479 24568 19524 24596
rect 19518 24556 19524 24568
rect 19576 24556 19582 24608
rect 20070 24596 20076 24608
rect 20031 24568 20076 24596
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20806 24596 20812 24608
rect 20767 24568 20812 24596
rect 20806 24556 20812 24568
rect 20864 24556 20870 24608
rect 22554 24556 22560 24608
rect 22612 24596 22618 24608
rect 23937 24599 23995 24605
rect 23937 24596 23949 24599
rect 22612 24568 23949 24596
rect 22612 24556 22618 24568
rect 23937 24565 23949 24568
rect 23983 24596 23995 24599
rect 24578 24596 24584 24608
rect 23983 24568 24584 24596
rect 23983 24565 23995 24568
rect 23937 24559 23995 24565
rect 24578 24556 24584 24568
rect 24636 24556 24642 24608
rect 25958 24596 25964 24608
rect 25919 24568 25964 24596
rect 25958 24556 25964 24568
rect 26016 24556 26022 24608
rect 26050 24556 26056 24608
rect 26108 24596 26114 24608
rect 27341 24599 27399 24605
rect 27341 24596 27353 24599
rect 26108 24568 27353 24596
rect 26108 24556 26114 24568
rect 27341 24565 27353 24568
rect 27387 24565 27399 24599
rect 27341 24559 27399 24565
rect 27985 24599 28043 24605
rect 27985 24565 27997 24599
rect 28031 24596 28043 24599
rect 28534 24596 28540 24608
rect 28031 24568 28540 24596
rect 28031 24565 28043 24568
rect 27985 24559 28043 24565
rect 28534 24556 28540 24568
rect 28592 24556 28598 24608
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 12161 24395 12219 24401
rect 12161 24361 12173 24395
rect 12207 24392 12219 24395
rect 13078 24392 13084 24404
rect 12207 24364 13084 24392
rect 12207 24361 12219 24364
rect 12161 24355 12219 24361
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 13633 24395 13691 24401
rect 13633 24361 13645 24395
rect 13679 24392 13691 24395
rect 14366 24392 14372 24404
rect 13679 24364 14372 24392
rect 13679 24361 13691 24364
rect 13633 24355 13691 24361
rect 14366 24352 14372 24364
rect 14424 24352 14430 24404
rect 17678 24352 17684 24404
rect 17736 24392 17742 24404
rect 20165 24395 20223 24401
rect 17736 24364 19288 24392
rect 17736 24352 17742 24364
rect 9858 24284 9864 24336
rect 9916 24324 9922 24336
rect 15381 24327 15439 24333
rect 9916 24296 12848 24324
rect 9916 24284 9922 24296
rect 8481 24259 8539 24265
rect 8481 24225 8493 24259
rect 8527 24256 8539 24259
rect 9401 24259 9459 24265
rect 9401 24256 9413 24259
rect 8527 24228 9413 24256
rect 8527 24225 8539 24228
rect 8481 24219 8539 24225
rect 9401 24225 9413 24228
rect 9447 24225 9459 24259
rect 9401 24219 9459 24225
rect 10318 24216 10324 24268
rect 10376 24256 10382 24268
rect 10965 24259 11023 24265
rect 10965 24256 10977 24259
rect 10376 24228 10977 24256
rect 10376 24216 10382 24228
rect 10965 24225 10977 24228
rect 11011 24225 11023 24259
rect 10965 24219 11023 24225
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 11974 24256 11980 24268
rect 11655 24228 11980 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 11974 24216 11980 24228
rect 12032 24216 12038 24268
rect 12360 24228 12664 24256
rect 8386 24188 8392 24200
rect 8347 24160 8392 24188
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 9214 24188 9220 24200
rect 9175 24160 9220 24188
rect 9214 24148 9220 24160
rect 9272 24148 9278 24200
rect 12360 24197 12388 24228
rect 12345 24191 12403 24197
rect 12345 24157 12357 24191
rect 12391 24157 12403 24191
rect 12345 24151 12403 24157
rect 11057 24123 11115 24129
rect 11057 24089 11069 24123
rect 11103 24089 11115 24123
rect 12636 24120 12664 24228
rect 12820 24200 12848 24296
rect 15381 24293 15393 24327
rect 15427 24324 15439 24327
rect 16298 24324 16304 24336
rect 15427 24296 16304 24324
rect 15427 24293 15439 24296
rect 15381 24287 15439 24293
rect 16298 24284 16304 24296
rect 16356 24284 16362 24336
rect 16853 24327 16911 24333
rect 16853 24293 16865 24327
rect 16899 24324 16911 24327
rect 19150 24324 19156 24336
rect 16899 24296 19156 24324
rect 16899 24293 16911 24296
rect 16853 24287 16911 24293
rect 19150 24284 19156 24296
rect 19208 24284 19214 24336
rect 19260 24324 19288 24364
rect 20165 24361 20177 24395
rect 20211 24392 20223 24395
rect 20990 24392 20996 24404
rect 20211 24364 20996 24392
rect 20211 24361 20223 24364
rect 20165 24355 20223 24361
rect 20990 24352 20996 24364
rect 21048 24352 21054 24404
rect 22186 24352 22192 24404
rect 22244 24392 22250 24404
rect 23569 24395 23627 24401
rect 23569 24392 23581 24395
rect 22244 24364 23581 24392
rect 22244 24352 22250 24364
rect 23569 24361 23581 24364
rect 23615 24361 23627 24395
rect 23569 24355 23627 24361
rect 24762 24352 24768 24404
rect 24820 24392 24826 24404
rect 24949 24395 25007 24401
rect 24949 24392 24961 24395
rect 24820 24364 24961 24392
rect 24820 24352 24826 24364
rect 24949 24361 24961 24364
rect 24995 24361 25007 24395
rect 27246 24392 27252 24404
rect 27207 24364 27252 24392
rect 24949 24355 25007 24361
rect 19610 24324 19616 24336
rect 19260 24296 19616 24324
rect 19610 24284 19616 24296
rect 19668 24284 19674 24336
rect 19794 24284 19800 24336
rect 19852 24324 19858 24336
rect 21453 24327 21511 24333
rect 21453 24324 21465 24327
rect 19852 24296 21465 24324
rect 19852 24284 19858 24296
rect 21453 24293 21465 24296
rect 21499 24293 21511 24327
rect 22922 24324 22928 24336
rect 22883 24296 22928 24324
rect 21453 24287 21511 24293
rect 22922 24284 22928 24296
rect 22980 24284 22986 24336
rect 23106 24284 23112 24336
rect 23164 24324 23170 24336
rect 24964 24324 24992 24355
rect 27246 24352 27252 24364
rect 27304 24352 27310 24404
rect 27706 24352 27712 24404
rect 27764 24392 27770 24404
rect 27893 24395 27951 24401
rect 27893 24392 27905 24395
rect 27764 24364 27905 24392
rect 27764 24352 27770 24364
rect 27893 24361 27905 24364
rect 27939 24361 27951 24395
rect 27893 24355 27951 24361
rect 23164 24296 24716 24324
rect 24964 24296 27200 24324
rect 23164 24284 23170 24296
rect 17405 24259 17463 24265
rect 17405 24225 17417 24259
rect 17451 24256 17463 24259
rect 19702 24256 19708 24268
rect 17451 24228 19708 24256
rect 17451 24225 17463 24228
rect 17405 24219 17463 24225
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 20070 24216 20076 24268
rect 20128 24256 20134 24268
rect 22557 24259 22615 24265
rect 20128 24228 21680 24256
rect 20128 24216 20134 24228
rect 12802 24188 12808 24200
rect 12763 24160 12808 24188
rect 12802 24148 12808 24160
rect 12860 24148 12866 24200
rect 13170 24148 13176 24200
rect 13228 24188 13234 24200
rect 13541 24191 13599 24197
rect 13541 24188 13553 24191
rect 13228 24160 13553 24188
rect 13228 24148 13234 24160
rect 13541 24157 13553 24160
rect 13587 24157 13599 24191
rect 13541 24151 13599 24157
rect 14921 24191 14979 24197
rect 14921 24157 14933 24191
rect 14967 24188 14979 24191
rect 15286 24188 15292 24200
rect 14967 24160 15292 24188
rect 14967 24157 14979 24160
rect 14921 24151 14979 24157
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24157 15623 24191
rect 16114 24188 16120 24200
rect 16075 24160 16120 24188
rect 15565 24151 15623 24157
rect 13188 24120 13216 24148
rect 15580 24120 15608 24151
rect 16114 24148 16120 24160
rect 16172 24148 16178 24200
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24157 16819 24191
rect 16761 24151 16819 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24188 17647 24191
rect 18138 24188 18144 24200
rect 17635 24160 18144 24188
rect 17635 24157 17647 24160
rect 17589 24151 17647 24157
rect 11057 24083 11115 24089
rect 12084 24092 12434 24120
rect 12636 24092 13216 24120
rect 14752 24092 15608 24120
rect 9861 24055 9919 24061
rect 9861 24021 9873 24055
rect 9907 24052 9919 24055
rect 10594 24052 10600 24064
rect 9907 24024 10600 24052
rect 9907 24021 9919 24024
rect 9861 24015 9919 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 11072 24052 11100 24083
rect 12084 24052 12112 24092
rect 11072 24024 12112 24052
rect 12406 24052 12434 24092
rect 12618 24052 12624 24064
rect 12406 24024 12624 24052
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 12894 24052 12900 24064
rect 12855 24024 12900 24052
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 14752 24061 14780 24092
rect 14737 24055 14795 24061
rect 14737 24021 14749 24055
rect 14783 24021 14795 24055
rect 14737 24015 14795 24021
rect 15194 24012 15200 24064
rect 15252 24052 15258 24064
rect 16209 24055 16267 24061
rect 16209 24052 16221 24055
rect 15252 24024 16221 24052
rect 15252 24012 15258 24024
rect 16209 24021 16221 24024
rect 16255 24021 16267 24055
rect 16776 24052 16804 24151
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 18782 24188 18788 24200
rect 18647 24160 18788 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 18782 24148 18788 24160
rect 18840 24148 18846 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19610 24188 19616 24200
rect 19475 24160 19616 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19610 24148 19616 24160
rect 19668 24148 19674 24200
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20349 24191 20407 24197
rect 20349 24188 20361 24191
rect 20036 24160 20361 24188
rect 20036 24148 20042 24160
rect 20349 24157 20361 24160
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24188 20867 24191
rect 21450 24188 21456 24200
rect 20855 24160 21456 24188
rect 20855 24157 20867 24160
rect 20809 24151 20867 24157
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 21652 24197 21680 24228
rect 22557 24225 22569 24259
rect 22603 24256 22615 24259
rect 23382 24256 23388 24268
rect 22603 24228 23388 24256
rect 22603 24225 22615 24228
rect 22557 24219 22615 24225
rect 23382 24216 23388 24228
rect 23440 24216 23446 24268
rect 24578 24256 24584 24268
rect 24539 24228 24584 24256
rect 24578 24216 24584 24228
rect 24636 24216 24642 24268
rect 24688 24256 24716 24296
rect 26050 24256 26056 24268
rect 24688 24228 25820 24256
rect 26011 24228 26056 24256
rect 21637 24191 21695 24197
rect 21637 24157 21649 24191
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 22373 24191 22431 24197
rect 22373 24157 22385 24191
rect 22419 24188 22431 24191
rect 23106 24188 23112 24200
rect 22419 24160 23112 24188
rect 22419 24157 22431 24160
rect 22373 24151 22431 24157
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23566 24188 23572 24200
rect 23523 24160 23572 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 23566 24148 23572 24160
rect 23624 24188 23630 24200
rect 23842 24188 23848 24200
rect 23624 24160 23848 24188
rect 23624 24148 23630 24160
rect 23842 24148 23848 24160
rect 23900 24148 23906 24200
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24188 24823 24191
rect 25682 24188 25688 24200
rect 24811 24160 25688 24188
rect 24811 24157 24823 24160
rect 24765 24151 24823 24157
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 18049 24123 18107 24129
rect 18049 24089 18061 24123
rect 18095 24120 18107 24123
rect 19521 24123 19579 24129
rect 18095 24092 19288 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18598 24052 18604 24064
rect 16776 24024 18604 24052
rect 16209 24015 16267 24021
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24052 18751 24055
rect 19150 24052 19156 24064
rect 18739 24024 19156 24052
rect 18739 24021 18751 24024
rect 18693 24015 18751 24021
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 19260 24052 19288 24092
rect 19521 24089 19533 24123
rect 19567 24120 19579 24123
rect 25498 24120 25504 24132
rect 19567 24092 25504 24120
rect 19567 24089 19579 24092
rect 19521 24083 19579 24089
rect 25498 24080 25504 24092
rect 25556 24080 25562 24132
rect 25792 24120 25820 24228
rect 26050 24216 26056 24228
rect 26108 24216 26114 24268
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24188 26295 24191
rect 26418 24188 26424 24200
rect 26283 24160 26424 24188
rect 26283 24157 26295 24160
rect 26237 24151 26295 24157
rect 26418 24148 26424 24160
rect 26476 24148 26482 24200
rect 27172 24197 27200 24296
rect 27157 24191 27215 24197
rect 27157 24157 27169 24191
rect 27203 24157 27215 24191
rect 27157 24151 27215 24157
rect 27801 24191 27859 24197
rect 27801 24157 27813 24191
rect 27847 24157 27859 24191
rect 27801 24151 27859 24157
rect 26697 24123 26755 24129
rect 26697 24120 26709 24123
rect 25792 24092 26709 24120
rect 26697 24089 26709 24092
rect 26743 24089 26755 24123
rect 26697 24083 26755 24089
rect 19610 24052 19616 24064
rect 19260 24024 19616 24052
rect 19610 24012 19616 24024
rect 19668 24012 19674 24064
rect 20438 24012 20444 24064
rect 20496 24052 20502 24064
rect 20901 24055 20959 24061
rect 20901 24052 20913 24055
rect 20496 24024 20913 24052
rect 20496 24012 20502 24024
rect 20901 24021 20913 24024
rect 20947 24021 20959 24055
rect 20901 24015 20959 24021
rect 22186 24012 22192 24064
rect 22244 24052 22250 24064
rect 25222 24052 25228 24064
rect 22244 24024 25228 24052
rect 22244 24012 22250 24024
rect 25222 24012 25228 24024
rect 25280 24012 25286 24064
rect 25314 24012 25320 24064
rect 25372 24052 25378 24064
rect 27816 24052 27844 24151
rect 25372 24024 27844 24052
rect 25372 24012 25378 24024
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 8021 23851 8079 23857
rect 8021 23817 8033 23851
rect 8067 23817 8079 23851
rect 8021 23811 8079 23817
rect 8036 23780 8064 23811
rect 9214 23808 9220 23860
rect 9272 23848 9278 23860
rect 9493 23851 9551 23857
rect 9493 23848 9505 23851
rect 9272 23820 9505 23848
rect 9272 23808 9278 23820
rect 9493 23817 9505 23820
rect 9539 23817 9551 23851
rect 9493 23811 9551 23817
rect 11164 23820 19288 23848
rect 8036 23752 8892 23780
rect 1762 23712 1768 23724
rect 1723 23684 1768 23712
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 8864 23721 8892 23752
rect 8205 23715 8263 23721
rect 8205 23681 8217 23715
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 8849 23715 8907 23721
rect 8849 23681 8861 23715
rect 8895 23681 8907 23715
rect 9306 23712 9312 23724
rect 9267 23684 9312 23712
rect 8849 23675 8907 23681
rect 8220 23644 8248 23675
rect 9306 23672 9312 23684
rect 9364 23672 9370 23724
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23712 10379 23715
rect 11054 23712 11060 23724
rect 10367 23684 11060 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 11164 23721 11192 23820
rect 12636 23721 12664 23820
rect 14737 23783 14795 23789
rect 14737 23780 14749 23783
rect 13740 23752 14749 23780
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 12161 23715 12219 23721
rect 12161 23681 12173 23715
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 8386 23644 8392 23656
rect 8220 23616 8392 23644
rect 8386 23604 8392 23616
rect 8444 23644 8450 23656
rect 12176 23644 12204 23675
rect 12894 23672 12900 23724
rect 12952 23712 12958 23724
rect 13633 23715 13691 23721
rect 13633 23712 13645 23715
rect 12952 23684 13645 23712
rect 12952 23672 12958 23684
rect 13633 23681 13645 23684
rect 13679 23681 13691 23715
rect 13633 23675 13691 23681
rect 8444 23616 10824 23644
rect 8444 23604 8450 23616
rect 1581 23579 1639 23585
rect 1581 23545 1593 23579
rect 1627 23576 1639 23579
rect 10686 23576 10692 23588
rect 1627 23548 10692 23576
rect 1627 23545 1639 23548
rect 1581 23539 1639 23545
rect 10686 23536 10692 23548
rect 10744 23536 10750 23588
rect 8665 23511 8723 23517
rect 8665 23477 8677 23511
rect 8711 23508 8723 23511
rect 10410 23508 10416 23520
rect 8711 23480 10416 23508
rect 8711 23477 8723 23480
rect 8665 23471 8723 23477
rect 10410 23468 10416 23480
rect 10468 23468 10474 23520
rect 10796 23508 10824 23616
rect 10980 23616 12204 23644
rect 10980 23585 11008 23616
rect 12986 23604 12992 23656
rect 13044 23644 13050 23656
rect 13449 23647 13507 23653
rect 13449 23644 13461 23647
rect 13044 23616 13461 23644
rect 13044 23604 13050 23616
rect 13449 23613 13461 23616
rect 13495 23613 13507 23647
rect 13449 23607 13507 23613
rect 10965 23579 11023 23585
rect 10965 23545 10977 23579
rect 11011 23545 11023 23579
rect 10965 23539 11023 23545
rect 11977 23579 12035 23585
rect 11977 23545 11989 23579
rect 12023 23576 12035 23579
rect 13740 23576 13768 23752
rect 14737 23749 14749 23752
rect 14783 23749 14795 23783
rect 14737 23743 14795 23749
rect 15289 23783 15347 23789
rect 15289 23749 15301 23783
rect 15335 23780 15347 23783
rect 15930 23780 15936 23792
rect 15335 23752 15936 23780
rect 15335 23749 15347 23752
rect 15289 23743 15347 23749
rect 15930 23740 15936 23752
rect 15988 23740 15994 23792
rect 18509 23783 18567 23789
rect 18509 23749 18521 23783
rect 18555 23780 18567 23783
rect 18874 23780 18880 23792
rect 18555 23752 18880 23780
rect 18555 23749 18567 23752
rect 18509 23743 18567 23749
rect 18874 23740 18880 23752
rect 18932 23740 18938 23792
rect 19150 23780 19156 23792
rect 19111 23752 19156 23780
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 19260 23780 19288 23820
rect 19702 23808 19708 23860
rect 19760 23848 19766 23860
rect 22646 23848 22652 23860
rect 19760 23820 22652 23848
rect 19760 23808 19766 23820
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 24118 23808 24124 23860
rect 24176 23848 24182 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 24176 23820 25145 23848
rect 24176 23808 24182 23820
rect 25133 23817 25145 23820
rect 25179 23817 25191 23851
rect 25682 23848 25688 23860
rect 25643 23820 25688 23848
rect 25133 23811 25191 23817
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 22462 23780 22468 23792
rect 19260 23752 22468 23780
rect 22462 23740 22468 23752
rect 22520 23740 22526 23792
rect 23290 23780 23296 23792
rect 23251 23752 23296 23780
rect 23290 23740 23296 23752
rect 23348 23740 23354 23792
rect 23385 23783 23443 23789
rect 23385 23749 23397 23783
rect 23431 23780 23443 23783
rect 24670 23780 24676 23792
rect 23431 23752 24676 23780
rect 23431 23749 23443 23752
rect 23385 23743 23443 23749
rect 24670 23740 24676 23752
rect 24728 23740 24734 23792
rect 25590 23780 25596 23792
rect 24872 23752 25596 23780
rect 15470 23672 15476 23724
rect 15528 23712 15534 23724
rect 15841 23715 15899 23721
rect 15841 23712 15853 23715
rect 15528 23684 15853 23712
rect 15528 23672 15534 23684
rect 15841 23681 15853 23684
rect 15887 23712 15899 23715
rect 16942 23712 16948 23724
rect 15887 23684 16948 23712
rect 15887 23681 15899 23684
rect 15841 23675 15899 23681
rect 16942 23672 16948 23684
rect 17000 23672 17006 23724
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 17678 23712 17684 23724
rect 17083 23684 17684 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 17678 23672 17684 23684
rect 17736 23672 17742 23724
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 18049 23715 18107 23721
rect 18049 23712 18061 23715
rect 18012 23684 18061 23712
rect 18012 23672 18018 23684
rect 18049 23681 18061 23684
rect 18095 23681 18107 23715
rect 20162 23712 20168 23724
rect 20123 23684 20168 23712
rect 18049 23675 18107 23681
rect 20162 23672 20168 23684
rect 20220 23672 20226 23724
rect 20809 23715 20867 23721
rect 20809 23681 20821 23715
rect 20855 23712 20867 23715
rect 21082 23712 21088 23724
rect 20855 23684 21088 23712
rect 20855 23681 20867 23684
rect 20809 23675 20867 23681
rect 21082 23672 21088 23684
rect 21140 23672 21146 23724
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 24872 23712 24900 23752
rect 25590 23740 25596 23752
rect 25648 23740 25654 23792
rect 25038 23712 25044 23724
rect 24443 23684 24900 23712
rect 24999 23684 25044 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 14642 23644 14648 23656
rect 14603 23616 14648 23644
rect 14642 23604 14648 23616
rect 14700 23604 14706 23656
rect 15378 23644 15384 23656
rect 15120 23616 15384 23644
rect 15120 23576 15148 23616
rect 15378 23604 15384 23616
rect 15436 23604 15442 23656
rect 16117 23647 16175 23653
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 16206 23644 16212 23656
rect 16163 23616 16212 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23613 17923 23647
rect 17865 23607 17923 23613
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23644 19119 23647
rect 19426 23644 19432 23656
rect 19107 23616 19432 23644
rect 19107 23613 19119 23616
rect 19061 23607 19119 23613
rect 17880 23576 17908 23607
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 19518 23604 19524 23656
rect 19576 23644 19582 23656
rect 19702 23644 19708 23656
rect 19576 23616 19708 23644
rect 19576 23604 19582 23616
rect 19702 23604 19708 23616
rect 19760 23604 19766 23656
rect 20530 23644 20536 23656
rect 19812 23616 20536 23644
rect 12023 23548 13768 23576
rect 14016 23548 15148 23576
rect 15304 23548 17908 23576
rect 12023 23545 12035 23548
rect 11977 23539 12035 23545
rect 11790 23508 11796 23520
rect 10796 23480 11796 23508
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 12713 23511 12771 23517
rect 12713 23477 12725 23511
rect 12759 23508 12771 23511
rect 14016 23508 14044 23548
rect 12759 23480 14044 23508
rect 14093 23511 14151 23517
rect 12759 23477 12771 23480
rect 12713 23471 12771 23477
rect 14093 23477 14105 23511
rect 14139 23508 14151 23511
rect 14918 23508 14924 23520
rect 14139 23480 14924 23508
rect 14139 23477 14151 23480
rect 14093 23471 14151 23477
rect 14918 23468 14924 23480
rect 14976 23508 14982 23520
rect 15304 23508 15332 23548
rect 18782 23536 18788 23588
rect 18840 23576 18846 23588
rect 19812 23576 19840 23616
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 22186 23644 22192 23656
rect 20947 23616 22192 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 22186 23604 22192 23616
rect 22244 23604 22250 23656
rect 22296 23644 22324 23675
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 25130 23672 25136 23724
rect 25188 23712 25194 23724
rect 25869 23715 25927 23721
rect 25869 23712 25881 23715
rect 25188 23684 25881 23712
rect 25188 23672 25194 23684
rect 25869 23681 25881 23684
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 26050 23672 26056 23724
rect 26108 23712 26114 23724
rect 26513 23715 26571 23721
rect 26513 23712 26525 23715
rect 26108 23684 26525 23712
rect 26108 23672 26114 23684
rect 26513 23681 26525 23684
rect 26559 23681 26571 23715
rect 28350 23712 28356 23724
rect 28311 23684 28356 23712
rect 26513 23675 26571 23681
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 24946 23644 24952 23656
rect 22296 23616 24952 23644
rect 24946 23604 24952 23616
rect 25004 23604 25010 23656
rect 18840 23548 19840 23576
rect 20257 23579 20315 23585
rect 18840 23536 18846 23548
rect 20257 23545 20269 23579
rect 20303 23576 20315 23579
rect 23474 23576 23480 23588
rect 20303 23548 23480 23576
rect 20303 23545 20315 23548
rect 20257 23539 20315 23545
rect 23474 23536 23480 23548
rect 23532 23536 23538 23588
rect 23845 23579 23903 23585
rect 23845 23545 23857 23579
rect 23891 23576 23903 23579
rect 24026 23576 24032 23588
rect 23891 23548 24032 23576
rect 23891 23545 23903 23548
rect 23845 23539 23903 23545
rect 24026 23536 24032 23548
rect 24084 23576 24090 23588
rect 27798 23576 27804 23588
rect 24084 23548 27804 23576
rect 24084 23536 24090 23548
rect 27798 23536 27804 23548
rect 27856 23536 27862 23588
rect 14976 23480 15332 23508
rect 16853 23511 16911 23517
rect 14976 23468 14982 23480
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 17494 23508 17500 23520
rect 16899 23480 17500 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 17770 23468 17776 23520
rect 17828 23508 17834 23520
rect 21266 23508 21272 23520
rect 17828 23480 21272 23508
rect 17828 23468 17834 23480
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 21358 23468 21364 23520
rect 21416 23508 21422 23520
rect 22373 23511 22431 23517
rect 22373 23508 22385 23511
rect 21416 23480 22385 23508
rect 21416 23468 21422 23480
rect 22373 23477 22385 23480
rect 22419 23477 22431 23511
rect 22373 23471 22431 23477
rect 22922 23468 22928 23520
rect 22980 23508 22986 23520
rect 24489 23511 24547 23517
rect 24489 23508 24501 23511
rect 22980 23480 24501 23508
rect 22980 23468 22986 23480
rect 24489 23477 24501 23480
rect 24535 23477 24547 23511
rect 24489 23471 24547 23477
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 26329 23511 26387 23517
rect 26329 23508 26341 23511
rect 26292 23480 26341 23508
rect 26292 23468 26298 23480
rect 26329 23477 26341 23480
rect 26375 23477 26387 23511
rect 26329 23471 26387 23477
rect 26602 23468 26608 23520
rect 26660 23508 26666 23520
rect 28169 23511 28227 23517
rect 28169 23508 28181 23511
rect 26660 23480 28181 23508
rect 26660 23468 26666 23480
rect 28169 23477 28181 23480
rect 28215 23477 28227 23511
rect 28169 23471 28227 23477
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 10594 23304 10600 23316
rect 10555 23276 10600 23304
rect 10594 23264 10600 23276
rect 10652 23304 10658 23316
rect 13998 23304 14004 23316
rect 10652 23276 14004 23304
rect 10652 23264 10658 23276
rect 13998 23264 14004 23276
rect 14056 23264 14062 23316
rect 14918 23304 14924 23316
rect 14879 23276 14924 23304
rect 14918 23264 14924 23276
rect 14976 23264 14982 23316
rect 18138 23264 18144 23316
rect 18196 23304 18202 23316
rect 18693 23307 18751 23313
rect 18693 23304 18705 23307
rect 18196 23276 18705 23304
rect 18196 23264 18202 23276
rect 18693 23273 18705 23276
rect 18739 23273 18751 23307
rect 19886 23304 19892 23316
rect 18693 23267 18751 23273
rect 18800 23276 19892 23304
rect 10410 23168 10416 23180
rect 10371 23140 10416 23168
rect 10410 23128 10416 23140
rect 10468 23128 10474 23180
rect 11054 23128 11060 23180
rect 11112 23168 11118 23180
rect 11333 23171 11391 23177
rect 11333 23168 11345 23171
rect 11112 23140 11345 23168
rect 11112 23128 11118 23140
rect 11333 23137 11345 23140
rect 11379 23137 11391 23171
rect 12434 23168 12440 23180
rect 12395 23140 12440 23168
rect 11333 23131 11391 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 12621 23171 12679 23177
rect 12621 23137 12633 23171
rect 12667 23137 12679 23171
rect 12621 23131 12679 23137
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 9585 23103 9643 23109
rect 9585 23100 9597 23103
rect 8352 23072 9597 23100
rect 8352 23060 8358 23072
rect 9585 23069 9597 23072
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 9677 22967 9735 22973
rect 9677 22933 9689 22967
rect 9723 22964 9735 22967
rect 10244 22964 10272 23063
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 11296 23072 11529 23100
rect 11296 23060 11302 23072
rect 11517 23069 11529 23072
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 11882 23060 11888 23112
rect 11940 23100 11946 23112
rect 12636 23100 12664 23131
rect 13906 23128 13912 23180
rect 13964 23168 13970 23180
rect 14461 23171 14519 23177
rect 14461 23168 14473 23171
rect 13964 23140 14473 23168
rect 13964 23128 13970 23140
rect 14461 23137 14473 23140
rect 14507 23137 14519 23171
rect 14461 23131 14519 23137
rect 15286 23128 15292 23180
rect 15344 23168 15350 23180
rect 18800 23168 18828 23276
rect 19886 23264 19892 23276
rect 19944 23264 19950 23316
rect 21266 23304 21272 23316
rect 21008 23276 21272 23304
rect 21008 23168 21036 23276
rect 21266 23264 21272 23276
rect 21324 23264 21330 23316
rect 24670 23304 24676 23316
rect 24631 23276 24676 23304
rect 24670 23264 24676 23276
rect 24728 23264 24734 23316
rect 26418 23304 26424 23316
rect 26379 23276 26424 23304
rect 26418 23264 26424 23276
rect 26476 23264 26482 23316
rect 15344 23140 18828 23168
rect 19306 23140 21036 23168
rect 15344 23128 15350 23140
rect 11940 23096 12388 23100
rect 12452 23096 12664 23100
rect 11940 23072 12664 23096
rect 13725 23103 13783 23109
rect 11940 23060 11946 23072
rect 12360 23068 12480 23072
rect 13725 23069 13737 23103
rect 13771 23100 13783 23103
rect 13814 23100 13820 23112
rect 13771 23072 13820 23100
rect 13771 23069 13783 23072
rect 13725 23063 13783 23069
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14366 23100 14372 23112
rect 14323 23072 14372 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 15396 23109 15424 23140
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23069 15439 23103
rect 17494 23100 17500 23112
rect 17455 23072 17500 23100
rect 15381 23063 15439 23069
rect 17494 23060 17500 23072
rect 17552 23060 17558 23112
rect 17678 23060 17684 23112
rect 17736 23100 17742 23112
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17736 23072 18153 23100
rect 17736 23060 17742 23072
rect 18141 23069 18153 23072
rect 18187 23100 18199 23103
rect 18601 23103 18659 23109
rect 18601 23100 18613 23103
rect 18187 23072 18613 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18601 23069 18613 23072
rect 18647 23100 18659 23103
rect 19150 23100 19156 23112
rect 18647 23072 19156 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 19150 23060 19156 23072
rect 19208 23060 19214 23112
rect 11977 23035 12035 23041
rect 11977 23001 11989 23035
rect 12023 23032 12035 23035
rect 13081 23035 13139 23041
rect 13081 23032 13093 23035
rect 12023 23004 13093 23032
rect 12023 23001 12035 23004
rect 11977 22995 12035 23001
rect 13081 23001 13093 23004
rect 13127 23032 13139 23035
rect 16209 23035 16267 23041
rect 16209 23032 16221 23035
rect 13127 23004 16221 23032
rect 13127 23001 13139 23004
rect 13081 22995 13139 23001
rect 16209 23001 16221 23004
rect 16255 23001 16267 23035
rect 16209 22995 16267 23001
rect 16298 22992 16304 23044
rect 16356 23032 16362 23044
rect 16850 23032 16856 23044
rect 16356 23004 16401 23032
rect 16811 23004 16856 23032
rect 16356 22992 16362 23004
rect 16850 22992 16856 23004
rect 16908 22992 16914 23044
rect 19306 23032 19334 23140
rect 21082 23128 21088 23180
rect 21140 23168 21146 23180
rect 21450 23168 21456 23180
rect 21140 23140 21456 23168
rect 21140 23128 21146 23140
rect 21450 23128 21456 23140
rect 21508 23168 21514 23180
rect 22649 23171 22707 23177
rect 21508 23140 21956 23168
rect 21508 23128 21514 23140
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 21174 23100 21180 23112
rect 20671 23072 21180 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21266 23060 21272 23112
rect 21324 23100 21330 23112
rect 21634 23100 21640 23112
rect 21324 23072 21640 23100
rect 21324 23060 21330 23072
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 21928 23109 21956 23140
rect 22649 23137 22661 23171
rect 22695 23168 22707 23171
rect 24946 23168 24952 23180
rect 22695 23140 24952 23168
rect 22695 23137 22707 23140
rect 22649 23131 22707 23137
rect 24946 23128 24952 23140
rect 25004 23128 25010 23180
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23069 21971 23103
rect 23750 23100 23756 23112
rect 21913 23063 21971 23069
rect 23492 23072 23756 23100
rect 19518 23032 19524 23044
rect 17236 23004 19334 23032
rect 19479 23004 19524 23032
rect 12066 22964 12072 22976
rect 9723 22936 12072 22964
rect 9723 22933 9735 22936
rect 9677 22927 9735 22933
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 13541 22967 13599 22973
rect 13541 22933 13553 22967
rect 13587 22964 13599 22967
rect 14734 22964 14740 22976
rect 13587 22936 14740 22964
rect 13587 22933 13599 22936
rect 13541 22927 13599 22933
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 15473 22967 15531 22973
rect 15473 22933 15485 22967
rect 15519 22964 15531 22967
rect 15746 22964 15752 22976
rect 15519 22936 15752 22964
rect 15519 22933 15531 22936
rect 15473 22927 15531 22933
rect 15746 22924 15752 22936
rect 15804 22924 15810 22976
rect 16482 22924 16488 22976
rect 16540 22964 16546 22976
rect 17236 22964 17264 23004
rect 19518 22992 19524 23004
rect 19576 22992 19582 23044
rect 19613 23035 19671 23041
rect 19613 23001 19625 23035
rect 19659 23001 19671 23035
rect 19613 22995 19671 23001
rect 16540 22936 17264 22964
rect 17313 22967 17371 22973
rect 16540 22924 16546 22936
rect 17313 22933 17325 22967
rect 17359 22964 17371 22967
rect 17862 22964 17868 22976
rect 17359 22936 17868 22964
rect 17359 22933 17371 22936
rect 17313 22927 17371 22933
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 17957 22967 18015 22973
rect 17957 22933 17969 22967
rect 18003 22964 18015 22967
rect 18874 22964 18880 22976
rect 18003 22936 18880 22964
rect 18003 22933 18015 22936
rect 17957 22927 18015 22933
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19628 22964 19656 22995
rect 19794 22992 19800 23044
rect 19852 23032 19858 23044
rect 20165 23035 20223 23041
rect 20165 23032 20177 23035
rect 19852 23004 20177 23032
rect 19852 22992 19858 23004
rect 20165 23001 20177 23004
rect 20211 23001 20223 23035
rect 20165 22995 20223 23001
rect 20717 23035 20775 23041
rect 20717 23001 20729 23035
rect 20763 23032 20775 23035
rect 21082 23032 21088 23044
rect 20763 23004 21088 23032
rect 20763 23001 20775 23004
rect 20717 22995 20775 23001
rect 21082 22992 21088 23004
rect 21140 22992 21146 23044
rect 22741 23035 22799 23041
rect 22741 23001 22753 23035
rect 22787 23032 22799 23035
rect 23492 23032 23520 23072
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 24486 23060 24492 23112
rect 24544 23100 24550 23112
rect 24581 23103 24639 23109
rect 24581 23100 24593 23103
rect 24544 23072 24593 23100
rect 24544 23060 24550 23072
rect 24581 23069 24593 23072
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 25869 23103 25927 23109
rect 25869 23069 25881 23103
rect 25915 23100 25927 23103
rect 26234 23100 26240 23112
rect 25915 23072 26240 23100
rect 25915 23069 25927 23072
rect 25869 23063 25927 23069
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 26329 23103 26387 23109
rect 26329 23069 26341 23103
rect 26375 23069 26387 23103
rect 26329 23063 26387 23069
rect 27985 23103 28043 23109
rect 27985 23069 27997 23103
rect 28031 23100 28043 23103
rect 28442 23100 28448 23112
rect 28031 23072 28448 23100
rect 28031 23069 28043 23072
rect 27985 23063 28043 23069
rect 23658 23032 23664 23044
rect 22787 23004 23520 23032
rect 23619 23004 23664 23032
rect 22787 23001 22799 23004
rect 22741 22995 22799 23001
rect 23658 22992 23664 23004
rect 23716 22992 23722 23044
rect 26344 23032 26372 23063
rect 28442 23060 28448 23072
rect 28500 23060 28506 23112
rect 25884 23004 26372 23032
rect 25884 22976 25912 23004
rect 19392 22936 19656 22964
rect 19392 22924 19398 22936
rect 20806 22924 20812 22976
rect 20864 22964 20870 22976
rect 21361 22967 21419 22973
rect 21361 22964 21373 22967
rect 20864 22936 21373 22964
rect 20864 22924 20870 22936
rect 21361 22933 21373 22936
rect 21407 22933 21419 22967
rect 21361 22927 21419 22933
rect 22005 22967 22063 22973
rect 22005 22933 22017 22967
rect 22051 22964 22063 22967
rect 23290 22964 23296 22976
rect 22051 22936 23296 22964
rect 22051 22933 22063 22936
rect 22005 22927 22063 22933
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 25682 22964 25688 22976
rect 25643 22936 25688 22964
rect 25682 22924 25688 22936
rect 25740 22924 25746 22976
rect 25866 22924 25872 22976
rect 25924 22924 25930 22976
rect 27798 22924 27804 22976
rect 27856 22964 27862 22976
rect 28077 22967 28135 22973
rect 28077 22964 28089 22967
rect 27856 22936 28089 22964
rect 27856 22924 27862 22936
rect 28077 22933 28089 22936
rect 28123 22933 28135 22967
rect 28077 22927 28135 22933
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 11882 22760 11888 22772
rect 11843 22732 11888 22760
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 18690 22760 18696 22772
rect 13372 22732 18696 22760
rect 1854 22652 1860 22704
rect 1912 22692 1918 22704
rect 13372 22701 13400 22732
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 19337 22763 19395 22769
rect 19337 22729 19349 22763
rect 19383 22760 19395 22763
rect 19426 22760 19432 22772
rect 19383 22732 19432 22760
rect 19383 22729 19395 22732
rect 19337 22723 19395 22729
rect 19426 22720 19432 22732
rect 19484 22760 19490 22772
rect 19794 22760 19800 22772
rect 19484 22732 19800 22760
rect 19484 22720 19490 22732
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 19886 22720 19892 22772
rect 19944 22760 19950 22772
rect 25682 22760 25688 22772
rect 19944 22732 23060 22760
rect 19944 22720 19950 22732
rect 13357 22695 13415 22701
rect 1912 22664 13124 22692
rect 1912 22652 1918 22664
rect 13096 22636 13124 22664
rect 13357 22661 13369 22695
rect 13403 22661 13415 22695
rect 15470 22692 15476 22704
rect 13357 22655 13415 22661
rect 13648 22664 15476 22692
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22593 8447 22627
rect 8389 22587 8447 22593
rect 9033 22627 9091 22633
rect 9033 22593 9045 22627
rect 9079 22624 9091 22627
rect 9677 22627 9735 22633
rect 9079 22596 9536 22624
rect 9079 22593 9091 22596
rect 9033 22587 9091 22593
rect 8404 22556 8432 22587
rect 9122 22556 9128 22568
rect 8404 22528 9128 22556
rect 9122 22516 9128 22528
rect 9180 22516 9186 22568
rect 9508 22497 9536 22596
rect 9677 22593 9689 22627
rect 9723 22593 9735 22627
rect 9677 22587 9735 22593
rect 9692 22556 9720 22587
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 10321 22627 10379 22633
rect 10321 22624 10333 22627
rect 9824 22596 10333 22624
rect 9824 22584 9830 22596
rect 10321 22593 10333 22596
rect 10367 22593 10379 22627
rect 10321 22587 10379 22593
rect 10962 22584 10968 22636
rect 11020 22624 11026 22636
rect 11149 22627 11207 22633
rect 11149 22624 11161 22627
rect 11020 22596 11161 22624
rect 11020 22584 11026 22596
rect 11149 22593 11161 22596
rect 11195 22593 11207 22627
rect 11790 22624 11796 22636
rect 11703 22596 11796 22624
rect 11149 22587 11207 22593
rect 11790 22584 11796 22596
rect 11848 22624 11854 22636
rect 12342 22624 12348 22636
rect 11848 22596 12348 22624
rect 11848 22584 11854 22596
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 13078 22624 13084 22636
rect 12991 22596 13084 22624
rect 13078 22584 13084 22596
rect 13136 22624 13142 22636
rect 13648 22624 13676 22664
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 15746 22692 15752 22704
rect 15707 22664 15752 22692
rect 15746 22652 15752 22664
rect 15804 22652 15810 22704
rect 16301 22695 16359 22701
rect 16301 22661 16313 22695
rect 16347 22692 16359 22695
rect 16850 22692 16856 22704
rect 16347 22664 16856 22692
rect 16347 22661 16359 22664
rect 16301 22655 16359 22661
rect 16850 22652 16856 22664
rect 16908 22692 16914 22704
rect 22738 22692 22744 22704
rect 16908 22664 22744 22692
rect 16908 22652 16914 22664
rect 22738 22652 22744 22664
rect 22796 22652 22802 22704
rect 13136 22596 13676 22624
rect 13136 22584 13142 22596
rect 13722 22584 13728 22636
rect 13780 22624 13786 22636
rect 14185 22627 14243 22633
rect 14185 22624 14197 22627
rect 13780 22596 14197 22624
rect 13780 22584 13786 22596
rect 14185 22593 14197 22596
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 14734 22584 14740 22636
rect 14792 22624 14798 22636
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14792 22596 15025 22624
rect 14792 22584 14798 22596
rect 15013 22593 15025 22596
rect 15059 22593 15071 22627
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 15013 22587 15071 22593
rect 17034 22584 17040 22596
rect 17092 22584 17098 22636
rect 17494 22624 17500 22636
rect 17455 22596 17500 22624
rect 17494 22584 17500 22596
rect 17552 22584 17558 22636
rect 17862 22584 17868 22636
rect 17920 22624 17926 22636
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 17920 22596 19993 22624
rect 17920 22584 17926 22596
rect 19981 22593 19993 22596
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 20901 22627 20959 22633
rect 20901 22593 20913 22627
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 11054 22556 11060 22568
rect 9692 22528 11060 22556
rect 11054 22516 11060 22528
rect 11112 22516 11118 22568
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22556 12495 22559
rect 12526 22556 12532 22568
rect 12483 22528 12532 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 12526 22516 12532 22528
rect 12584 22516 12590 22568
rect 13998 22516 14004 22568
rect 14056 22556 14062 22568
rect 15657 22559 15715 22565
rect 15657 22556 15669 22559
rect 14056 22528 15669 22556
rect 14056 22516 14062 22528
rect 15657 22525 15669 22528
rect 15703 22525 15715 22559
rect 18693 22559 18751 22565
rect 18693 22556 18705 22559
rect 15657 22519 15715 22525
rect 15764 22528 18705 22556
rect 9493 22491 9551 22497
rect 9493 22457 9505 22491
rect 9539 22457 9551 22491
rect 9493 22451 9551 22457
rect 10413 22491 10471 22497
rect 10413 22457 10425 22491
rect 10459 22488 10471 22491
rect 11698 22488 11704 22500
rect 10459 22460 11704 22488
rect 10459 22457 10471 22460
rect 10413 22451 10471 22457
rect 11698 22448 11704 22460
rect 11756 22448 11762 22500
rect 13630 22448 13636 22500
rect 13688 22488 13694 22500
rect 14366 22488 14372 22500
rect 13688 22460 14372 22488
rect 13688 22448 13694 22460
rect 14366 22448 14372 22460
rect 14424 22488 14430 22500
rect 15764 22488 15792 22528
rect 18693 22525 18705 22528
rect 18739 22556 18751 22559
rect 18782 22556 18788 22568
rect 18739 22528 18788 22556
rect 18739 22525 18751 22528
rect 18693 22519 18751 22525
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 18877 22559 18935 22565
rect 18877 22525 18889 22559
rect 18923 22556 18935 22559
rect 19426 22556 19432 22568
rect 18923 22528 19432 22556
rect 18923 22525 18935 22528
rect 18877 22519 18935 22525
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22556 19855 22559
rect 20254 22556 20260 22568
rect 19843 22528 20260 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 20254 22516 20260 22528
rect 20312 22516 20318 22568
rect 20916 22556 20944 22587
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21048 22596 22017 22624
rect 21048 22584 21054 22596
rect 22005 22593 22017 22596
rect 22051 22624 22063 22627
rect 22554 22624 22560 22636
rect 22051 22596 22560 22624
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 22922 22624 22928 22636
rect 22883 22596 22928 22624
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 21266 22556 21272 22568
rect 20916 22528 21272 22556
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 23032 22556 23060 22732
rect 23124 22732 25688 22760
rect 23124 22633 23152 22732
rect 25682 22720 25688 22732
rect 25740 22720 25746 22772
rect 23842 22652 23848 22704
rect 23900 22692 23906 22704
rect 24305 22695 24363 22701
rect 24305 22692 24317 22695
rect 23900 22664 24317 22692
rect 23900 22652 23906 22664
rect 24305 22661 24317 22664
rect 24351 22661 24363 22695
rect 25590 22692 25596 22704
rect 25530 22664 25596 22692
rect 24305 22655 24363 22661
rect 25590 22652 25596 22664
rect 25648 22652 25654 22704
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23109 22587 23167 22593
rect 23952 22596 24041 22624
rect 23566 22556 23572 22568
rect 23032 22528 23572 22556
rect 23566 22516 23572 22528
rect 23624 22516 23630 22568
rect 14424 22460 15792 22488
rect 17589 22491 17647 22497
rect 14424 22448 14430 22460
rect 17589 22457 17601 22491
rect 17635 22488 17647 22491
rect 19886 22488 19892 22500
rect 17635 22460 19892 22488
rect 17635 22457 17647 22460
rect 17589 22451 17647 22457
rect 19886 22448 19892 22460
rect 19944 22448 19950 22500
rect 20070 22448 20076 22500
rect 20128 22488 20134 22500
rect 21174 22488 21180 22500
rect 20128 22460 21180 22488
rect 20128 22448 20134 22460
rect 21174 22448 21180 22460
rect 21232 22448 21238 22500
rect 8205 22423 8263 22429
rect 8205 22389 8217 22423
rect 8251 22420 8263 22423
rect 8754 22420 8760 22432
rect 8251 22392 8760 22420
rect 8251 22389 8263 22392
rect 8205 22383 8263 22389
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 8849 22423 8907 22429
rect 8849 22389 8861 22423
rect 8895 22420 8907 22423
rect 10318 22420 10324 22432
rect 8895 22392 10324 22420
rect 8895 22389 8907 22392
rect 8849 22383 8907 22389
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 10502 22380 10508 22432
rect 10560 22420 10566 22432
rect 10965 22423 11023 22429
rect 10965 22420 10977 22423
rect 10560 22392 10977 22420
rect 10560 22380 10566 22392
rect 10965 22389 10977 22392
rect 11011 22389 11023 22423
rect 14274 22420 14280 22432
rect 14235 22392 14280 22420
rect 10965 22383 11023 22389
rect 14274 22380 14280 22392
rect 14332 22380 14338 22432
rect 14734 22380 14740 22432
rect 14792 22420 14798 22432
rect 14829 22423 14887 22429
rect 14829 22420 14841 22423
rect 14792 22392 14841 22420
rect 14792 22380 14798 22392
rect 14829 22389 14841 22392
rect 14875 22389 14887 22423
rect 14829 22383 14887 22389
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 16816 22392 16865 22420
rect 16816 22380 16822 22392
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 16853 22383 16911 22389
rect 18874 22380 18880 22432
rect 18932 22420 18938 22432
rect 19518 22420 19524 22432
rect 18932 22392 19524 22420
rect 18932 22380 18938 22392
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 19610 22380 19616 22432
rect 19668 22420 19674 22432
rect 20165 22423 20223 22429
rect 20165 22420 20177 22423
rect 19668 22392 20177 22420
rect 19668 22380 19674 22392
rect 20165 22389 20177 22392
rect 20211 22389 20223 22423
rect 20165 22383 20223 22389
rect 20898 22380 20904 22432
rect 20956 22420 20962 22432
rect 20993 22423 21051 22429
rect 20993 22420 21005 22423
rect 20956 22392 21005 22420
rect 20956 22380 20962 22392
rect 20993 22389 21005 22392
rect 21039 22389 21051 22423
rect 20993 22383 21051 22389
rect 22097 22423 22155 22429
rect 22097 22389 22109 22423
rect 22143 22420 22155 22423
rect 22186 22420 22192 22432
rect 22143 22392 22192 22420
rect 22143 22389 22155 22392
rect 22097 22383 22155 22389
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 22738 22380 22744 22432
rect 22796 22420 22802 22432
rect 23293 22423 23351 22429
rect 23293 22420 23305 22423
rect 22796 22392 23305 22420
rect 22796 22380 22802 22392
rect 23293 22389 23305 22392
rect 23339 22389 23351 22423
rect 23952 22420 23980 22596
rect 24029 22593 24041 22596
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 27890 22584 27896 22636
rect 27948 22624 27954 22636
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 27948 22596 28089 22624
rect 27948 22584 27954 22596
rect 28077 22593 28089 22596
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 28258 22488 28264 22500
rect 28219 22460 28264 22488
rect 28258 22448 28264 22460
rect 28316 22448 28322 22500
rect 24670 22420 24676 22432
rect 23952 22392 24676 22420
rect 23293 22383 23351 22389
rect 24670 22380 24676 22392
rect 24728 22380 24734 22432
rect 25682 22380 25688 22432
rect 25740 22420 25746 22432
rect 25777 22423 25835 22429
rect 25777 22420 25789 22423
rect 25740 22392 25789 22420
rect 25740 22380 25746 22392
rect 25777 22389 25789 22392
rect 25823 22389 25835 22423
rect 25777 22383 25835 22389
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 10870 22176 10876 22228
rect 10928 22216 10934 22228
rect 13722 22216 13728 22228
rect 10928 22188 13728 22216
rect 10928 22176 10934 22188
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 14182 22176 14188 22228
rect 14240 22216 14246 22228
rect 18782 22216 18788 22228
rect 14240 22188 18788 22216
rect 14240 22176 14246 22188
rect 18782 22176 18788 22188
rect 18840 22176 18846 22228
rect 18874 22176 18880 22228
rect 18932 22216 18938 22228
rect 19150 22216 19156 22228
rect 18932 22188 19156 22216
rect 18932 22176 18938 22188
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 19426 22216 19432 22228
rect 19387 22188 19432 22216
rect 19426 22176 19432 22188
rect 19484 22176 19490 22228
rect 19886 22176 19892 22228
rect 19944 22216 19950 22228
rect 19944 22188 23520 22216
rect 19944 22176 19950 22188
rect 9122 22108 9128 22160
rect 9180 22148 9186 22160
rect 13814 22148 13820 22160
rect 9180 22120 13820 22148
rect 9180 22108 9186 22120
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 15194 22148 15200 22160
rect 14660 22120 15200 22148
rect 10318 22040 10324 22092
rect 10376 22080 10382 22092
rect 11057 22083 11115 22089
rect 11057 22080 11069 22083
rect 10376 22052 11069 22080
rect 10376 22040 10382 22052
rect 11057 22049 11069 22052
rect 11103 22049 11115 22083
rect 11057 22043 11115 22049
rect 13265 22083 13323 22089
rect 13265 22049 13277 22083
rect 13311 22080 13323 22083
rect 14274 22080 14280 22092
rect 13311 22052 14280 22080
rect 13311 22049 13323 22052
rect 13265 22043 13323 22049
rect 14274 22040 14280 22052
rect 14332 22040 14338 22092
rect 1762 22012 1768 22024
rect 1723 21984 1768 22012
rect 1762 21972 1768 21984
rect 1820 21972 1826 22024
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 8812 21984 9505 22012
rect 8812 21972 8818 21984
rect 9493 21981 9505 21984
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 10502 22012 10508 22024
rect 10459 21984 10508 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 10873 22015 10931 22021
rect 10873 21981 10885 22015
rect 10919 21981 10931 22015
rect 10873 21975 10931 21981
rect 7374 21904 7380 21956
rect 7432 21944 7438 21956
rect 10888 21944 10916 21975
rect 11238 21972 11244 22024
rect 11296 22012 11302 22024
rect 11974 22012 11980 22024
rect 11296 21984 11980 22012
rect 11296 21972 11302 21984
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12158 22012 12164 22024
rect 12119 21984 12164 22012
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 13081 22015 13139 22021
rect 13081 22012 13093 22015
rect 12492 21984 13093 22012
rect 12492 21972 12498 21984
rect 13081 21981 13093 21984
rect 13127 22012 13139 22015
rect 14660 22012 14688 22120
rect 15194 22108 15200 22120
rect 15252 22108 15258 22160
rect 16850 22108 16856 22160
rect 16908 22148 16914 22160
rect 17037 22151 17095 22157
rect 17037 22148 17049 22151
rect 16908 22120 17049 22148
rect 16908 22108 16914 22120
rect 17037 22117 17049 22120
rect 17083 22148 17095 22151
rect 20070 22148 20076 22160
rect 17083 22120 20076 22148
rect 17083 22117 17095 22120
rect 17037 22111 17095 22117
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 20254 22108 20260 22160
rect 20312 22148 20318 22160
rect 20714 22148 20720 22160
rect 20312 22120 20720 22148
rect 20312 22108 20318 22120
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 21174 22108 21180 22160
rect 21232 22148 21238 22160
rect 22738 22148 22744 22160
rect 21232 22120 22744 22148
rect 21232 22108 21238 22120
rect 22738 22108 22744 22120
rect 22796 22108 22802 22160
rect 23492 22148 23520 22188
rect 23566 22176 23572 22228
rect 23624 22216 23630 22228
rect 24394 22216 24400 22228
rect 23624 22188 24400 22216
rect 23624 22176 23630 22188
rect 24394 22176 24400 22188
rect 24452 22176 24458 22228
rect 27614 22216 27620 22228
rect 24504 22188 27620 22216
rect 24504 22148 24532 22188
rect 27614 22176 27620 22188
rect 27672 22176 27678 22228
rect 23032 22120 23428 22148
rect 23492 22120 24532 22148
rect 15010 22040 15016 22092
rect 15068 22080 15074 22092
rect 15289 22083 15347 22089
rect 15289 22080 15301 22083
rect 15068 22052 15301 22080
rect 15068 22040 15074 22052
rect 15289 22049 15301 22052
rect 15335 22049 15347 22083
rect 15930 22080 15936 22092
rect 15891 22052 15936 22080
rect 15289 22043 15347 22049
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 16577 22083 16635 22089
rect 16577 22049 16589 22083
rect 16623 22080 16635 22083
rect 18046 22080 18052 22092
rect 16623 22052 18052 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 20990 22080 20996 22092
rect 18279 22052 20996 22080
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 22922 22080 22928 22092
rect 22883 22052 22928 22080
rect 22922 22040 22928 22052
rect 22980 22040 22986 22092
rect 13127 21984 14688 22012
rect 14745 22015 14803 22021
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 14745 21981 14757 22015
rect 14791 22012 14803 22015
rect 14791 21984 15148 22012
rect 14791 21981 14803 21984
rect 14745 21975 14803 21981
rect 7432 21916 10916 21944
rect 7432 21904 7438 21916
rect 11146 21904 11152 21956
rect 11204 21944 11210 21956
rect 14366 21944 14372 21956
rect 11204 21916 14372 21944
rect 11204 21904 11210 21916
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 15010 21944 15016 21956
rect 14476 21916 15016 21944
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 8754 21876 8760 21888
rect 1627 21848 8760 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 10042 21876 10048 21888
rect 9355 21848 10048 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10229 21879 10287 21885
rect 10229 21845 10241 21879
rect 10275 21876 10287 21879
rect 11054 21876 11060 21888
rect 10275 21848 11060 21876
rect 10275 21845 10287 21848
rect 10229 21839 10287 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11517 21879 11575 21885
rect 11517 21845 11529 21879
rect 11563 21876 11575 21879
rect 12618 21876 12624 21888
rect 11563 21848 12624 21876
rect 11563 21845 11575 21848
rect 11517 21839 11575 21845
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 13722 21876 13728 21888
rect 13683 21848 13728 21876
rect 13722 21836 13728 21848
rect 13780 21876 13786 21888
rect 14476 21876 14504 21916
rect 15010 21904 15016 21916
rect 15068 21904 15074 21956
rect 13780 21848 14504 21876
rect 14553 21879 14611 21885
rect 13780 21836 13786 21848
rect 14553 21845 14565 21879
rect 14599 21876 14611 21879
rect 14642 21876 14648 21888
rect 14599 21848 14648 21876
rect 14599 21845 14611 21848
rect 14553 21839 14611 21845
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 15120 21876 15148 21984
rect 16022 21972 16028 22024
rect 16080 22012 16086 22024
rect 16393 22015 16451 22021
rect 16393 22012 16405 22015
rect 16080 21984 16405 22012
rect 16080 21972 16086 21984
rect 16393 21981 16405 21984
rect 16439 21981 16451 22015
rect 18690 22012 18696 22024
rect 18651 21984 18696 22012
rect 16393 21975 16451 21981
rect 18690 21972 18696 21984
rect 18748 21972 18754 22024
rect 19518 21972 19524 22024
rect 19576 22012 19582 22024
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 19576 21984 19625 22012
rect 19576 21972 19582 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 22554 21972 22560 22024
rect 22612 22012 22618 22024
rect 22833 22015 22891 22021
rect 22833 22012 22845 22015
rect 22612 21984 22845 22012
rect 22612 21972 22618 21984
rect 22833 21981 22845 21984
rect 22879 22012 22891 22015
rect 23032 22012 23060 22120
rect 23400 22080 23428 22120
rect 23400 22052 25268 22080
rect 22879 21984 23060 22012
rect 23477 22015 23535 22021
rect 22879 21981 22891 21984
rect 22833 21975 22891 21981
rect 23477 21981 23489 22015
rect 23523 22012 23535 22015
rect 23523 21984 23612 22012
rect 23523 21981 23535 21984
rect 23477 21975 23535 21981
rect 15378 21904 15384 21956
rect 15436 21944 15442 21956
rect 15436 21916 15481 21944
rect 15436 21904 15442 21916
rect 15562 21904 15568 21956
rect 15620 21944 15626 21956
rect 17589 21947 17647 21953
rect 17589 21944 17601 21947
rect 15620 21916 17601 21944
rect 15620 21904 15626 21916
rect 17589 21913 17601 21916
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 17681 21947 17739 21953
rect 17681 21913 17693 21947
rect 17727 21913 17739 21947
rect 17681 21907 17739 21913
rect 16482 21876 16488 21888
rect 15120 21848 16488 21876
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 17696 21876 17724 21907
rect 17770 21904 17776 21956
rect 17828 21944 17834 21956
rect 20533 21947 20591 21953
rect 20533 21944 20545 21947
rect 17828 21916 20545 21944
rect 17828 21904 17834 21916
rect 20533 21913 20545 21916
rect 20579 21913 20591 21947
rect 20533 21907 20591 21913
rect 20625 21947 20683 21953
rect 20625 21913 20637 21947
rect 20671 21944 20683 21947
rect 20806 21944 20812 21956
rect 20671 21916 20812 21944
rect 20671 21913 20683 21916
rect 20625 21907 20683 21913
rect 20806 21904 20812 21916
rect 20864 21904 20870 21956
rect 21358 21904 21364 21956
rect 21416 21944 21422 21956
rect 21729 21947 21787 21953
rect 21729 21944 21741 21947
rect 21416 21916 21741 21944
rect 21416 21904 21422 21916
rect 21729 21913 21741 21916
rect 21775 21913 21787 21947
rect 21729 21907 21787 21913
rect 21821 21947 21879 21953
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 22370 21944 22376 21956
rect 21867 21916 22094 21944
rect 22331 21916 22376 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 16632 21848 17724 21876
rect 18785 21879 18843 21885
rect 16632 21836 16638 21848
rect 18785 21845 18797 21879
rect 18831 21876 18843 21879
rect 21082 21876 21088 21888
rect 18831 21848 21088 21876
rect 18831 21845 18843 21848
rect 18785 21839 18843 21845
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 22066 21876 22094 21916
rect 22370 21904 22376 21916
rect 22428 21904 22434 21956
rect 22480 21916 23336 21944
rect 22480 21876 22508 21916
rect 22066 21848 22508 21876
rect 23308 21876 23336 21916
rect 23382 21904 23388 21956
rect 23440 21944 23446 21956
rect 23584 21944 23612 21984
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 25240 22021 25268 22052
rect 27706 22040 27712 22092
rect 27764 22040 27770 22092
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24176 21984 24777 22012
rect 24176 21972 24182 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 22012 25283 22015
rect 25590 22012 25596 22024
rect 25271 21984 25596 22012
rect 25271 21981 25283 21984
rect 25225 21975 25283 21981
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 26234 22012 26240 22024
rect 26195 21984 26240 22012
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 27724 22012 27752 22040
rect 27646 21984 27752 22012
rect 24210 21944 24216 21956
rect 23440 21916 24216 21944
rect 23440 21904 23446 21916
rect 24210 21904 24216 21916
rect 24268 21904 24274 21956
rect 25314 21944 25320 21956
rect 25275 21916 25320 21944
rect 25314 21904 25320 21916
rect 25372 21904 25378 21956
rect 26510 21944 26516 21956
rect 26471 21916 26516 21944
rect 26510 21904 26516 21916
rect 26568 21904 26574 21956
rect 23569 21879 23627 21885
rect 23569 21876 23581 21879
rect 23308 21848 23581 21876
rect 23569 21845 23581 21848
rect 23615 21845 23627 21879
rect 24578 21876 24584 21888
rect 24539 21848 24584 21876
rect 23569 21839 23627 21845
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 25096 21848 27997 21876
rect 25096 21836 25102 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 27985 21839 28043 21845
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 7374 21672 7380 21684
rect 7335 21644 7380 21672
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 12710 21672 12716 21684
rect 11808 21644 12716 21672
rect 7282 21536 7288 21548
rect 7243 21508 7288 21536
rect 7282 21496 7288 21508
rect 7340 21496 7346 21548
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9950 21536 9956 21548
rect 9631 21508 9956 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21505 10563 21539
rect 10962 21536 10968 21548
rect 10923 21508 10968 21536
rect 10505 21499 10563 21505
rect 10520 21468 10548 21499
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11808 21545 11836 21644
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 20254 21672 20260 21684
rect 14424 21644 20260 21672
rect 14424 21632 14430 21644
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 20809 21675 20867 21681
rect 20809 21672 20821 21675
rect 20772 21644 20821 21672
rect 20772 21632 20778 21644
rect 20809 21641 20821 21644
rect 20855 21641 20867 21675
rect 24670 21672 24676 21684
rect 20809 21635 20867 21641
rect 22848 21644 24676 21672
rect 12618 21564 12624 21616
rect 12676 21604 12682 21616
rect 15746 21604 15752 21616
rect 12676 21576 15424 21604
rect 15659 21576 15752 21604
rect 12676 21564 12682 21576
rect 11793 21539 11851 21545
rect 11793 21505 11805 21539
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 13538 21536 13544 21548
rect 11931 21508 13544 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 13814 21536 13820 21548
rect 13727 21508 13820 21536
rect 13814 21496 13820 21508
rect 13872 21536 13878 21548
rect 14458 21536 14464 21548
rect 13872 21508 14464 21536
rect 13872 21496 13878 21508
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 14645 21539 14703 21545
rect 14645 21505 14657 21539
rect 14691 21536 14703 21539
rect 15010 21536 15016 21548
rect 14691 21508 15016 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 9416 21440 10548 21468
rect 9416 21409 9444 21440
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 12621 21471 12679 21477
rect 12492 21440 12537 21468
rect 12492 21428 12498 21440
rect 12621 21437 12633 21471
rect 12667 21437 12679 21471
rect 15102 21468 15108 21480
rect 15063 21440 15108 21468
rect 12621 21431 12679 21437
rect 9401 21403 9459 21409
rect 9401 21369 9413 21403
rect 9447 21369 9459 21403
rect 9401 21363 9459 21369
rect 11057 21403 11115 21409
rect 11057 21369 11069 21403
rect 11103 21400 11115 21403
rect 12636 21400 12664 21431
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 15212 21440 15301 21468
rect 11103 21372 12664 21400
rect 13909 21403 13967 21409
rect 11103 21369 11115 21372
rect 11057 21363 11115 21369
rect 13909 21369 13921 21403
rect 13955 21400 13967 21403
rect 15212 21400 15240 21440
rect 15289 21437 15301 21440
rect 15335 21437 15347 21471
rect 15396 21468 15424 21576
rect 15746 21564 15752 21576
rect 15804 21604 15810 21616
rect 17770 21604 17776 21616
rect 15804 21576 17776 21604
rect 15804 21564 15810 21576
rect 17770 21564 17776 21576
rect 17828 21564 17834 21616
rect 18506 21604 18512 21616
rect 17880 21576 18512 21604
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 17880 21536 17908 21576
rect 18506 21564 18512 21576
rect 18564 21564 18570 21616
rect 22186 21604 22192 21616
rect 19458 21576 22192 21604
rect 22186 21564 22192 21576
rect 22244 21564 22250 21616
rect 22848 21604 22876 21644
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 24854 21632 24860 21684
rect 24912 21672 24918 21684
rect 26513 21675 26571 21681
rect 26513 21672 26525 21675
rect 24912 21644 26525 21672
rect 24912 21632 24918 21644
rect 26513 21641 26525 21644
rect 26559 21641 26571 21675
rect 26513 21635 26571 21641
rect 23014 21604 23020 21616
rect 22756 21576 22876 21604
rect 22975 21576 23020 21604
rect 16899 21508 17908 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 17788 21480 17816 21508
rect 20070 21496 20076 21548
rect 20128 21536 20134 21548
rect 20165 21539 20223 21545
rect 20165 21536 20177 21539
rect 20128 21508 20177 21536
rect 20128 21496 20134 21508
rect 20165 21505 20177 21508
rect 20211 21505 20223 21539
rect 20165 21499 20223 21505
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 22554 21536 22560 21548
rect 22051 21508 22560 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 22756 21545 22784 21576
rect 23014 21564 23020 21576
rect 23072 21564 23078 21616
rect 23474 21564 23480 21616
rect 23532 21564 23538 21616
rect 24486 21564 24492 21616
rect 24544 21564 24550 21616
rect 24578 21564 24584 21616
rect 24636 21604 24642 21616
rect 24636 21576 28120 21604
rect 24636 21564 24642 21576
rect 22741 21539 22799 21545
rect 22741 21505 22753 21539
rect 22787 21505 22799 21539
rect 24504 21536 24532 21564
rect 24504 21508 24624 21536
rect 22741 21499 22799 21505
rect 17678 21468 17684 21480
rect 15396 21440 17684 21468
rect 15289 21431 15347 21437
rect 17678 21428 17684 21440
rect 17736 21428 17742 21480
rect 17770 21428 17776 21480
rect 17828 21428 17834 21480
rect 17954 21468 17960 21480
rect 17915 21440 17960 21468
rect 17954 21428 17960 21440
rect 18012 21428 18018 21480
rect 18230 21468 18236 21480
rect 18191 21440 18236 21468
rect 18230 21428 18236 21440
rect 18288 21468 18294 21480
rect 18966 21468 18972 21480
rect 18288 21440 18972 21468
rect 18288 21428 18294 21440
rect 18966 21428 18972 21440
rect 19024 21428 19030 21480
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 23382 21468 23388 21480
rect 19300 21440 23388 21468
rect 19300 21428 19306 21440
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 23566 21428 23572 21480
rect 23624 21468 23630 21480
rect 24486 21468 24492 21480
rect 23624 21440 24492 21468
rect 23624 21428 23630 21440
rect 24486 21428 24492 21440
rect 24544 21428 24550 21480
rect 24596 21468 24624 21508
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 26234 21536 26240 21548
rect 24728 21508 26240 21536
rect 24728 21496 24734 21508
rect 26234 21496 26240 21508
rect 26292 21496 26298 21548
rect 26421 21539 26479 21545
rect 26421 21505 26433 21539
rect 26467 21505 26479 21539
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 26421 21499 26479 21505
rect 24762 21468 24768 21480
rect 24596 21440 24768 21468
rect 24762 21428 24768 21440
rect 24820 21428 24826 21480
rect 26436 21468 26464 21499
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 28092 21545 28120 21576
rect 28077 21539 28135 21545
rect 28077 21505 28089 21539
rect 28123 21505 28135 21539
rect 28077 21499 28135 21505
rect 28166 21468 28172 21480
rect 26436 21440 28172 21468
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 13955 21372 15240 21400
rect 13955 21369 13967 21372
rect 13909 21363 13967 21369
rect 19610 21360 19616 21412
rect 19668 21400 19674 21412
rect 19668 21372 22876 21400
rect 19668 21360 19674 21372
rect 10318 21332 10324 21344
rect 10279 21304 10324 21332
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 11882 21292 11888 21344
rect 11940 21332 11946 21344
rect 12250 21332 12256 21344
rect 11940 21304 12256 21332
rect 11940 21292 11946 21304
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12805 21335 12863 21341
rect 12805 21332 12817 21335
rect 12492 21304 12817 21332
rect 12492 21292 12498 21304
rect 12805 21301 12817 21304
rect 12851 21301 12863 21335
rect 12805 21295 12863 21301
rect 14461 21335 14519 21341
rect 14461 21301 14473 21335
rect 14507 21332 14519 21335
rect 15654 21332 15660 21344
rect 14507 21304 15660 21332
rect 14507 21301 14519 21304
rect 14461 21295 14519 21301
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17862 21332 17868 21344
rect 16991 21304 17868 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 19702 21332 19708 21344
rect 19663 21304 19708 21332
rect 19702 21292 19708 21304
rect 19760 21292 19766 21344
rect 20254 21332 20260 21344
rect 20215 21304 20260 21332
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21332 22155 21335
rect 22278 21332 22284 21344
rect 22143 21304 22284 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 22848 21332 22876 21372
rect 24210 21360 24216 21412
rect 24268 21400 24274 21412
rect 25774 21400 25780 21412
rect 24268 21372 25780 21400
rect 24268 21360 24274 21372
rect 25774 21360 25780 21372
rect 25832 21360 25838 21412
rect 24026 21332 24032 21344
rect 22848 21304 24032 21332
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 27249 21335 27307 21341
rect 27249 21301 27261 21335
rect 27295 21332 27307 21335
rect 28074 21332 28080 21344
rect 27295 21304 28080 21332
rect 27295 21301 27307 21304
rect 27249 21295 27307 21301
rect 28074 21292 28080 21304
rect 28132 21292 28138 21344
rect 28258 21332 28264 21344
rect 28219 21304 28264 21332
rect 28258 21292 28264 21304
rect 28316 21292 28322 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 11149 21131 11207 21137
rect 11149 21097 11161 21131
rect 11195 21128 11207 21131
rect 12158 21128 12164 21140
rect 11195 21100 12164 21128
rect 11195 21097 11207 21100
rect 11149 21091 11207 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 15105 21131 15163 21137
rect 15105 21097 15117 21131
rect 15151 21128 15163 21131
rect 15746 21128 15752 21140
rect 15151 21100 15752 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 15933 21131 15991 21137
rect 15933 21097 15945 21131
rect 15979 21128 15991 21131
rect 16574 21128 16580 21140
rect 15979 21100 16580 21128
rect 15979 21097 15991 21100
rect 15933 21091 15991 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17034 21088 17040 21140
rect 17092 21128 17098 21140
rect 17773 21131 17831 21137
rect 17773 21128 17785 21131
rect 17092 21100 17785 21128
rect 17092 21088 17098 21100
rect 17773 21097 17785 21100
rect 17819 21097 17831 21131
rect 19610 21128 19616 21140
rect 17773 21091 17831 21097
rect 17880 21100 19616 21128
rect 13354 21020 13360 21072
rect 13412 21060 13418 21072
rect 13449 21063 13507 21069
rect 13449 21060 13461 21063
rect 13412 21032 13461 21060
rect 13412 21020 13418 21032
rect 13449 21029 13461 21032
rect 13495 21029 13507 21063
rect 15194 21060 15200 21072
rect 13449 21023 13507 21029
rect 14568 21032 15200 21060
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 14568 21001 14596 21032
rect 15194 21020 15200 21032
rect 15252 21020 15258 21072
rect 17221 21063 17279 21069
rect 17221 21029 17233 21063
rect 17267 21060 17279 21063
rect 17880 21060 17908 21100
rect 19610 21088 19616 21100
rect 19668 21088 19674 21140
rect 20162 21088 20168 21140
rect 20220 21128 20226 21140
rect 20514 21131 20572 21137
rect 20514 21128 20526 21131
rect 20220 21100 20526 21128
rect 20220 21088 20226 21100
rect 20514 21097 20526 21100
rect 20560 21097 20572 21131
rect 20514 21091 20572 21097
rect 20622 21088 20628 21140
rect 20680 21128 20686 21140
rect 23106 21128 23112 21140
rect 20680 21100 21588 21128
rect 23067 21100 23112 21128
rect 20680 21088 20686 21100
rect 21560 21060 21588 21100
rect 23106 21088 23112 21100
rect 23164 21088 23170 21140
rect 24118 21128 24124 21140
rect 23768 21100 24124 21128
rect 22005 21063 22063 21069
rect 22005 21060 22017 21063
rect 17267 21032 17908 21060
rect 17972 21032 20392 21060
rect 21560 21032 22017 21060
rect 17267 21029 17279 21032
rect 17221 21023 17279 21029
rect 13265 20995 13323 21001
rect 13265 20992 13277 20995
rect 10376 20964 13277 20992
rect 10376 20952 10382 20964
rect 13265 20961 13277 20964
rect 13311 20961 13323 20995
rect 13265 20955 13323 20961
rect 14553 20995 14611 21001
rect 14553 20961 14565 20995
rect 14599 20961 14611 20995
rect 14734 20992 14740 21004
rect 14695 20964 14740 20992
rect 14553 20955 14611 20961
rect 14734 20952 14740 20964
rect 14792 20952 14798 21004
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 6086 20924 6092 20936
rect 6047 20896 6092 20924
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 10226 20924 10232 20936
rect 10187 20896 10232 20924
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 11057 20927 11115 20933
rect 11057 20893 11069 20927
rect 11103 20924 11115 20927
rect 11146 20924 11152 20936
rect 11103 20896 11152 20924
rect 11103 20893 11115 20896
rect 11057 20887 11115 20893
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11940 20896 11989 20924
rect 11940 20884 11946 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 12158 20924 12164 20936
rect 12119 20896 12164 20924
rect 11977 20887 12035 20893
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 12526 20884 12532 20936
rect 12584 20924 12590 20936
rect 13081 20927 13139 20933
rect 13081 20924 13093 20927
rect 12584 20896 13093 20924
rect 12584 20884 12590 20896
rect 13081 20893 13093 20896
rect 13127 20893 13139 20927
rect 13081 20887 13139 20893
rect 14642 20884 14648 20936
rect 14700 20924 14706 20936
rect 17972 20933 18000 21032
rect 19242 20952 19248 21004
rect 19300 20992 19306 21004
rect 20257 20995 20315 21001
rect 20257 20992 20269 20995
rect 19300 20964 20269 20992
rect 19300 20952 19306 20964
rect 20257 20961 20269 20964
rect 20303 20961 20315 20995
rect 20364 20992 20392 21032
rect 22005 21029 22017 21032
rect 22051 21029 22063 21063
rect 22005 21023 22063 21029
rect 23661 21063 23719 21069
rect 23661 21029 23673 21063
rect 23707 21060 23719 21063
rect 23768 21060 23796 21100
rect 24118 21088 24124 21100
rect 24176 21088 24182 21140
rect 23707 21032 23796 21060
rect 23707 21029 23719 21032
rect 23661 21023 23719 21029
rect 20364 20964 21772 20992
rect 20257 20955 20315 20961
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 14700 20896 16129 20924
rect 14700 20884 14706 20896
rect 16117 20893 16129 20896
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 17957 20927 18015 20933
rect 17957 20893 17969 20927
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20924 18475 20927
rect 18690 20924 18696 20936
rect 18463 20896 18696 20924
rect 18463 20893 18475 20896
rect 18417 20887 18475 20893
rect 18690 20884 18696 20896
rect 18748 20924 18754 20936
rect 19334 20924 19340 20936
rect 18748 20896 19340 20924
rect 18748 20884 18754 20896
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20926 19487 20927
rect 19518 20926 19524 20936
rect 19475 20898 19524 20926
rect 19475 20893 19487 20898
rect 19429 20887 19487 20893
rect 19518 20884 19524 20898
rect 19576 20884 19582 20936
rect 21744 20924 21772 20964
rect 21818 20952 21824 21004
rect 21876 20992 21882 21004
rect 22465 20995 22523 21001
rect 22465 20992 22477 20995
rect 21876 20964 22477 20992
rect 21876 20952 21882 20964
rect 22465 20961 22477 20964
rect 22511 20961 22523 20995
rect 22465 20955 22523 20961
rect 22649 20995 22707 21001
rect 22649 20961 22661 20995
rect 22695 20992 22707 20995
rect 22830 20992 22836 21004
rect 22695 20964 22836 20992
rect 22695 20961 22707 20964
rect 22649 20955 22707 20961
rect 22830 20952 22836 20964
rect 22888 20952 22894 21004
rect 24762 20992 24768 21004
rect 22940 20964 24768 20992
rect 22940 20924 22968 20964
rect 24762 20952 24768 20964
rect 24820 20952 24826 21004
rect 26234 20952 26240 21004
rect 26292 20992 26298 21004
rect 26329 20995 26387 21001
rect 26329 20992 26341 20995
rect 26292 20964 26341 20992
rect 26292 20952 26298 20964
rect 26329 20961 26341 20964
rect 26375 20961 26387 20995
rect 26329 20955 26387 20961
rect 21744 20896 22968 20924
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 24026 20924 24032 20936
rect 23615 20896 24032 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 24026 20884 24032 20896
rect 24084 20884 24090 20936
rect 15562 20856 15568 20868
rect 12406 20828 15568 20856
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 3970 20788 3976 20800
rect 1627 20760 3976 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 3970 20748 3976 20760
rect 4028 20748 4034 20800
rect 6178 20788 6184 20800
rect 6139 20760 6184 20788
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20788 9643 20791
rect 9858 20788 9864 20800
rect 9631 20760 9864 20788
rect 9631 20757 9643 20760
rect 9585 20751 9643 20757
rect 9858 20748 9864 20760
rect 9916 20748 9922 20800
rect 10318 20788 10324 20800
rect 10279 20760 10324 20788
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 10502 20748 10508 20800
rect 10560 20788 10566 20800
rect 12406 20788 12434 20828
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 16666 20856 16672 20868
rect 16627 20828 16672 20856
rect 16666 20816 16672 20828
rect 16724 20816 16730 20868
rect 16758 20816 16764 20868
rect 16816 20856 16822 20868
rect 16816 20828 16861 20856
rect 16960 20828 19288 20856
rect 16816 20816 16822 20828
rect 10560 20760 12434 20788
rect 12621 20791 12679 20797
rect 10560 20748 10566 20760
rect 12621 20757 12633 20791
rect 12667 20788 12679 20791
rect 12802 20788 12808 20800
rect 12667 20760 12808 20788
rect 12667 20757 12679 20760
rect 12621 20751 12679 20757
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15378 20788 15384 20800
rect 15252 20760 15384 20788
rect 15252 20748 15258 20760
rect 15378 20748 15384 20760
rect 15436 20788 15442 20800
rect 16960 20788 16988 20828
rect 15436 20760 16988 20788
rect 18509 20791 18567 20797
rect 15436 20748 15442 20760
rect 18509 20757 18521 20791
rect 18555 20788 18567 20791
rect 19150 20788 19156 20800
rect 18555 20760 19156 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 19150 20748 19156 20760
rect 19208 20748 19214 20800
rect 19260 20788 19288 20828
rect 21082 20816 21088 20868
rect 21140 20816 21146 20868
rect 26605 20859 26663 20865
rect 26605 20856 26617 20859
rect 23216 20828 26617 20856
rect 19521 20791 19579 20797
rect 19521 20788 19533 20791
rect 19260 20760 19533 20788
rect 19521 20757 19533 20760
rect 19567 20757 19579 20791
rect 19521 20751 19579 20757
rect 22830 20748 22836 20800
rect 22888 20788 22894 20800
rect 23216 20788 23244 20828
rect 26605 20825 26617 20828
rect 26651 20825 26663 20859
rect 26605 20819 26663 20825
rect 27614 20816 27620 20868
rect 27672 20816 27678 20868
rect 28258 20816 28264 20868
rect 28316 20856 28322 20868
rect 28353 20859 28411 20865
rect 28353 20856 28365 20859
rect 28316 20828 28365 20856
rect 28316 20816 28322 20828
rect 28353 20825 28365 20828
rect 28399 20825 28411 20859
rect 28353 20819 28411 20825
rect 22888 20760 23244 20788
rect 22888 20748 22894 20760
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 10502 20584 10508 20596
rect 10463 20556 10508 20584
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 10962 20544 10968 20596
rect 11020 20584 11026 20596
rect 11020 20556 12434 20584
rect 11020 20544 11026 20556
rect 12406 20516 12434 20556
rect 12986 20544 12992 20596
rect 13044 20584 13050 20596
rect 18138 20584 18144 20596
rect 13044 20556 18144 20584
rect 13044 20544 13050 20556
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 21358 20584 21364 20596
rect 18288 20556 21364 20584
rect 18288 20544 18294 20556
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 21692 20556 22017 20584
rect 21692 20544 21698 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 22462 20544 22468 20596
rect 22520 20584 22526 20596
rect 26418 20584 26424 20596
rect 22520 20556 26424 20584
rect 22520 20544 22526 20556
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 27890 20584 27896 20596
rect 27851 20556 27896 20584
rect 27890 20544 27896 20556
rect 27948 20544 27954 20596
rect 18325 20519 18383 20525
rect 18325 20516 18337 20519
rect 12406 20488 18337 20516
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 9858 20448 9864 20460
rect 9819 20420 9864 20448
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 10042 20448 10048 20460
rect 10003 20420 10048 20448
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 11020 20420 11161 20448
rect 11020 20408 11026 20420
rect 11149 20417 11161 20420
rect 11195 20417 11207 20451
rect 11698 20448 11704 20460
rect 11659 20420 11704 20448
rect 11149 20411 11207 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20448 12863 20451
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 12851 20420 14565 20448
rect 12851 20417 12863 20420
rect 12805 20411 12863 20417
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15712 20420 16037 20448
rect 15712 20408 15718 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20448 16911 20451
rect 17126 20448 17132 20460
rect 16899 20420 17132 20448
rect 16899 20417 16911 20420
rect 16853 20411 16911 20417
rect 17126 20408 17132 20420
rect 17184 20448 17190 20460
rect 17494 20448 17500 20460
rect 17184 20420 17500 20448
rect 17184 20408 17190 20420
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 4617 20383 4675 20389
rect 4617 20349 4629 20383
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 4801 20383 4859 20389
rect 4801 20349 4813 20383
rect 4847 20380 4859 20383
rect 6086 20380 6092 20392
rect 4847 20352 6092 20380
rect 4847 20349 4859 20352
rect 4801 20343 4859 20349
rect 4632 20312 4660 20343
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 11885 20383 11943 20389
rect 11885 20380 11897 20383
rect 11112 20352 11897 20380
rect 11112 20340 11118 20352
rect 11885 20349 11897 20352
rect 11931 20349 11943 20383
rect 13446 20380 13452 20392
rect 13407 20352 13452 20380
rect 11885 20343 11943 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13538 20340 13544 20392
rect 13596 20380 13602 20392
rect 13633 20383 13691 20389
rect 13633 20380 13645 20383
rect 13596 20352 13645 20380
rect 13596 20340 13602 20352
rect 13633 20349 13645 20352
rect 13679 20349 13691 20383
rect 14734 20380 14740 20392
rect 14695 20352 14740 20380
rect 13633 20343 13691 20349
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 17880 20380 17908 20488
rect 18325 20485 18337 20488
rect 18371 20485 18383 20519
rect 18325 20479 18383 20485
rect 19702 20476 19708 20528
rect 19760 20516 19766 20528
rect 19760 20488 21036 20516
rect 19760 20476 19766 20488
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 18012 20420 18061 20448
rect 18012 20408 18018 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 19426 20408 19432 20460
rect 19484 20408 19490 20460
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 20901 20451 20959 20457
rect 20901 20448 20913 20451
rect 19668 20420 20913 20448
rect 19668 20408 19674 20420
rect 20901 20417 20913 20420
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 20257 20383 20315 20389
rect 17880 20352 20208 20380
rect 5074 20312 5080 20324
rect 4632 20284 5080 20312
rect 5074 20272 5080 20284
rect 5132 20272 5138 20324
rect 14093 20315 14151 20321
rect 14093 20281 14105 20315
rect 14139 20312 14151 20315
rect 15194 20312 15200 20324
rect 14139 20284 15200 20312
rect 14139 20281 14151 20284
rect 14093 20275 14151 20281
rect 15194 20272 15200 20284
rect 15252 20272 15258 20324
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 20070 20312 20076 20324
rect 19484 20284 20076 20312
rect 19484 20272 19490 20284
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 5718 20244 5724 20256
rect 5307 20216 5724 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 7800 20216 8861 20244
rect 7800 20204 7806 20216
rect 8849 20213 8861 20216
rect 8895 20213 8907 20247
rect 8849 20207 8907 20213
rect 10965 20247 11023 20253
rect 10965 20213 10977 20247
rect 11011 20244 11023 20247
rect 11698 20244 11704 20256
rect 11011 20216 11704 20244
rect 11011 20213 11023 20216
rect 10965 20207 11023 20213
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 12345 20247 12403 20253
rect 12345 20213 12357 20247
rect 12391 20244 12403 20247
rect 12434 20244 12440 20256
rect 12391 20216 12440 20244
rect 12391 20213 12403 20216
rect 12345 20207 12403 20213
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 14366 20204 14372 20256
rect 14424 20244 14430 20256
rect 14921 20247 14979 20253
rect 14921 20244 14933 20247
rect 14424 20216 14933 20244
rect 14424 20204 14430 20216
rect 14921 20213 14933 20216
rect 14967 20213 14979 20247
rect 14921 20207 14979 20213
rect 15841 20247 15899 20253
rect 15841 20213 15853 20247
rect 15887 20244 15899 20247
rect 16758 20244 16764 20256
rect 15887 20216 16764 20244
rect 15887 20213 15899 20216
rect 15841 20207 15899 20213
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 16945 20247 17003 20253
rect 16945 20213 16957 20247
rect 16991 20244 17003 20247
rect 19058 20244 19064 20256
rect 16991 20216 19064 20244
rect 16991 20213 17003 20216
rect 16945 20207 17003 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19797 20247 19855 20253
rect 19797 20244 19809 20247
rect 19392 20216 19809 20244
rect 19392 20204 19398 20216
rect 19797 20213 19809 20216
rect 19843 20213 19855 20247
rect 20180 20244 20208 20352
rect 20257 20349 20269 20383
rect 20303 20349 20315 20383
rect 20438 20380 20444 20392
rect 20399 20352 20444 20380
rect 20257 20343 20315 20349
rect 20272 20312 20300 20343
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 21008 20380 21036 20488
rect 23474 20476 23480 20528
rect 23532 20516 23538 20528
rect 23532 20488 23966 20516
rect 23532 20476 23538 20488
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 28074 20448 28080 20460
rect 21692 20446 21864 20448
rect 21928 20446 23244 20448
rect 21692 20420 23244 20446
rect 28035 20420 28080 20448
rect 21692 20408 21698 20420
rect 21836 20418 21956 20420
rect 22002 20380 22008 20392
rect 21008 20352 22008 20380
rect 22002 20340 22008 20352
rect 22060 20340 22066 20392
rect 23216 20389 23244 20420
rect 28074 20408 28080 20420
rect 28132 20408 28138 20460
rect 23201 20383 23259 20389
rect 23201 20349 23213 20383
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 23477 20383 23535 20389
rect 23477 20349 23489 20383
rect 23523 20380 23535 20383
rect 23566 20380 23572 20392
rect 23523 20352 23572 20380
rect 23523 20349 23535 20352
rect 23477 20343 23535 20349
rect 23106 20312 23112 20324
rect 20272 20284 23112 20312
rect 23106 20272 23112 20284
rect 23164 20272 23170 20324
rect 20714 20244 20720 20256
rect 20180 20216 20720 20244
rect 19797 20207 19855 20213
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21358 20204 21364 20256
rect 21416 20244 21422 20256
rect 23014 20244 23020 20256
rect 21416 20216 23020 20244
rect 21416 20204 21422 20216
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 23216 20244 23244 20343
rect 23566 20340 23572 20352
rect 23624 20340 23630 20392
rect 25038 20340 25044 20392
rect 25096 20380 25102 20392
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 25096 20352 25237 20380
rect 25096 20340 25102 20352
rect 25225 20349 25237 20352
rect 25271 20349 25283 20383
rect 25225 20343 25283 20349
rect 24670 20244 24676 20256
rect 23216 20216 24676 20244
rect 24670 20204 24676 20216
rect 24728 20204 24734 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 5074 20040 5080 20052
rect 5035 20012 5080 20040
rect 5074 20000 5080 20012
rect 5132 20000 5138 20052
rect 6086 20000 6092 20052
rect 6144 20040 6150 20052
rect 6181 20043 6239 20049
rect 6181 20040 6193 20043
rect 6144 20012 6193 20040
rect 6144 20000 6150 20012
rect 6181 20009 6193 20012
rect 6227 20009 6239 20043
rect 6181 20003 6239 20009
rect 11057 20043 11115 20049
rect 11057 20009 11069 20043
rect 11103 20040 11115 20043
rect 12158 20040 12164 20052
rect 11103 20012 12164 20040
rect 11103 20009 11115 20012
rect 11057 20003 11115 20009
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 12897 20043 12955 20049
rect 12897 20009 12909 20043
rect 12943 20040 12955 20043
rect 14734 20040 14740 20052
rect 12943 20012 14740 20040
rect 12943 20009 12955 20012
rect 12897 20003 12955 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 17770 20040 17776 20052
rect 16172 20012 17776 20040
rect 16172 20000 16178 20012
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18414 20040 18420 20052
rect 18012 20012 18420 20040
rect 18012 20000 18018 20012
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 22186 20040 22192 20052
rect 19306 20012 22192 20040
rect 18230 19972 18236 19984
rect 15212 19944 18236 19972
rect 1762 19836 1768 19848
rect 1723 19808 1768 19836
rect 1762 19796 1768 19808
rect 1820 19796 1826 19848
rect 4062 19796 4068 19848
rect 4120 19836 4126 19848
rect 5077 19839 5135 19845
rect 5077 19836 5089 19839
rect 4120 19808 5089 19836
rect 4120 19796 4126 19808
rect 5077 19805 5089 19808
rect 5123 19805 5135 19839
rect 5077 19799 5135 19805
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19836 6147 19839
rect 6730 19836 6736 19848
rect 6135 19808 6736 19836
rect 6135 19805 6147 19808
rect 6089 19799 6147 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 9122 19836 9128 19848
rect 9083 19808 9128 19836
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19836 10563 19839
rect 10778 19836 10784 19848
rect 10551 19808 10784 19836
rect 10551 19805 10563 19808
rect 10505 19799 10563 19805
rect 10778 19796 10784 19808
rect 10836 19836 10842 19848
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 10836 19808 10977 19836
rect 10836 19796 10842 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11609 19839 11667 19845
rect 11609 19805 11621 19839
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 11624 19768 11652 19799
rect 11974 19796 11980 19848
rect 12032 19836 12038 19848
rect 13081 19839 13139 19845
rect 13081 19836 13093 19839
rect 12032 19808 13093 19836
rect 12032 19796 12038 19808
rect 13081 19805 13093 19808
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 14090 19836 14096 19848
rect 13771 19808 14096 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 15212 19836 15240 19944
rect 18230 19932 18236 19944
rect 18288 19932 18294 19984
rect 19306 19972 19334 20012
rect 22186 20000 22192 20012
rect 22244 20040 22250 20052
rect 22244 20012 23060 20040
rect 22244 20000 22250 20012
rect 18340 19944 19334 19972
rect 21269 19975 21327 19981
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 16850 19904 16856 19916
rect 15335 19876 16856 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 18340 19904 18368 19944
rect 21269 19941 21281 19975
rect 21315 19972 21327 19975
rect 21542 19972 21548 19984
rect 21315 19944 21548 19972
rect 21315 19941 21327 19944
rect 21269 19935 21327 19941
rect 21542 19932 21548 19944
rect 21600 19932 21606 19984
rect 23032 19972 23060 20012
rect 23106 20000 23112 20052
rect 23164 20040 23170 20052
rect 25958 20040 25964 20052
rect 23164 20012 25964 20040
rect 23164 20000 23170 20012
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 28166 20040 28172 20052
rect 28127 20012 28172 20040
rect 28166 20000 28172 20012
rect 28224 20000 28230 20052
rect 23032 19944 24808 19972
rect 18248 19876 18368 19904
rect 14875 19808 15240 19836
rect 15473 19839 15531 19845
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15473 19805 15485 19839
rect 15519 19836 15531 19839
rect 16022 19836 16028 19848
rect 15519 19808 16028 19836
rect 15519 19805 15531 19808
rect 15473 19799 15531 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 17770 19836 17776 19848
rect 17731 19808 17776 19836
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19836 17923 19839
rect 18138 19836 18144 19848
rect 17911 19808 18144 19836
rect 17911 19805 17923 19808
rect 17865 19799 17923 19805
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18248 19836 18276 19876
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 19242 19904 19248 19916
rect 18656 19876 19248 19904
rect 18656 19864 18662 19876
rect 19242 19864 19248 19876
rect 19300 19904 19306 19916
rect 19521 19907 19579 19913
rect 19521 19904 19533 19907
rect 19300 19876 19533 19904
rect 19300 19864 19306 19876
rect 19521 19873 19533 19876
rect 19567 19904 19579 19907
rect 21634 19904 21640 19916
rect 19567 19876 21640 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 21634 19864 21640 19876
rect 21692 19904 21698 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 21692 19876 21741 19904
rect 21692 19864 21698 19876
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 22002 19904 22008 19916
rect 21963 19876 22008 19904
rect 21729 19867 21787 19873
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 24670 19904 24676 19916
rect 24631 19876 24676 19904
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 24780 19904 24808 19944
rect 26050 19932 26056 19984
rect 26108 19932 26114 19984
rect 26068 19904 26096 19932
rect 24780 19876 26096 19904
rect 18409 19849 18467 19855
rect 18409 19846 18421 19849
rect 18340 19836 18421 19846
rect 18248 19818 18421 19836
rect 18248 19808 18368 19818
rect 18409 19815 18421 19818
rect 18455 19815 18467 19849
rect 18409 19809 18467 19815
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19426 19836 19432 19848
rect 18748 19808 19432 19836
rect 18748 19796 18754 19808
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 21266 19836 21272 19848
rect 20930 19808 21272 19836
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 28350 19836 28356 19848
rect 28311 19808 28356 19836
rect 28350 19796 28356 19808
rect 28408 19796 28414 19848
rect 13262 19768 13268 19780
rect 11624 19740 13268 19768
rect 13262 19728 13268 19740
rect 13320 19768 13326 19780
rect 15933 19771 15991 19777
rect 15933 19768 15945 19771
rect 13320 19740 15945 19768
rect 13320 19728 13326 19740
rect 15933 19737 15945 19740
rect 15979 19737 15991 19771
rect 15933 19731 15991 19737
rect 16669 19771 16727 19777
rect 16669 19737 16681 19771
rect 16715 19737 16727 19771
rect 16669 19731 16727 19737
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 3694 19700 3700 19712
rect 1627 19672 3700 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 3694 19660 3700 19672
rect 3752 19660 3758 19712
rect 9214 19700 9220 19712
rect 9175 19672 9220 19700
rect 9214 19660 9220 19672
rect 9272 19660 9278 19712
rect 10321 19703 10379 19709
rect 10321 19669 10333 19703
rect 10367 19700 10379 19703
rect 10502 19700 10508 19712
rect 10367 19672 10508 19700
rect 10367 19669 10379 19672
rect 10321 19663 10379 19669
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 11146 19660 11152 19712
rect 11204 19700 11210 19712
rect 11701 19703 11759 19709
rect 11701 19700 11713 19703
rect 11204 19672 11713 19700
rect 11204 19660 11210 19672
rect 11701 19669 11713 19672
rect 11747 19669 11759 19703
rect 11701 19663 11759 19669
rect 12253 19703 12311 19709
rect 12253 19669 12265 19703
rect 12299 19700 12311 19703
rect 12618 19700 12624 19712
rect 12299 19672 12624 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13538 19700 13544 19712
rect 13499 19672 13544 19700
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 14645 19703 14703 19709
rect 14645 19669 14657 19703
rect 14691 19700 14703 19703
rect 15654 19700 15660 19712
rect 14691 19672 15660 19700
rect 14691 19669 14703 19672
rect 14645 19663 14703 19669
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 16684 19700 16712 19731
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17313 19771 17371 19777
rect 16816 19740 16861 19768
rect 16816 19728 16822 19740
rect 17313 19737 17325 19771
rect 17359 19768 17371 19771
rect 19797 19771 19855 19777
rect 17359 19740 19748 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 17494 19700 17500 19712
rect 16684 19672 17500 19700
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18104 19672 18521 19700
rect 18104 19660 18110 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 18690 19660 18696 19712
rect 18748 19700 18754 19712
rect 19610 19700 19616 19712
rect 18748 19672 19616 19700
rect 18748 19660 18754 19672
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 19720 19700 19748 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 19886 19768 19892 19780
rect 19843 19740 19892 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 21910 19768 21916 19780
rect 21192 19740 21916 19768
rect 21192 19700 21220 19740
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22462 19728 22468 19780
rect 22520 19728 22526 19780
rect 23290 19728 23296 19780
rect 23348 19768 23354 19780
rect 23348 19740 23612 19768
rect 23348 19728 23354 19740
rect 19720 19672 21220 19700
rect 21358 19660 21364 19712
rect 21416 19700 21422 19712
rect 23477 19703 23535 19709
rect 23477 19700 23489 19703
rect 21416 19672 23489 19700
rect 21416 19660 21422 19672
rect 23477 19669 23489 19672
rect 23523 19669 23535 19703
rect 23584 19700 23612 19740
rect 24486 19728 24492 19780
rect 24544 19768 24550 19780
rect 24949 19771 25007 19777
rect 24949 19768 24961 19771
rect 24544 19740 24961 19768
rect 24544 19728 24550 19740
rect 24949 19737 24961 19740
rect 24995 19737 25007 19771
rect 26694 19768 26700 19780
rect 24949 19731 25007 19737
rect 25056 19740 25438 19768
rect 26655 19740 26700 19768
rect 25056 19700 25084 19740
rect 26694 19728 26700 19740
rect 26752 19728 26758 19780
rect 23584 19672 25084 19700
rect 23477 19663 23535 19669
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 6549 19499 6607 19505
rect 6549 19465 6561 19499
rect 6595 19465 6607 19499
rect 6549 19459 6607 19465
rect 10321 19499 10379 19505
rect 10321 19465 10333 19499
rect 10367 19465 10379 19499
rect 10962 19496 10968 19508
rect 10923 19468 10968 19496
rect 10321 19459 10379 19465
rect 6564 19428 6592 19459
rect 10336 19428 10364 19459
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11974 19496 11980 19508
rect 11935 19468 11980 19496
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 13262 19496 13268 19508
rect 13223 19468 13268 19496
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 14366 19496 14372 19508
rect 14327 19468 14372 19496
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 14829 19499 14887 19505
rect 14829 19496 14841 19499
rect 14608 19468 14841 19496
rect 14608 19456 14614 19468
rect 14829 19465 14841 19468
rect 14875 19465 14887 19499
rect 16022 19496 16028 19508
rect 15983 19468 16028 19496
rect 14829 19459 14887 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 17589 19499 17647 19505
rect 17589 19465 17601 19499
rect 17635 19496 17647 19499
rect 22462 19496 22468 19508
rect 17635 19468 22468 19496
rect 17635 19465 17647 19468
rect 17589 19459 17647 19465
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 23014 19456 23020 19508
rect 23072 19496 23078 19508
rect 24121 19499 24179 19505
rect 24121 19496 24133 19499
rect 23072 19468 24133 19496
rect 23072 19456 23078 19468
rect 24121 19465 24133 19468
rect 24167 19465 24179 19499
rect 24121 19459 24179 19465
rect 26418 19456 26424 19508
rect 26476 19496 26482 19508
rect 26513 19499 26571 19505
rect 26513 19496 26525 19499
rect 26476 19468 26525 19496
rect 26476 19456 26482 19468
rect 26513 19465 26525 19468
rect 26559 19465 26571 19499
rect 26513 19459 26571 19465
rect 11054 19428 11060 19440
rect 6564 19400 7604 19428
rect 10336 19400 11060 19428
rect 6730 19360 6736 19372
rect 6691 19332 6736 19360
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 7576 19369 7604 19400
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 11164 19400 13308 19428
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 9950 19360 9956 19372
rect 9907 19332 9956 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 10502 19360 10508 19372
rect 10463 19332 10508 19360
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 11164 19369 11192 19400
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 12161 19363 12219 19369
rect 12161 19334 12173 19363
rect 11149 19323 11207 19329
rect 12084 19329 12173 19334
rect 12207 19329 12219 19363
rect 12618 19360 12624 19372
rect 12579 19332 12624 19360
rect 12084 19323 12219 19329
rect 12084 19306 12204 19323
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 13280 19360 13308 19400
rect 13354 19388 13360 19440
rect 13412 19428 13418 19440
rect 18690 19428 18696 19440
rect 13412 19400 18696 19428
rect 13412 19388 13418 19400
rect 18690 19388 18696 19400
rect 18748 19388 18754 19440
rect 20990 19428 20996 19440
rect 19642 19400 20996 19428
rect 20990 19388 20996 19400
rect 21048 19388 21054 19440
rect 21542 19388 21548 19440
rect 21600 19428 21606 19440
rect 22649 19431 22707 19437
rect 22649 19428 22661 19431
rect 21600 19400 22661 19428
rect 21600 19388 21606 19400
rect 22649 19397 22661 19400
rect 22695 19397 22707 19431
rect 22649 19391 22707 19397
rect 25130 19388 25136 19440
rect 25188 19428 25194 19440
rect 25188 19400 25530 19428
rect 25188 19388 25194 19400
rect 13280 19332 13492 19360
rect 12084 19224 12112 19306
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12268 19264 12817 19292
rect 12158 19224 12164 19236
rect 12084 19196 12164 19224
rect 12158 19184 12164 19196
rect 12216 19184 12222 19236
rect 7374 19156 7380 19168
rect 7335 19128 7380 19156
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 9677 19159 9735 19165
rect 9677 19125 9689 19159
rect 9723 19156 9735 19159
rect 9858 19156 9864 19168
rect 9723 19128 9864 19156
rect 9723 19125 9735 19128
rect 9677 19119 9735 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 11698 19116 11704 19168
rect 11756 19156 11762 19168
rect 12268 19156 12296 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13464 19224 13492 19332
rect 13538 19320 13544 19372
rect 13596 19360 13602 19372
rect 15013 19363 15071 19369
rect 15013 19360 15025 19363
rect 13596 19332 15025 19360
rect 13596 19320 13602 19332
rect 15013 19329 15025 19332
rect 15059 19329 15071 19363
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15013 19323 15071 19329
rect 15120 19332 15945 19360
rect 13630 19252 13636 19304
rect 13688 19292 13694 19304
rect 13725 19295 13783 19301
rect 13725 19292 13737 19295
rect 13688 19264 13737 19292
rect 13688 19252 13694 19264
rect 13725 19261 13737 19264
rect 13771 19261 13783 19295
rect 13906 19292 13912 19304
rect 13867 19264 13912 19292
rect 13725 19255 13783 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 15120 19224 15148 19332
rect 15933 19329 15945 19332
rect 15979 19360 15991 19363
rect 17402 19360 17408 19372
rect 15979 19332 17408 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19360 17555 19363
rect 17586 19360 17592 19372
rect 17543 19332 17592 19360
rect 17543 19329 17555 19332
rect 17497 19323 17555 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18141 19363 18199 19369
rect 18141 19360 18153 19363
rect 18012 19332 18153 19360
rect 18012 19320 18018 19332
rect 18141 19329 18153 19332
rect 18187 19329 18199 19363
rect 18141 19323 18199 19329
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19360 20407 19363
rect 20806 19360 20812 19372
rect 20395 19332 20812 19360
rect 20395 19329 20407 19332
rect 20349 19323 20407 19329
rect 20806 19320 20812 19332
rect 20864 19360 20870 19372
rect 21450 19360 21456 19372
rect 20864 19332 21456 19360
rect 20864 19320 20870 19332
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 21634 19320 21640 19372
rect 21692 19360 21698 19372
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 21692 19332 22385 19360
rect 21692 19320 21698 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 23750 19320 23756 19372
rect 23808 19320 23814 19372
rect 24670 19320 24676 19372
rect 24728 19360 24734 19372
rect 24765 19363 24823 19369
rect 24765 19360 24777 19363
rect 24728 19332 24777 19360
rect 24728 19320 24734 19332
rect 24765 19329 24777 19332
rect 24811 19329 24823 19363
rect 24765 19323 24823 19329
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19292 16911 19295
rect 16942 19292 16948 19304
rect 16899 19264 16948 19292
rect 16899 19261 16911 19264
rect 16853 19255 16911 19261
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19292 18475 19295
rect 19978 19292 19984 19304
rect 18463 19264 19984 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 23198 19292 23204 19304
rect 22066 19264 23204 19292
rect 22066 19224 22094 19264
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 23290 19252 23296 19304
rect 23348 19292 23354 19304
rect 25038 19292 25044 19304
rect 23348 19264 25044 19292
rect 23348 19252 23354 19264
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 27614 19224 27620 19236
rect 13464 19196 15148 19224
rect 19444 19196 22094 19224
rect 26068 19196 27620 19224
rect 11756 19128 12296 19156
rect 11756 19116 11762 19128
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 19444 19156 19472 19196
rect 19886 19156 19892 19168
rect 16356 19128 19472 19156
rect 19847 19128 19892 19156
rect 16356 19116 16362 19128
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 20438 19156 20444 19168
rect 20399 19128 20444 19156
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 22830 19156 22836 19168
rect 20772 19128 22836 19156
rect 20772 19116 20778 19128
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 23198 19116 23204 19168
rect 23256 19156 23262 19168
rect 26068 19156 26096 19196
rect 27614 19184 27620 19196
rect 27672 19184 27678 19236
rect 23256 19128 26096 19156
rect 23256 19116 23262 19128
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 10410 18952 10416 18964
rect 9999 18924 10416 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 17773 18955 17831 18961
rect 17773 18921 17785 18955
rect 17819 18952 17831 18955
rect 22830 18952 22836 18964
rect 17819 18924 22692 18952
rect 22791 18924 22836 18952
rect 17819 18921 17831 18924
rect 17773 18915 17831 18921
rect 6730 18844 6736 18896
rect 6788 18884 6794 18896
rect 17954 18884 17960 18896
rect 6788 18856 17960 18884
rect 6788 18844 6794 18856
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 7147 18788 8493 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 8481 18785 8493 18788
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 6822 18748 6828 18760
rect 1627 18720 6828 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 6917 18751 6975 18757
rect 6917 18717 6929 18751
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 8588 18748 8616 18856
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 19058 18844 19064 18896
rect 19116 18884 19122 18896
rect 22664 18884 22692 18924
rect 22830 18912 22836 18924
rect 22888 18912 22894 18964
rect 26234 18952 26240 18964
rect 22940 18924 26240 18952
rect 22940 18884 22968 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 27982 18912 27988 18964
rect 28040 18952 28046 18964
rect 28169 18955 28227 18961
rect 28169 18952 28181 18955
rect 28040 18924 28181 18952
rect 28040 18912 28046 18924
rect 28169 18921 28181 18924
rect 28215 18921 28227 18955
rect 28169 18915 28227 18921
rect 19116 18856 21220 18884
rect 22664 18856 22968 18884
rect 19116 18844 19122 18856
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 9272 18788 9505 18816
rect 9272 18776 9278 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 10376 18788 11621 18816
rect 10376 18776 10382 18788
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18816 12311 18819
rect 13262 18816 13268 18828
rect 12299 18788 13268 18816
rect 12299 18785 12311 18788
rect 12253 18779 12311 18785
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 14366 18776 14372 18828
rect 14424 18816 14430 18828
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 14424 18788 14841 18816
rect 14424 18776 14430 18788
rect 14829 18785 14841 18788
rect 14875 18785 14887 18819
rect 15930 18816 15936 18828
rect 15891 18788 15936 18816
rect 14829 18779 14887 18785
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 18966 18816 18972 18828
rect 16040 18788 18972 18816
rect 9306 18748 9312 18760
rect 8435 18720 8616 18748
rect 9267 18720 9312 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 6932 18680 6960 18711
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 11790 18748 11796 18760
rect 11751 18720 11796 18748
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 11940 18720 13185 18748
rect 11940 18708 11946 18720
rect 13173 18717 13185 18720
rect 13219 18748 13231 18751
rect 14550 18748 14556 18760
rect 13219 18720 14556 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 16040 18748 16068 18788
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19242 18776 19248 18828
rect 19300 18816 19306 18828
rect 21085 18819 21143 18825
rect 21085 18816 21097 18819
rect 19300 18788 21097 18816
rect 19300 18776 19306 18788
rect 21085 18785 21097 18788
rect 21131 18785 21143 18819
rect 21192 18816 21220 18856
rect 23382 18844 23388 18896
rect 23440 18884 23446 18896
rect 23440 18856 24716 18884
rect 23440 18844 23446 18856
rect 24578 18816 24584 18828
rect 21192 18788 22968 18816
rect 24539 18788 24584 18816
rect 21085 18779 21143 18785
rect 15528 18720 16068 18748
rect 16117 18751 16175 18757
rect 15528 18708 15534 18720
rect 16117 18717 16129 18751
rect 16163 18717 16175 18751
rect 16117 18711 16175 18717
rect 7098 18680 7104 18692
rect 6932 18652 7104 18680
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 14921 18683 14979 18689
rect 14921 18680 14933 18683
rect 13688 18652 14933 18680
rect 13688 18640 13694 18652
rect 14921 18649 14933 18652
rect 14967 18649 14979 18683
rect 14921 18643 14979 18649
rect 15562 18640 15568 18692
rect 15620 18680 15626 18692
rect 16132 18680 16160 18711
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 16264 18720 17049 18748
rect 16264 18708 16270 18720
rect 17037 18717 17049 18720
rect 17083 18748 17095 18751
rect 17681 18751 17739 18757
rect 17083 18720 17632 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 15620 18652 16160 18680
rect 15620 18640 15626 18652
rect 1762 18612 1768 18624
rect 1723 18584 1768 18612
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 7561 18615 7619 18621
rect 7561 18581 7573 18615
rect 7607 18612 7619 18615
rect 8294 18612 8300 18624
rect 7607 18584 8300 18612
rect 7607 18581 7619 18584
rect 7561 18575 7619 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 10965 18615 11023 18621
rect 10965 18581 10977 18615
rect 11011 18612 11023 18615
rect 12250 18612 12256 18624
rect 11011 18584 12256 18612
rect 11011 18581 11023 18584
rect 10965 18575 11023 18581
rect 12250 18572 12256 18584
rect 12308 18572 12314 18624
rect 13265 18615 13323 18621
rect 13265 18581 13277 18615
rect 13311 18612 13323 18615
rect 14458 18612 14464 18624
rect 13311 18584 14464 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 16206 18572 16212 18624
rect 16264 18612 16270 18624
rect 16577 18615 16635 18621
rect 16577 18612 16589 18615
rect 16264 18584 16589 18612
rect 16264 18572 16270 18584
rect 16577 18581 16589 18584
rect 16623 18581 16635 18615
rect 16577 18575 16635 18581
rect 17129 18615 17187 18621
rect 17129 18581 17141 18615
rect 17175 18612 17187 18615
rect 17402 18612 17408 18624
rect 17175 18584 17408 18612
rect 17175 18581 17187 18584
rect 17129 18575 17187 18581
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 17604 18612 17632 18720
rect 17681 18717 17693 18751
rect 17727 18748 17739 18751
rect 18138 18748 18144 18760
rect 17727 18720 18144 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 18138 18708 18144 18720
rect 18196 18748 18202 18760
rect 18317 18753 18375 18759
rect 18317 18750 18329 18753
rect 18248 18748 18329 18750
rect 18196 18722 18329 18748
rect 18196 18720 18276 18722
rect 18196 18708 18202 18720
rect 18317 18719 18329 18722
rect 18363 18719 18375 18753
rect 18317 18713 18375 18719
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 20898 18748 20904 18760
rect 18472 18720 20904 18748
rect 18472 18708 18478 18720
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 19886 18680 19892 18692
rect 17920 18652 19892 18680
rect 17920 18640 17926 18652
rect 19886 18640 19892 18652
rect 19944 18640 19950 18692
rect 21266 18640 21272 18692
rect 21324 18680 21330 18692
rect 21361 18683 21419 18689
rect 21361 18680 21373 18683
rect 21324 18652 21373 18680
rect 21324 18640 21330 18652
rect 21361 18649 21373 18652
rect 21407 18649 21419 18683
rect 22830 18680 22836 18692
rect 22586 18652 22836 18680
rect 21361 18643 21419 18649
rect 22830 18640 22836 18652
rect 22888 18640 22894 18692
rect 22940 18680 22968 18788
rect 24578 18776 24584 18788
rect 24636 18776 24642 18828
rect 24688 18816 24716 18856
rect 26510 18844 26516 18896
rect 26568 18884 26574 18896
rect 27062 18884 27068 18896
rect 26568 18856 27068 18884
rect 26568 18844 26574 18856
rect 27062 18844 27068 18856
rect 27120 18844 27126 18896
rect 26605 18819 26663 18825
rect 26605 18816 26617 18819
rect 24688 18788 26617 18816
rect 26605 18785 26617 18788
rect 26651 18785 26663 18819
rect 26605 18779 26663 18785
rect 28353 18751 28411 18757
rect 28353 18717 28365 18751
rect 28399 18748 28411 18751
rect 29914 18748 29920 18760
rect 28399 18720 29920 18748
rect 28399 18717 28411 18720
rect 28353 18711 28411 18717
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 22940 18652 23244 18680
rect 18322 18612 18328 18624
rect 17604 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 23106 18612 23112 18624
rect 18463 18584 23112 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 23106 18572 23112 18584
rect 23164 18572 23170 18624
rect 23216 18612 23244 18652
rect 24210 18640 24216 18692
rect 24268 18680 24274 18692
rect 24857 18683 24915 18689
rect 24857 18680 24869 18683
rect 24268 18652 24869 18680
rect 24268 18640 24274 18652
rect 24857 18649 24869 18652
rect 24903 18649 24915 18683
rect 24857 18643 24915 18649
rect 25043 18652 25346 18680
rect 25043 18612 25071 18652
rect 23216 18584 25071 18612
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 8294 18408 8300 18420
rect 8255 18380 8300 18408
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 13725 18411 13783 18417
rect 12216 18380 13676 18408
rect 12216 18368 12222 18380
rect 6730 18340 6736 18352
rect 4448 18312 6736 18340
rect 4448 18281 4476 18312
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 10888 18312 12434 18340
rect 10888 18284 10916 18312
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18241 5319 18275
rect 5261 18235 5319 18241
rect 5276 18204 5304 18235
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7432 18244 7849 18272
rect 7432 18232 7438 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 8444 18244 9229 18272
rect 8444 18232 8450 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9217 18235 9275 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18272 10563 18275
rect 10870 18272 10876 18284
rect 10551 18244 10876 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11882 18272 11888 18284
rect 11195 18244 11888 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12250 18272 12256 18284
rect 12211 18244 12256 18272
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 12406 18272 12434 18312
rect 13648 18281 13676 18380
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 13906 18408 13912 18420
rect 13771 18380 13912 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 15473 18411 15531 18417
rect 15473 18377 15485 18411
rect 15519 18408 15531 18411
rect 15562 18408 15568 18420
rect 15519 18380 15568 18408
rect 15519 18377 15531 18380
rect 15473 18371 15531 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 19518 18408 19524 18420
rect 16224 18380 19524 18408
rect 14458 18340 14464 18352
rect 14419 18312 14464 18340
rect 14458 18300 14464 18312
rect 14516 18300 14522 18352
rect 14550 18300 14556 18352
rect 14608 18340 14614 18352
rect 16224 18340 16252 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 19978 18408 19984 18420
rect 19939 18380 19984 18408
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20438 18368 20444 18420
rect 20496 18408 20502 18420
rect 23198 18408 23204 18420
rect 20496 18380 23204 18408
rect 20496 18368 20502 18380
rect 23198 18368 23204 18380
rect 23256 18368 23262 18420
rect 23566 18368 23572 18420
rect 23624 18408 23630 18420
rect 25130 18408 25136 18420
rect 23624 18380 25136 18408
rect 23624 18368 23630 18380
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 16942 18340 16948 18352
rect 14608 18312 16252 18340
rect 16903 18312 16948 18340
rect 14608 18300 14614 18312
rect 16942 18300 16948 18312
rect 17000 18300 17006 18352
rect 17034 18300 17040 18352
rect 17092 18340 17098 18352
rect 17092 18312 17137 18340
rect 17092 18300 17098 18312
rect 17402 18300 17408 18352
rect 17460 18340 17466 18352
rect 17460 18312 18998 18340
rect 17460 18300 17466 18312
rect 19886 18300 19892 18352
rect 19944 18340 19950 18352
rect 25593 18343 25651 18349
rect 19944 18312 24334 18340
rect 19944 18300 19950 18312
rect 25593 18309 25605 18343
rect 25639 18340 25651 18343
rect 25866 18340 25872 18352
rect 25639 18312 25872 18340
rect 25639 18309 25651 18312
rect 25593 18303 25651 18309
rect 25866 18300 25872 18312
rect 25924 18300 25930 18352
rect 13633 18275 13691 18281
rect 12406 18244 13584 18272
rect 4264 18176 5304 18204
rect 4264 18145 4292 18176
rect 7466 18164 7472 18216
rect 7524 18204 7530 18216
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7524 18176 7665 18204
rect 7524 18164 7530 18176
rect 7653 18173 7665 18176
rect 7699 18204 7711 18207
rect 8570 18204 8576 18216
rect 7699 18176 8576 18204
rect 7699 18173 7711 18176
rect 7653 18167 7711 18173
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 11112 18176 12449 18204
rect 11112 18164 11118 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 4249 18139 4307 18145
rect 4249 18105 4261 18139
rect 4295 18105 4307 18139
rect 4249 18099 4307 18105
rect 9033 18139 9091 18145
rect 9033 18105 9045 18139
rect 9079 18136 9091 18139
rect 9858 18136 9864 18148
rect 9079 18108 9864 18136
rect 9079 18105 9091 18108
rect 9033 18099 9091 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 10321 18139 10379 18145
rect 10321 18105 10333 18139
rect 10367 18136 10379 18139
rect 11882 18136 11888 18148
rect 10367 18108 11888 18136
rect 10367 18105 10379 18108
rect 10321 18099 10379 18105
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 13556 18136 13584 18244
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 13906 18272 13912 18284
rect 13679 18244 13912 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 13906 18232 13912 18244
rect 13964 18232 13970 18284
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18272 15071 18275
rect 15470 18272 15476 18284
rect 15059 18244 15476 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 15654 18272 15660 18284
rect 15615 18244 15660 18272
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16114 18272 16120 18284
rect 15988 18244 16120 18272
rect 15988 18232 15994 18244
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 16209 18275 16267 18281
rect 16209 18241 16221 18275
rect 16255 18272 16267 18275
rect 16298 18272 16304 18284
rect 16255 18244 16304 18272
rect 16255 18241 16267 18244
rect 16209 18235 16267 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 14366 18204 14372 18216
rect 14327 18176 14372 18204
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 17218 18204 17224 18216
rect 14476 18176 16344 18204
rect 17179 18176 17224 18204
rect 14476 18136 14504 18176
rect 13556 18108 14504 18136
rect 5077 18071 5135 18077
rect 5077 18037 5089 18071
rect 5123 18068 5135 18071
rect 5534 18068 5540 18080
rect 5123 18040 5540 18068
rect 5123 18037 5135 18040
rect 5077 18031 5135 18037
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 10965 18071 11023 18077
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 11974 18068 11980 18080
rect 11011 18040 11980 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 16316 18068 16344 18176
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 18046 18164 18052 18216
rect 18104 18204 18110 18216
rect 18233 18207 18291 18213
rect 18233 18204 18245 18207
rect 18104 18176 18245 18204
rect 18104 18164 18110 18176
rect 18233 18173 18245 18176
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 18874 18204 18880 18216
rect 18555 18176 18880 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 23569 18207 23627 18213
rect 23569 18173 23581 18207
rect 23615 18204 23627 18207
rect 23845 18207 23903 18213
rect 23615 18176 23704 18204
rect 23615 18173 23627 18176
rect 23569 18167 23627 18173
rect 23290 18136 23296 18148
rect 19536 18108 23296 18136
rect 19536 18068 19564 18108
rect 23290 18096 23296 18108
rect 23348 18096 23354 18148
rect 16316 18040 19564 18068
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 23566 18068 23572 18080
rect 19668 18040 23572 18068
rect 19668 18028 19674 18040
rect 23566 18028 23572 18040
rect 23624 18028 23630 18080
rect 23676 18068 23704 18176
rect 23845 18173 23857 18207
rect 23891 18204 23903 18207
rect 23934 18204 23940 18216
rect 23891 18176 23940 18204
rect 23891 18173 23903 18176
rect 23845 18167 23903 18173
rect 23934 18164 23940 18176
rect 23992 18164 23998 18216
rect 24578 18068 24584 18080
rect 23676 18040 24584 18068
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 6822 17824 6828 17876
rect 6880 17864 6886 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 6880 17836 7757 17864
rect 6880 17824 6886 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 8386 17864 8392 17876
rect 8347 17836 8392 17864
rect 7745 17827 7803 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9306 17864 9312 17876
rect 9267 17836 9312 17864
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 11793 17867 11851 17873
rect 9456 17836 10180 17864
rect 9456 17824 9462 17836
rect 9398 17728 9404 17740
rect 8588 17700 9404 17728
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 5350 17484 5356 17536
rect 5408 17524 5414 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5408 17496 5825 17524
rect 5408 17484 5414 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 7944 17524 7972 17623
rect 8386 17620 8392 17672
rect 8444 17660 8450 17672
rect 8588 17669 8616 17700
rect 9398 17688 9404 17700
rect 9456 17688 9462 17740
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9732 17700 10057 17728
rect 9732 17688 9738 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10152 17728 10180 17836
rect 11793 17833 11805 17867
rect 11839 17864 11851 17867
rect 13630 17864 13636 17876
rect 11839 17836 13636 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 24302 17864 24308 17876
rect 13740 17836 24308 17864
rect 13740 17728 13768 17836
rect 24302 17824 24308 17836
rect 24360 17824 24366 17876
rect 24394 17824 24400 17876
rect 24452 17864 24458 17876
rect 27065 17867 27123 17873
rect 27065 17864 27077 17867
rect 24452 17836 27077 17864
rect 24452 17824 24458 17836
rect 27065 17833 27077 17836
rect 27111 17833 27123 17867
rect 27065 17827 27123 17833
rect 15194 17796 15200 17808
rect 15155 17768 15200 17796
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 15933 17799 15991 17805
rect 15933 17765 15945 17799
rect 15979 17796 15991 17799
rect 17034 17796 17040 17808
rect 15979 17768 17040 17796
rect 15979 17765 15991 17768
rect 15933 17759 15991 17765
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 17954 17756 17960 17808
rect 18012 17796 18018 17808
rect 18012 17768 19564 17796
rect 18012 17756 18018 17768
rect 10152 17700 13768 17728
rect 10045 17691 10103 17697
rect 15838 17688 15844 17740
rect 15896 17728 15902 17740
rect 15896 17700 17724 17728
rect 15896 17688 15902 17700
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 8444 17632 8585 17660
rect 8444 17620 8450 17632
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 9214 17660 9220 17672
rect 9175 17632 9220 17660
rect 8573 17623 8631 17629
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17660 9919 17663
rect 10060 17660 10180 17662
rect 11238 17660 11244 17672
rect 9907 17634 11244 17660
rect 9907 17632 10088 17634
rect 10152 17632 11244 17634
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17629 11391 17663
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11333 17623 11391 17629
rect 10505 17595 10563 17601
rect 10505 17561 10517 17595
rect 10551 17592 10563 17595
rect 11054 17592 11060 17604
rect 10551 17564 11060 17592
rect 10551 17561 10563 17564
rect 10505 17555 10563 17561
rect 11054 17552 11060 17564
rect 11112 17552 11118 17604
rect 10962 17524 10968 17536
rect 7944 17496 10968 17524
rect 5813 17487 5871 17493
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11146 17524 11152 17536
rect 11107 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 11348 17524 11376 17623
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12400 17632 12633 17660
rect 12400 17620 12406 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 12894 17620 12900 17672
rect 12952 17660 12958 17672
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12952 17632 13093 17660
rect 12952 17620 12958 17632
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17629 13323 17663
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13265 17623 13323 17629
rect 12986 17552 12992 17604
rect 13044 17592 13050 17604
rect 13280 17592 13308 17623
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14332 17632 14841 17660
rect 14332 17620 14338 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17629 15071 17663
rect 16114 17660 16120 17672
rect 16075 17632 16120 17660
rect 15013 17623 15071 17629
rect 15028 17592 15056 17623
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 16574 17660 16580 17672
rect 16535 17632 16580 17660
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17586 17660 17592 17672
rect 17543 17632 17592 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 17696 17660 17724 17700
rect 18046 17688 18052 17740
rect 18104 17728 18110 17740
rect 18690 17728 18696 17740
rect 18104 17700 18696 17728
rect 18104 17688 18110 17700
rect 18690 17688 18696 17700
rect 18748 17728 18754 17740
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 18748 17700 19441 17728
rect 18748 17688 18754 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19536 17728 19564 17768
rect 20732 17768 21772 17796
rect 20732 17728 20760 17768
rect 21634 17728 21640 17740
rect 19536 17700 20760 17728
rect 21595 17700 21640 17728
rect 19429 17691 19487 17697
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 21744 17728 21772 17768
rect 24946 17756 24952 17808
rect 25004 17796 25010 17808
rect 25041 17799 25099 17805
rect 25041 17796 25053 17799
rect 25004 17768 25053 17796
rect 25004 17756 25010 17768
rect 25041 17765 25053 17768
rect 25087 17796 25099 17799
rect 25087 17768 25452 17796
rect 25087 17765 25099 17768
rect 25041 17759 25099 17765
rect 24486 17728 24492 17740
rect 21744 17700 24492 17728
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 24578 17688 24584 17740
rect 24636 17728 24642 17740
rect 25317 17731 25375 17737
rect 25317 17728 25329 17731
rect 24636 17700 25329 17728
rect 24636 17688 24642 17700
rect 25317 17697 25329 17700
rect 25363 17697 25375 17731
rect 25424 17728 25452 17768
rect 25593 17731 25651 17737
rect 25593 17728 25605 17731
rect 25424 17700 25605 17728
rect 25317 17691 25375 17697
rect 25593 17697 25605 17700
rect 25639 17728 25651 17731
rect 27890 17728 27896 17740
rect 25639 17700 27896 17728
rect 25639 17697 25651 17700
rect 25593 17691 25651 17697
rect 27890 17688 27896 17700
rect 27948 17688 27954 17740
rect 18141 17663 18199 17669
rect 17696 17632 18092 17660
rect 13044 17564 13308 17592
rect 13648 17564 15056 17592
rect 16853 17595 16911 17601
rect 13044 17552 13050 17564
rect 11974 17524 11980 17536
rect 11348 17496 11980 17524
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12437 17527 12495 17533
rect 12437 17493 12449 17527
rect 12483 17524 12495 17527
rect 13648 17524 13676 17564
rect 16853 17561 16865 17595
rect 16899 17592 16911 17595
rect 17954 17592 17960 17604
rect 16899 17564 17960 17592
rect 16899 17561 16911 17564
rect 16853 17555 16911 17561
rect 17954 17552 17960 17564
rect 18012 17552 18018 17604
rect 17586 17524 17592 17536
rect 12483 17496 13676 17524
rect 17547 17496 17592 17524
rect 12483 17493 12495 17496
rect 12437 17487 12495 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 18064 17524 18092 17632
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 18230 17660 18236 17672
rect 18187 17632 18236 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18156 17592 18184 17623
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 18156 17564 19717 17592
rect 19705 17561 19717 17564
rect 19751 17592 19763 17595
rect 19751 17564 20024 17592
rect 20930 17564 21312 17592
rect 19751 17561 19763 17564
rect 19705 17555 19763 17561
rect 18233 17527 18291 17533
rect 18233 17524 18245 17527
rect 18064 17496 18245 17524
rect 18233 17493 18245 17496
rect 18279 17493 18291 17527
rect 18233 17487 18291 17493
rect 18782 17484 18788 17536
rect 18840 17524 18846 17536
rect 19886 17524 19892 17536
rect 18840 17496 19892 17524
rect 18840 17484 18846 17496
rect 19886 17484 19892 17496
rect 19944 17484 19950 17536
rect 19996 17524 20024 17564
rect 20622 17524 20628 17536
rect 19996 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 21284 17524 21312 17564
rect 21542 17552 21548 17604
rect 21600 17592 21606 17604
rect 21913 17595 21971 17601
rect 21913 17592 21925 17595
rect 21600 17564 21925 17592
rect 21600 17552 21606 17564
rect 21913 17561 21925 17564
rect 21959 17592 21971 17595
rect 22002 17592 22008 17604
rect 21959 17564 22008 17592
rect 21959 17561 21971 17564
rect 21913 17555 21971 17561
rect 22002 17552 22008 17564
rect 22060 17552 22066 17604
rect 22370 17552 22376 17604
rect 22428 17552 22434 17604
rect 23566 17592 23572 17604
rect 23216 17564 23572 17592
rect 23216 17524 23244 17564
rect 23566 17552 23572 17564
rect 23624 17552 23630 17604
rect 26234 17552 26240 17604
rect 26292 17552 26298 17604
rect 23382 17524 23388 17536
rect 21284 17496 23244 17524
rect 23343 17496 23388 17524
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 24302 17484 24308 17536
rect 24360 17524 24366 17536
rect 28166 17524 28172 17536
rect 24360 17496 28172 17524
rect 24360 17484 24366 17496
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17289 6699 17323
rect 6641 17283 6699 17289
rect 6656 17252 6684 17283
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 10965 17323 11023 17329
rect 6972 17292 8708 17320
rect 6972 17280 6978 17292
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 6656 17224 7481 17252
rect 7469 17221 7481 17224
rect 7515 17221 7527 17255
rect 7469 17215 7527 17221
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 8680 17261 8708 17292
rect 10965 17289 10977 17323
rect 11011 17320 11023 17323
rect 11790 17320 11796 17332
rect 11011 17292 11796 17320
rect 11011 17289 11023 17292
rect 10965 17283 11023 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12342 17320 12348 17332
rect 12303 17292 12348 17320
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 13354 17320 13360 17332
rect 13096 17292 13360 17320
rect 13096 17261 13124 17292
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 16022 17320 16028 17332
rect 15488 17292 16028 17320
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 8352 17224 8585 17252
rect 8352 17212 8358 17224
rect 8573 17221 8585 17224
rect 8619 17221 8631 17255
rect 8573 17215 8631 17221
rect 8665 17255 8723 17261
rect 8665 17221 8677 17255
rect 8711 17221 8723 17255
rect 13081 17255 13139 17261
rect 8665 17215 8723 17221
rect 10336 17224 12664 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 5166 17184 5172 17196
rect 1627 17156 5172 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5350 17184 5356 17196
rect 5311 17156 5356 17184
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5534 17184 5540 17196
rect 5495 17156 5540 17184
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7190 17184 7196 17196
rect 6871 17156 7196 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 10336 17193 10364 17224
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17153 10379 17187
rect 11146 17184 11152 17196
rect 11107 17156 11152 17184
rect 10321 17147 10379 17153
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 11882 17184 11888 17196
rect 11843 17156 11888 17184
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 12526 17184 12532 17196
rect 12487 17156 12532 17184
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12636 17184 12664 17224
rect 13081 17221 13093 17255
rect 13127 17221 13139 17255
rect 13081 17215 13139 17221
rect 13182 17255 13240 17261
rect 13182 17221 13194 17255
rect 13228 17252 13240 17255
rect 13446 17252 13452 17264
rect 13228 17224 13452 17252
rect 13228 17221 13240 17224
rect 13182 17215 13240 17221
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 15488 17261 15516 17292
rect 16022 17280 16028 17292
rect 16080 17320 16086 17332
rect 16080 17292 17448 17320
rect 16080 17280 16086 17292
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 14240 17224 14933 17252
rect 14240 17212 14246 17224
rect 14921 17221 14933 17224
rect 14967 17221 14979 17255
rect 14921 17215 14979 17221
rect 15473 17255 15531 17261
rect 15473 17221 15485 17255
rect 15519 17221 15531 17255
rect 17126 17252 17132 17264
rect 15473 17215 15531 17221
rect 16132 17224 17132 17252
rect 16132 17193 16160 17224
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 17420 17252 17448 17292
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17644 17292 19840 17320
rect 17644 17280 17650 17292
rect 18598 17252 18604 17264
rect 17420 17224 18604 17252
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 19812 17252 19840 17292
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20622 17320 20628 17332
rect 20220 17292 20628 17320
rect 20220 17280 20226 17292
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 21358 17320 21364 17332
rect 20772 17292 21364 17320
rect 20772 17280 20778 17292
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 21450 17280 21456 17332
rect 21508 17320 21514 17332
rect 21818 17320 21824 17332
rect 21508 17292 21824 17320
rect 21508 17280 21514 17292
rect 21818 17280 21824 17292
rect 21876 17320 21882 17332
rect 26513 17323 26571 17329
rect 26513 17320 26525 17323
rect 21876 17292 26525 17320
rect 21876 17280 21882 17292
rect 26513 17289 26525 17292
rect 26559 17289 26571 17323
rect 26513 17283 26571 17289
rect 19812 17224 23322 17252
rect 25130 17212 25136 17264
rect 25188 17252 25194 17264
rect 25188 17224 25530 17252
rect 25188 17212 25194 17224
rect 16117 17187 16175 17193
rect 12636 17156 12848 17184
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 5736 17088 7389 17116
rect 5736 17060 5764 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 7524 17088 7665 17116
rect 7524 17076 7530 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 1762 17048 1768 17060
rect 1723 17020 1768 17048
rect 1762 17008 1768 17020
rect 1820 17008 1826 17060
rect 5718 17048 5724 17060
rect 5679 17020 5724 17048
rect 5718 17008 5724 17020
rect 5776 17008 5782 17060
rect 7668 17048 7696 17079
rect 8018 17076 8024 17128
rect 8076 17116 8082 17128
rect 12618 17116 12624 17128
rect 8076 17088 12624 17116
rect 8076 17076 8082 17088
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 12820 17116 12848 17156
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16632 17156 16865 17184
rect 16632 17144 16638 17156
rect 16853 17153 16865 17156
rect 16899 17184 16911 17187
rect 17402 17184 17408 17196
rect 16899 17156 17408 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17402 17144 17408 17156
rect 17460 17144 17466 17196
rect 18046 17184 18052 17196
rect 18007 17156 18052 17184
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 20257 17187 20315 17193
rect 13354 17116 13360 17128
rect 12820 17088 13124 17116
rect 13315 17088 13360 17116
rect 9125 17051 9183 17057
rect 9125 17048 9137 17051
rect 7668 17020 9137 17048
rect 9125 17017 9137 17020
rect 9171 17017 9183 17051
rect 9125 17011 9183 17017
rect 10137 17051 10195 17057
rect 10137 17017 10149 17051
rect 10183 17048 10195 17051
rect 11238 17048 11244 17060
rect 10183 17020 11244 17048
rect 10183 17017 10195 17020
rect 10137 17011 10195 17017
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 11701 17051 11759 17057
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 12986 17048 12992 17060
rect 11747 17020 12992 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 12986 17008 12992 17020
rect 13044 17008 13050 17060
rect 13096 17048 13124 17088
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 17862 17116 17868 17128
rect 17175 17088 17868 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 14550 17048 14556 17060
rect 13096 17020 14556 17048
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 14844 17048 14872 17079
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 18325 17119 18383 17125
rect 18325 17085 18337 17119
rect 18371 17116 18383 17119
rect 19444 17116 19472 17170
rect 20257 17153 20269 17187
rect 20303 17184 20315 17187
rect 20806 17184 20812 17196
rect 20303 17156 20812 17184
rect 20303 17153 20315 17156
rect 20257 17147 20315 17153
rect 20806 17144 20812 17156
rect 20864 17184 20870 17196
rect 21082 17184 21088 17196
rect 20864 17156 21088 17184
rect 20864 17144 20870 17156
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 21634 17144 21640 17196
rect 21692 17184 21698 17196
rect 22557 17187 22615 17193
rect 22557 17184 22569 17187
rect 21692 17156 22569 17184
rect 21692 17144 21698 17156
rect 22557 17153 22569 17156
rect 22603 17153 22615 17187
rect 22557 17147 22615 17153
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 24765 17187 24823 17193
rect 24765 17184 24777 17187
rect 24636 17156 24777 17184
rect 24636 17144 24642 17156
rect 24765 17153 24777 17156
rect 24811 17153 24823 17187
rect 28350 17184 28356 17196
rect 28311 17156 28356 17184
rect 24765 17147 24823 17153
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 22278 17116 22284 17128
rect 18371 17088 19380 17116
rect 19444 17088 22284 17116
rect 18371 17085 18383 17088
rect 18325 17079 18383 17085
rect 14792 17020 14872 17048
rect 19352 17048 19380 17088
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 22462 17076 22468 17128
rect 22520 17116 22526 17128
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 22520 17088 22845 17116
rect 22520 17076 22526 17088
rect 22833 17085 22845 17088
rect 22879 17085 22891 17119
rect 22833 17079 22891 17085
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 24176 17088 24317 17116
rect 24176 17076 24182 17088
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 24305 17079 24363 17085
rect 24486 17076 24492 17128
rect 24544 17116 24550 17128
rect 25041 17119 25099 17125
rect 25041 17116 25053 17119
rect 24544 17088 25053 17116
rect 24544 17076 24550 17088
rect 25041 17085 25053 17088
rect 25087 17116 25099 17119
rect 26694 17116 26700 17128
rect 25087 17088 26700 17116
rect 25087 17085 25099 17088
rect 25041 17079 25099 17085
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 21910 17048 21916 17060
rect 19352 17020 21916 17048
rect 14792 17008 14798 17020
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 22002 17008 22008 17060
rect 22060 17048 22066 17060
rect 22060 17020 22692 17048
rect 22060 17008 22066 17020
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 19702 16980 19708 16992
rect 16255 16952 19708 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 19886 16980 19892 16992
rect 19843 16952 19892 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 22554 16980 22560 16992
rect 20395 16952 22560 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 22664 16980 22692 17020
rect 24026 16980 24032 16992
rect 22664 16952 24032 16980
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 27982 16940 27988 16992
rect 28040 16980 28046 16992
rect 28169 16983 28227 16989
rect 28169 16980 28181 16983
rect 28040 16952 28181 16980
rect 28040 16940 28046 16952
rect 28169 16949 28181 16952
rect 28215 16949 28227 16983
rect 28169 16943 28227 16949
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 5224 16748 5457 16776
rect 5224 16736 5230 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 5445 16739 5503 16745
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7745 16779 7803 16785
rect 7745 16776 7757 16779
rect 7248 16748 7757 16776
rect 7248 16736 7254 16748
rect 7745 16745 7757 16748
rect 7791 16745 7803 16779
rect 12526 16776 12532 16788
rect 7745 16739 7803 16745
rect 8404 16748 12532 16776
rect 3970 16668 3976 16720
rect 4028 16708 4034 16720
rect 7006 16708 7012 16720
rect 4028 16680 7012 16708
rect 4028 16668 4034 16680
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 6288 16612 7972 16640
rect 6288 16581 6316 16612
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 7006 16572 7012 16584
rect 6967 16544 7012 16572
rect 6273 16535 6331 16541
rect 5644 16504 5672 16535
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7098 16532 7104 16584
rect 7156 16572 7162 16584
rect 7944 16581 7972 16612
rect 7929 16575 7987 16581
rect 7156 16544 7201 16572
rect 7156 16532 7162 16544
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8018 16572 8024 16584
rect 7975 16544 8024 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 8404 16581 8432 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 21450 16776 21456 16788
rect 12676 16748 21456 16776
rect 12676 16736 12682 16748
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 23382 16776 23388 16788
rect 21744 16748 23388 16776
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 8628 16680 9720 16708
rect 8628 16668 8634 16680
rect 9692 16649 9720 16680
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 11756 16680 12940 16708
rect 11756 16668 11762 16680
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9858 16640 9864 16652
rect 9819 16612 9864 16640
rect 9677 16603 9735 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 12912 16649 12940 16680
rect 14550 16668 14556 16720
rect 14608 16708 14614 16720
rect 18966 16708 18972 16720
rect 14608 16680 18972 16708
rect 14608 16668 14614 16680
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 19334 16668 19340 16720
rect 19392 16708 19398 16720
rect 19392 16680 19564 16708
rect 19392 16668 19398 16680
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12492 16612 12633 16640
rect 12492 16600 12498 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16609 12955 16643
rect 14274 16640 14280 16652
rect 14235 16612 14280 16640
rect 12897 16603 12955 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 15436 16612 15577 16640
rect 15436 16600 15442 16612
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 15838 16640 15844 16652
rect 15795 16612 15844 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 15930 16600 15936 16652
rect 15988 16640 15994 16652
rect 16298 16640 16304 16652
rect 15988 16612 16304 16640
rect 15988 16600 15994 16612
rect 16298 16600 16304 16612
rect 16356 16640 16362 16652
rect 16356 16612 18276 16640
rect 16356 16600 16362 16612
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 11296 16544 11529 16572
rect 11296 16532 11302 16544
rect 11517 16541 11529 16544
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 15105 16575 15163 16581
rect 15105 16541 15117 16575
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16572 17095 16575
rect 17126 16572 17132 16584
rect 17083 16544 17132 16572
rect 17083 16541 17095 16544
rect 17037 16535 17095 16541
rect 8481 16507 8539 16513
rect 8481 16504 8493 16507
rect 5644 16476 8493 16504
rect 8481 16473 8493 16476
rect 8527 16473 8539 16507
rect 8481 16467 8539 16473
rect 12066 16464 12072 16516
rect 12124 16504 12130 16516
rect 12713 16507 12771 16513
rect 12124 16476 12572 16504
rect 12124 16464 12130 16476
rect 6365 16439 6423 16445
rect 6365 16405 6377 16439
rect 6411 16436 6423 16439
rect 6914 16436 6920 16448
rect 6411 16408 6920 16436
rect 6411 16405 6423 16408
rect 6365 16399 6423 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10962 16436 10968 16448
rect 10367 16408 10968 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 11333 16439 11391 16445
rect 11333 16405 11345 16439
rect 11379 16436 11391 16439
rect 12434 16436 12440 16448
rect 11379 16408 12440 16436
rect 11379 16405 11391 16408
rect 11333 16399 11391 16405
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 12544 16436 12572 16476
rect 12713 16473 12725 16507
rect 12759 16473 12771 16507
rect 15120 16504 15148 16535
rect 17126 16532 17132 16544
rect 17184 16572 17190 16584
rect 17586 16572 17592 16584
rect 17184 16544 17592 16572
rect 17184 16532 17190 16544
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 17954 16572 17960 16584
rect 17727 16544 17960 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 17954 16532 17960 16544
rect 18012 16572 18018 16584
rect 18138 16572 18144 16584
rect 18012 16544 18144 16572
rect 18012 16532 18018 16544
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18248 16572 18276 16612
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19429 16643 19487 16649
rect 19429 16640 19441 16643
rect 19300 16612 19441 16640
rect 19300 16600 19306 16612
rect 19429 16609 19441 16612
rect 19475 16609 19487 16643
rect 19536 16640 19564 16680
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 21744 16708 21772 16748
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 20772 16680 21772 16708
rect 20772 16668 20778 16680
rect 19705 16643 19763 16649
rect 19705 16640 19717 16643
rect 19536 16612 19717 16640
rect 19429 16603 19487 16609
rect 19705 16609 19717 16612
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 20070 16600 20076 16652
rect 20128 16640 20134 16652
rect 21634 16640 21640 16652
rect 20128 16612 20944 16640
rect 21595 16612 21640 16640
rect 20128 16600 20134 16612
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18248 16544 18337 16572
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 20916 16572 20944 16612
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 21910 16600 21916 16652
rect 21968 16640 21974 16652
rect 22462 16640 22468 16652
rect 21968 16612 22468 16640
rect 21968 16600 21974 16612
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 23750 16640 23756 16652
rect 22612 16612 23756 16640
rect 22612 16600 22618 16612
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 26329 16643 26387 16649
rect 26329 16640 26341 16643
rect 24636 16612 26341 16640
rect 24636 16600 24642 16612
rect 26329 16609 26341 16612
rect 26375 16609 26387 16643
rect 26602 16640 26608 16652
rect 26563 16612 26608 16640
rect 26329 16603 26387 16609
rect 26602 16600 26608 16612
rect 26660 16600 26666 16652
rect 20916 16544 21680 16572
rect 18325 16535 18383 16541
rect 21652 16516 21680 16544
rect 19610 16504 19616 16516
rect 15120 16476 19616 16504
rect 12713 16467 12771 16473
rect 12728 16436 12756 16467
rect 19610 16464 19616 16476
rect 19668 16464 19674 16516
rect 21266 16504 21272 16516
rect 20930 16476 21272 16504
rect 21266 16464 21272 16476
rect 21324 16464 21330 16516
rect 21634 16464 21640 16516
rect 21692 16464 21698 16516
rect 21818 16464 21824 16516
rect 21876 16504 21882 16516
rect 21913 16507 21971 16513
rect 21913 16504 21925 16507
rect 21876 16476 21925 16504
rect 21876 16464 21882 16476
rect 21913 16473 21925 16476
rect 21959 16473 21971 16507
rect 21913 16467 21971 16473
rect 22370 16464 22376 16516
rect 22428 16464 22434 16516
rect 23198 16464 23204 16516
rect 23256 16504 23262 16516
rect 25130 16504 25136 16516
rect 23256 16476 25136 16504
rect 23256 16464 23262 16476
rect 25130 16464 25136 16476
rect 25188 16464 25194 16516
rect 27614 16464 27620 16516
rect 27672 16464 27678 16516
rect 28074 16464 28080 16516
rect 28132 16504 28138 16516
rect 28353 16507 28411 16513
rect 28353 16504 28365 16507
rect 28132 16476 28365 16504
rect 28132 16464 28138 16476
rect 28353 16473 28365 16476
rect 28399 16473 28411 16507
rect 28353 16467 28411 16473
rect 12544 16408 12756 16436
rect 14921 16439 14979 16445
rect 14921 16405 14933 16439
rect 14967 16436 14979 16439
rect 16114 16436 16120 16448
rect 14967 16408 16120 16436
rect 14967 16405 14979 16408
rect 14921 16399 14979 16405
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 16206 16396 16212 16448
rect 16264 16436 16270 16448
rect 17126 16436 17132 16448
rect 16264 16408 16309 16436
rect 17087 16408 17132 16436
rect 16264 16396 16270 16408
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 17770 16436 17776 16448
rect 17731 16408 17776 16436
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16436 18475 16439
rect 20346 16436 20352 16448
rect 18463 16408 20352 16436
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 20496 16408 21189 16436
rect 20496 16396 20502 16408
rect 21177 16405 21189 16408
rect 21223 16405 21235 16439
rect 21177 16399 21235 16405
rect 21542 16396 21548 16448
rect 21600 16436 21606 16448
rect 23385 16439 23443 16445
rect 23385 16436 23397 16439
rect 21600 16408 23397 16436
rect 21600 16396 21606 16408
rect 23385 16405 23397 16408
rect 23431 16405 23443 16439
rect 23385 16399 23443 16405
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 9766 16232 9772 16244
rect 7156 16204 9772 16232
rect 7156 16192 7162 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12345 16235 12403 16241
rect 12345 16232 12357 16235
rect 12124 16204 12357 16232
rect 12124 16192 12130 16204
rect 12345 16201 12357 16204
rect 12391 16201 12403 16235
rect 12345 16195 12403 16201
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 13446 16232 13452 16244
rect 12492 16204 13452 16232
rect 12492 16192 12498 16204
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 14182 16232 14188 16244
rect 14143 16204 14188 16232
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 14734 16192 14740 16244
rect 14792 16232 14798 16244
rect 14829 16235 14887 16241
rect 14829 16232 14841 16235
rect 14792 16204 14841 16232
rect 14792 16192 14798 16204
rect 14829 16201 14841 16204
rect 14875 16201 14887 16235
rect 14829 16195 14887 16201
rect 15473 16235 15531 16241
rect 15473 16201 15485 16235
rect 15519 16201 15531 16235
rect 15473 16195 15531 16201
rect 9125 16167 9183 16173
rect 9125 16133 9137 16167
rect 9171 16164 9183 16167
rect 10594 16164 10600 16176
rect 9171 16136 10600 16164
rect 9171 16133 9183 16136
rect 9125 16127 9183 16133
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 13630 16164 13636 16176
rect 12406 16136 13636 16164
rect 1762 16096 1768 16108
rect 1723 16068 1768 16096
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 4893 16099 4951 16105
rect 4893 16096 4905 16099
rect 3752 16068 4905 16096
rect 3752 16056 3758 16068
rect 4893 16065 4905 16068
rect 4939 16065 4951 16099
rect 8386 16096 8392 16108
rect 8347 16068 8392 16096
rect 4893 16059 4951 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 9030 16096 9036 16108
rect 8991 16068 9036 16096
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9364 16068 9873 16096
rect 9364 16056 9370 16068
rect 9861 16065 9873 16068
rect 9907 16096 9919 16099
rect 11238 16096 11244 16108
rect 9907 16068 11244 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 12250 16096 12256 16108
rect 12211 16068 12256 16096
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 9214 16028 9220 16040
rect 2746 16000 9220 16028
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 2746 15960 2774 16000
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 9824 16000 10333 16028
rect 9824 15988 9830 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 1627 15932 2774 15960
rect 8481 15963 8539 15969
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 8481 15929 8493 15963
rect 8527 15960 8539 15963
rect 10226 15960 10232 15972
rect 8527 15932 10232 15960
rect 8527 15929 8539 15932
rect 8481 15923 8539 15929
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 10336 15960 10364 15991
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 12406 16028 12434 16136
rect 13630 16124 13636 16136
rect 13688 16124 13694 16176
rect 15488 16164 15516 16195
rect 17126 16192 17132 16244
rect 17184 16232 17190 16244
rect 21910 16232 21916 16244
rect 17184 16204 21916 16232
rect 17184 16192 17190 16204
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 22204 16204 24440 16232
rect 17494 16164 17500 16176
rect 15488 16136 17356 16164
rect 17455 16136 17500 16164
rect 12710 16056 12716 16108
rect 12768 16096 12774 16108
rect 13081 16099 13139 16105
rect 13081 16096 13093 16099
rect 12768 16068 13093 16096
rect 12768 16056 12774 16068
rect 13081 16065 13093 16068
rect 13127 16096 13139 16099
rect 13170 16096 13176 16108
rect 13127 16068 13176 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 14369 16099 14427 16105
rect 14369 16065 14381 16099
rect 14415 16096 14427 16099
rect 15470 16096 15476 16108
rect 14415 16068 15476 16096
rect 14415 16065 14427 16068
rect 14369 16059 14427 16065
rect 13740 16028 13768 16059
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15654 16096 15660 16108
rect 15615 16068 15660 16096
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 10560 16000 10605 16028
rect 10796 16000 12434 16028
rect 12912 16000 13768 16028
rect 16117 16031 16175 16037
rect 10560 15988 10566 16000
rect 10796 15960 10824 16000
rect 11054 15960 11060 15972
rect 10336 15932 10824 15960
rect 10888 15932 11060 15960
rect 4985 15895 5043 15901
rect 4985 15861 4997 15895
rect 5031 15892 5043 15895
rect 6546 15892 6552 15904
rect 5031 15864 6552 15892
rect 5031 15861 5043 15864
rect 4985 15855 5043 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 9677 15895 9735 15901
rect 9677 15861 9689 15895
rect 9723 15892 9735 15895
rect 10888 15892 10916 15932
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 12912 15969 12940 16000
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 16163 16000 16865 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 16853 15997 16865 16000
rect 16899 15997 16911 16031
rect 17034 16028 17040 16040
rect 16995 16000 17040 16028
rect 16853 15991 16911 15997
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17328 16028 17356 16136
rect 17494 16124 17500 16136
rect 17552 16124 17558 16176
rect 19242 16164 19248 16176
rect 18156 16136 19248 16164
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 18156 16105 18184 16136
rect 19242 16124 19248 16136
rect 19300 16124 19306 16176
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17920 16068 18153 16096
rect 17920 16056 17926 16068
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 18141 16059 18199 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 20990 16096 20996 16108
rect 20102 16068 20996 16096
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21082 16056 21088 16108
rect 21140 16096 21146 16108
rect 22204 16105 22232 16204
rect 22462 16124 22468 16176
rect 22520 16164 22526 16176
rect 24412 16164 24440 16204
rect 24486 16192 24492 16244
rect 24544 16232 24550 16244
rect 24544 16204 24716 16232
rect 24544 16192 24550 16204
rect 24578 16164 24584 16176
rect 22520 16136 22954 16164
rect 24412 16136 24584 16164
rect 22520 16124 22526 16136
rect 24412 16105 24440 16136
rect 24578 16124 24584 16136
rect 24636 16124 24642 16176
rect 24688 16173 24716 16204
rect 24673 16167 24731 16173
rect 24673 16133 24685 16167
rect 24719 16133 24731 16167
rect 24673 16127 24731 16133
rect 25130 16124 25136 16176
rect 25188 16124 25194 16176
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 21140 16068 21281 16096
rect 21140 16056 21146 16068
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 24397 16099 24455 16105
rect 24397 16065 24409 16099
rect 24443 16065 24455 16099
rect 24397 16059 24455 16065
rect 28077 16099 28135 16105
rect 28077 16065 28089 16099
rect 28123 16096 28135 16099
rect 28534 16096 28540 16108
rect 28123 16068 28540 16096
rect 28123 16065 28135 16068
rect 28077 16059 28135 16065
rect 18966 16028 18972 16040
rect 17328 16000 18092 16028
rect 18927 16000 18972 16028
rect 12897 15963 12955 15969
rect 12897 15929 12909 15963
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 15654 15920 15660 15972
rect 15712 15960 15718 15972
rect 15712 15932 17908 15960
rect 15712 15920 15718 15932
rect 9723 15864 10916 15892
rect 9723 15861 9735 15864
rect 9677 15855 9735 15861
rect 10962 15852 10968 15904
rect 11020 15892 11026 15904
rect 13538 15892 13544 15904
rect 11020 15864 11065 15892
rect 13499 15864 13544 15892
rect 11020 15852 11026 15864
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 17880 15892 17908 15932
rect 17957 15895 18015 15901
rect 17957 15892 17969 15895
rect 17880 15864 17969 15892
rect 17957 15861 17969 15864
rect 18003 15861 18015 15895
rect 18064 15892 18092 16000
rect 18966 15988 18972 16000
rect 19024 16028 19030 16040
rect 19518 16028 19524 16040
rect 19024 16000 19524 16028
rect 19024 15988 19030 16000
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 20254 15988 20260 16040
rect 20312 16028 20318 16040
rect 20312 16000 21864 16028
rect 20312 15988 20318 16000
rect 21726 15960 21732 15972
rect 20364 15932 21732 15960
rect 20364 15892 20392 15932
rect 21726 15920 21732 15932
rect 21784 15920 21790 15972
rect 21836 15960 21864 16000
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 22204 16028 22232 16059
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 22462 16028 22468 16040
rect 22152 16000 22232 16028
rect 22277 16000 22468 16028
rect 22152 15988 22158 16000
rect 22277 15960 22305 16000
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 24026 16028 24032 16040
rect 22612 16000 24032 16028
rect 22612 15988 22618 16000
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 26418 16028 26424 16040
rect 26379 16000 26424 16028
rect 26418 15988 26424 16000
rect 26476 15988 26482 16040
rect 21836 15932 22305 15960
rect 18064 15864 20392 15892
rect 17957 15855 18015 15861
rect 20438 15852 20444 15904
rect 20496 15892 20502 15904
rect 21361 15895 21419 15901
rect 20496 15864 20541 15892
rect 20496 15852 20502 15864
rect 21361 15861 21373 15895
rect 21407 15892 21419 15895
rect 21634 15892 21640 15904
rect 21407 15864 21640 15892
rect 21407 15861 21419 15864
rect 21361 15855 21419 15861
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 23934 15892 23940 15904
rect 22244 15864 23940 15892
rect 22244 15852 22250 15864
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 26694 15892 26700 15904
rect 24820 15864 26700 15892
rect 24820 15852 24826 15864
rect 26694 15852 26700 15864
rect 26752 15852 26758 15904
rect 28258 15892 28264 15904
rect 28219 15864 28264 15892
rect 28258 15852 28264 15864
rect 28316 15852 28322 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 6917 15691 6975 15697
rect 6917 15657 6929 15691
rect 6963 15688 6975 15691
rect 9950 15688 9956 15700
rect 6963 15660 9956 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 11057 15691 11115 15697
rect 11057 15657 11069 15691
rect 11103 15688 11115 15691
rect 11146 15688 11152 15700
rect 11103 15660 11152 15688
rect 11103 15657 11115 15660
rect 11057 15651 11115 15657
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 21542 15688 21548 15700
rect 11296 15660 21548 15688
rect 11296 15648 11302 15660
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22094 15688 22100 15700
rect 21744 15660 22100 15688
rect 7742 15580 7748 15632
rect 7800 15580 7806 15632
rect 9861 15623 9919 15629
rect 9861 15589 9873 15623
rect 9907 15620 9919 15623
rect 11164 15620 11192 15648
rect 9907 15592 11100 15620
rect 11164 15592 11652 15620
rect 9907 15589 9919 15592
rect 9861 15583 9919 15589
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 6273 15555 6331 15561
rect 6273 15552 6285 15555
rect 6236 15524 6285 15552
rect 6236 15512 6242 15524
rect 6273 15521 6285 15524
rect 6319 15521 6331 15555
rect 7760 15552 7788 15580
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 7760 15524 7941 15552
rect 6273 15515 6331 15521
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15552 9275 15555
rect 9263 15524 10732 15552
rect 9263 15521 9275 15524
rect 9217 15515 9275 15521
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15484 6515 15487
rect 7742 15484 7748 15496
rect 6503 15456 7748 15484
rect 6503 15453 6515 15456
rect 6457 15447 6515 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9306 15484 9312 15496
rect 9171 15456 9312 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 9876 15456 10425 15484
rect 8021 15419 8079 15425
rect 8021 15385 8033 15419
rect 8067 15416 8079 15419
rect 8386 15416 8392 15428
rect 8067 15388 8392 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 8573 15419 8631 15425
rect 8573 15385 8585 15419
rect 8619 15416 8631 15419
rect 9030 15416 9036 15428
rect 8619 15388 9036 15416
rect 8619 15385 8631 15388
rect 8573 15379 8631 15385
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 9876 15348 9904 15456
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10413 15447 10471 15453
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 10704 15416 10732 15524
rect 11072 15484 11100 15592
rect 11624 15561 11652 15592
rect 16942 15580 16948 15632
rect 17000 15620 17006 15632
rect 17221 15623 17279 15629
rect 17221 15620 17233 15623
rect 17000 15592 17233 15620
rect 17000 15580 17006 15592
rect 17221 15589 17233 15592
rect 17267 15589 17279 15623
rect 21744 15620 21772 15660
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22278 15648 22284 15700
rect 22336 15688 22342 15700
rect 24210 15688 24216 15700
rect 22336 15660 24216 15688
rect 22336 15648 22342 15660
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 26326 15648 26332 15700
rect 26384 15648 26390 15700
rect 17221 15583 17279 15589
rect 21560 15592 21772 15620
rect 11609 15555 11667 15561
rect 11609 15521 11621 15555
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 13538 15512 13544 15564
rect 13596 15552 13602 15564
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 13596 15524 17049 15552
rect 13596 15512 13602 15524
rect 17037 15521 17049 15524
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 18690 15552 18696 15564
rect 18288 15524 18696 15552
rect 18288 15512 18294 15524
rect 18690 15512 18696 15524
rect 18748 15552 18754 15564
rect 19242 15552 19248 15564
rect 18748 15524 19248 15552
rect 18748 15512 18754 15524
rect 19242 15512 19248 15524
rect 19300 15552 19306 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19300 15524 19441 15552
rect 19300 15512 19306 15524
rect 19429 15521 19441 15524
rect 19475 15552 19487 15555
rect 21560 15552 21588 15592
rect 21652 15561 21680 15592
rect 23014 15580 23020 15632
rect 23072 15620 23078 15632
rect 23385 15623 23443 15629
rect 23385 15620 23397 15623
rect 23072 15592 23397 15620
rect 23072 15580 23078 15592
rect 23385 15589 23397 15592
rect 23431 15589 23443 15623
rect 23385 15583 23443 15589
rect 24578 15580 24584 15632
rect 24636 15620 24642 15632
rect 24636 15592 26280 15620
rect 24636 15580 24642 15592
rect 19475 15524 21588 15552
rect 21637 15555 21695 15561
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 21637 15521 21649 15555
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 22922 15512 22928 15564
rect 22980 15552 22986 15564
rect 26252 15561 26280 15592
rect 26237 15555 26295 15561
rect 22980 15524 23244 15552
rect 22980 15512 22986 15524
rect 11146 15484 11152 15496
rect 11072 15456 11152 15484
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 12710 15444 12716 15496
rect 12768 15484 12774 15496
rect 12894 15484 12900 15496
rect 12768 15456 12900 15484
rect 12768 15444 12774 15456
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13078 15484 13084 15496
rect 13039 15456 13084 15484
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15896 15456 15945 15484
rect 15896 15444 15902 15456
rect 15933 15453 15945 15456
rect 15979 15453 15991 15487
rect 16853 15487 16911 15493
rect 16853 15484 16865 15487
rect 15933 15447 15991 15453
rect 16132 15456 16865 15484
rect 11701 15419 11759 15425
rect 11701 15416 11713 15419
rect 10704 15388 11713 15416
rect 11701 15385 11713 15388
rect 11747 15385 11759 15419
rect 11701 15379 11759 15385
rect 12253 15419 12311 15425
rect 12253 15385 12265 15419
rect 12299 15416 12311 15419
rect 13354 15416 13360 15428
rect 12299 15388 13360 15416
rect 12299 15385 12311 15388
rect 12253 15379 12311 15385
rect 8352 15320 9904 15348
rect 8352 15308 8358 15320
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 12406 15348 12434 15388
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 14645 15419 14703 15425
rect 14645 15385 14657 15419
rect 14691 15385 14703 15419
rect 14645 15379 14703 15385
rect 12216 15320 12434 15348
rect 12216 15308 12222 15320
rect 13262 15308 13268 15360
rect 13320 15348 13326 15360
rect 13538 15348 13544 15360
rect 13320 15320 13544 15348
rect 13320 15308 13326 15320
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 14660 15348 14688 15379
rect 14734 15376 14740 15428
rect 14792 15416 14798 15428
rect 15289 15419 15347 15425
rect 14792 15388 14837 15416
rect 14792 15376 14798 15388
rect 15289 15385 15301 15419
rect 15335 15385 15347 15419
rect 15289 15379 15347 15385
rect 15194 15348 15200 15360
rect 14660 15320 15200 15348
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 15304 15348 15332 15379
rect 15378 15376 15384 15428
rect 15436 15416 15442 15428
rect 16132 15416 16160 15456
rect 16853 15453 16865 15456
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 17586 15444 17592 15496
rect 17644 15484 17650 15496
rect 17862 15484 17868 15496
rect 17644 15456 17868 15484
rect 17644 15444 17650 15456
rect 17862 15444 17868 15456
rect 17920 15484 17926 15496
rect 17957 15487 18015 15493
rect 17957 15484 17969 15487
rect 17920 15456 17969 15484
rect 17920 15444 17926 15456
rect 17957 15453 17969 15456
rect 18003 15453 18015 15487
rect 17957 15447 18015 15453
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18196 15456 18613 15484
rect 18196 15444 18202 15456
rect 18601 15453 18613 15456
rect 18647 15484 18659 15487
rect 18782 15484 18788 15496
rect 18647 15456 18788 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 15436 15388 16160 15416
rect 16209 15419 16267 15425
rect 15436 15376 15442 15388
rect 16209 15385 16221 15419
rect 16255 15416 16267 15419
rect 16298 15416 16304 15428
rect 16255 15388 16304 15416
rect 16255 15385 16267 15388
rect 16209 15379 16267 15385
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 16390 15376 16396 15428
rect 16448 15416 16454 15428
rect 19334 15416 19340 15428
rect 16448 15388 19340 15416
rect 16448 15376 16454 15388
rect 19334 15376 19340 15388
rect 19392 15376 19398 15428
rect 19610 15376 19616 15428
rect 19668 15416 19674 15428
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 19668 15388 19717 15416
rect 19668 15376 19674 15388
rect 19705 15385 19717 15388
rect 19751 15385 19763 15419
rect 19705 15379 19763 15385
rect 20714 15376 20720 15428
rect 20772 15376 20778 15428
rect 21818 15416 21824 15428
rect 21100 15388 21824 15416
rect 16574 15348 16580 15360
rect 15304 15320 16580 15348
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 18049 15351 18107 15357
rect 18049 15317 18061 15351
rect 18095 15348 18107 15351
rect 18598 15348 18604 15360
rect 18095 15320 18604 15348
rect 18095 15317 18107 15320
rect 18049 15311 18107 15317
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 18693 15351 18751 15357
rect 18693 15317 18705 15351
rect 18739 15348 18751 15351
rect 21100 15348 21128 15388
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 21910 15376 21916 15428
rect 21968 15416 21974 15428
rect 21968 15388 22013 15416
rect 21968 15376 21974 15388
rect 22370 15376 22376 15428
rect 22428 15376 22434 15428
rect 23216 15416 23244 15524
rect 26237 15521 26249 15555
rect 26283 15521 26295 15555
rect 26344 15552 26372 15648
rect 26513 15555 26571 15561
rect 26513 15552 26525 15555
rect 26344 15524 26525 15552
rect 26237 15515 26295 15521
rect 26513 15521 26525 15524
rect 26559 15521 26571 15555
rect 26513 15515 26571 15521
rect 27706 15512 27712 15564
rect 27764 15512 27770 15564
rect 27724 15484 27752 15512
rect 27646 15456 27752 15484
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 23216 15388 24685 15416
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 24673 15379 24731 15385
rect 24765 15419 24823 15425
rect 24765 15385 24777 15419
rect 24811 15385 24823 15419
rect 24765 15379 24823 15385
rect 25317 15419 25375 15425
rect 25317 15385 25329 15419
rect 25363 15416 25375 15419
rect 25866 15416 25872 15428
rect 25363 15388 25872 15416
rect 25363 15385 25375 15388
rect 25317 15379 25375 15385
rect 18739 15320 21128 15348
rect 21177 15351 21235 15357
rect 18739 15317 18751 15320
rect 18693 15311 18751 15317
rect 21177 15317 21189 15351
rect 21223 15348 21235 15351
rect 21542 15348 21548 15360
rect 21223 15320 21548 15348
rect 21223 15317 21235 15320
rect 21177 15311 21235 15317
rect 21542 15308 21548 15320
rect 21600 15308 21606 15360
rect 21726 15308 21732 15360
rect 21784 15348 21790 15360
rect 24780 15348 24808 15379
rect 25866 15376 25872 15388
rect 25924 15376 25930 15428
rect 27798 15376 27804 15428
rect 27856 15416 27862 15428
rect 28261 15419 28319 15425
rect 28261 15416 28273 15419
rect 27856 15388 28273 15416
rect 27856 15376 27862 15388
rect 28261 15385 28273 15388
rect 28307 15385 28319 15419
rect 28261 15379 28319 15385
rect 21784 15320 24808 15348
rect 21784 15308 21790 15320
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 9033 15147 9091 15153
rect 9033 15144 9045 15147
rect 7800 15116 9045 15144
rect 7800 15104 7806 15116
rect 9033 15113 9045 15116
rect 9079 15113 9091 15147
rect 10870 15144 10876 15156
rect 10831 15116 10876 15144
rect 9033 15107 9091 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 11204 15116 13400 15144
rect 11204 15104 11210 15116
rect 12250 15076 12256 15088
rect 10428 15048 12256 15076
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 15008 8999 15011
rect 9306 15008 9312 15020
rect 8987 14980 9312 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9306 14968 9312 14980
rect 9364 15008 9370 15020
rect 10428 15017 10456 15048
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 9364 14980 9781 15008
rect 9364 14968 9370 14980
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 14977 10471 15011
rect 11054 15008 11060 15020
rect 11015 14980 11060 15008
rect 10413 14971 10471 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 15008 12219 15011
rect 12986 15008 12992 15020
rect 12207 14980 12992 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 13372 15017 13400 15116
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 15749 15147 15807 15153
rect 13504 15116 14320 15144
rect 13504 15104 13510 15116
rect 14292 15076 14320 15116
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 17034 15144 17040 15156
rect 15795 15116 17040 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 19981 15147 20039 15153
rect 18524 15116 19932 15144
rect 14461 15079 14519 15085
rect 14461 15076 14473 15079
rect 14292 15048 14473 15076
rect 14461 15045 14473 15048
rect 14507 15045 14519 15079
rect 14461 15039 14519 15045
rect 16482 15036 16488 15088
rect 16540 15076 16546 15088
rect 18524 15076 18552 15116
rect 16540 15048 18552 15076
rect 16540 15036 16546 15048
rect 18598 15036 18604 15088
rect 18656 15076 18662 15088
rect 19904 15076 19932 15116
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20438 15144 20444 15156
rect 20027 15116 20444 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15113 20591 15147
rect 20533 15107 20591 15113
rect 21361 15147 21419 15153
rect 21361 15113 21373 15147
rect 21407 15144 21419 15147
rect 22370 15144 22376 15156
rect 21407 15116 22376 15144
rect 21407 15113 21419 15116
rect 21361 15107 21419 15113
rect 20346 15076 20352 15088
rect 18656 15048 18998 15076
rect 19904 15048 20352 15076
rect 18656 15036 18662 15048
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 20548 15076 20576 15107
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 22830 15104 22836 15156
rect 22888 15104 22894 15156
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23532 15116 24133 15144
rect 23532 15104 23538 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 25038 15104 25044 15156
rect 25096 15104 25102 15156
rect 22848 15076 22876 15104
rect 20548 15048 22876 15076
rect 23106 15036 23112 15088
rect 23164 15036 23170 15088
rect 24946 15076 24952 15088
rect 23952 15048 24952 15076
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 14977 13231 15011
rect 13173 14971 13231 14977
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 14977 13415 15011
rect 15930 15008 15936 15020
rect 15891 14980 15936 15008
rect 13357 14971 13415 14977
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 9732 14844 10241 14872
rect 9732 14832 9738 14844
rect 10229 14841 10241 14844
rect 10275 14841 10287 14875
rect 12360 14872 12388 14903
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13188 14940 13216 14971
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 18230 15008 18236 15020
rect 16040 14980 17540 15008
rect 18191 14980 18236 15008
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 12492 14912 14381 14940
rect 12492 14900 12498 14912
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14516 14912 14657 14940
rect 14516 14900 14522 14912
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 16040 14940 16068 14980
rect 14884 14912 16068 14940
rect 14884 14900 14890 14912
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 17037 14943 17095 14949
rect 17037 14940 17049 14943
rect 16908 14912 17049 14940
rect 16908 14900 16914 14912
rect 17037 14909 17049 14912
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 13446 14872 13452 14884
rect 12360 14844 13452 14872
rect 10229 14835 10287 14841
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 13648 14844 14504 14872
rect 9585 14807 9643 14813
rect 9585 14773 9597 14807
rect 9631 14804 9643 14807
rect 10134 14804 10140 14816
rect 9631 14776 10140 14804
rect 9631 14773 9643 14776
rect 9585 14767 9643 14773
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 13648 14804 13676 14844
rect 13814 14804 13820 14816
rect 12492 14776 13676 14804
rect 13775 14776 13820 14804
rect 12492 14764 12498 14776
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14476 14804 14504 14844
rect 14550 14832 14556 14884
rect 14608 14872 14614 14884
rect 17236 14872 17264 14903
rect 14608 14844 17264 14872
rect 14608 14832 14614 14844
rect 16482 14804 16488 14816
rect 14476 14776 16488 14804
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 16724 14776 17417 14804
rect 16724 14764 16730 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 17512 14804 17540 14980
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20128 14980 20453 15008
rect 20128 14968 20134 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20622 14968 20628 15020
rect 20680 15008 20686 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 20680 14980 21281 15008
rect 20680 14968 20686 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21358 14968 21364 15020
rect 21416 15008 21422 15020
rect 21416 14980 22094 15008
rect 21416 14968 21422 14980
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18196 14912 18521 14940
rect 18196 14900 18202 14912
rect 18509 14909 18521 14912
rect 18555 14940 18567 14943
rect 19058 14940 19064 14952
rect 18555 14912 19064 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 22066 14940 22094 14980
rect 22186 14968 22192 15020
rect 22244 15008 22250 15020
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 22244 14980 22385 15008
rect 22244 14968 22250 14980
rect 22373 14977 22385 14980
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 22649 14943 22707 14949
rect 22649 14940 22661 14943
rect 22066 14912 22661 14940
rect 22649 14909 22661 14912
rect 22695 14940 22707 14943
rect 23952 14940 23980 15048
rect 24946 15036 24952 15048
rect 25004 15036 25010 15088
rect 25056 15076 25084 15104
rect 25056 15048 25346 15076
rect 27154 15008 27160 15020
rect 27115 14980 27160 15008
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 27982 15008 27988 15020
rect 27943 14980 27988 15008
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 24578 14940 24584 14952
rect 22695 14912 23980 14940
rect 24539 14912 24584 14940
rect 22695 14909 22707 14912
rect 22649 14903 22707 14909
rect 24578 14900 24584 14912
rect 24636 14900 24642 14952
rect 24854 14940 24860 14952
rect 24815 14912 24860 14940
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 26602 14940 26608 14952
rect 26563 14912 26608 14940
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 19610 14832 19616 14884
rect 19668 14872 19674 14884
rect 22278 14872 22284 14884
rect 19668 14844 22284 14872
rect 19668 14832 19674 14844
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 23676 14844 24256 14872
rect 20162 14804 20168 14816
rect 17512 14776 20168 14804
rect 17405 14767 17463 14773
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 23676 14804 23704 14844
rect 20588 14776 23704 14804
rect 24228 14804 24256 14844
rect 24854 14804 24860 14816
rect 24228 14776 24860 14804
rect 20588 14764 20594 14776
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 26234 14764 26240 14816
rect 26292 14804 26298 14816
rect 27249 14807 27307 14813
rect 27249 14804 27261 14807
rect 26292 14776 27261 14804
rect 26292 14764 26298 14776
rect 27249 14773 27261 14776
rect 27295 14773 27307 14807
rect 27249 14767 27307 14773
rect 27614 14764 27620 14816
rect 27672 14804 27678 14816
rect 28077 14807 28135 14813
rect 28077 14804 28089 14807
rect 27672 14776 28089 14804
rect 27672 14764 27678 14776
rect 28077 14773 28089 14776
rect 28123 14773 28135 14807
rect 28077 14767 28135 14773
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 8444 14572 9689 14600
rect 8444 14560 8450 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10502 14600 10508 14612
rect 10008 14572 10508 14600
rect 10008 14560 10014 14572
rect 10502 14560 10508 14572
rect 10560 14600 10566 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 10560 14572 12633 14600
rect 10560 14560 10566 14572
rect 12621 14569 12633 14572
rect 12667 14569 12679 14603
rect 12621 14563 12679 14569
rect 13541 14603 13599 14609
rect 13541 14569 13553 14603
rect 13587 14600 13599 14603
rect 15933 14603 15991 14609
rect 13587 14572 15516 14600
rect 13587 14569 13599 14572
rect 13541 14563 13599 14569
rect 10965 14535 11023 14541
rect 10965 14501 10977 14535
rect 11011 14532 11023 14535
rect 14645 14535 14703 14541
rect 14645 14532 14657 14535
rect 11011 14504 12480 14532
rect 11011 14501 11023 14504
rect 10965 14495 11023 14501
rect 10134 14424 10140 14476
rect 10192 14464 10198 14476
rect 12452 14473 12480 14504
rect 13372 14504 14657 14532
rect 12437 14467 12495 14473
rect 10192 14436 11192 14464
rect 10192 14424 10198 14436
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5810 14396 5816 14408
rect 4939 14368 5816 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 9585 14399 9643 14405
rect 9585 14365 9597 14399
rect 9631 14396 9643 14399
rect 10410 14396 10416 14408
rect 9631 14368 10416 14396
rect 9631 14365 9643 14368
rect 9585 14359 9643 14365
rect 10410 14356 10416 14368
rect 10468 14356 10474 14408
rect 11164 14405 11192 14436
rect 12437 14433 12449 14467
rect 12483 14433 12495 14467
rect 12437 14427 12495 14433
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 11974 14396 11980 14408
rect 11655 14368 11980 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 13372 14396 13400 14504
rect 14645 14501 14657 14504
rect 14691 14501 14703 14535
rect 14645 14495 14703 14501
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 15488 14473 15516 14572
rect 15933 14569 15945 14603
rect 15979 14600 15991 14603
rect 16666 14600 16672 14612
rect 15979 14572 16672 14600
rect 15979 14569 15991 14572
rect 15933 14563 15991 14569
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 21174 14600 21180 14612
rect 16776 14572 21180 14600
rect 15654 14492 15660 14544
rect 15712 14532 15718 14544
rect 16776 14532 16804 14572
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 23566 14560 23572 14612
rect 23624 14600 23630 14612
rect 26786 14600 26792 14612
rect 23624 14572 23669 14600
rect 23768 14572 26792 14600
rect 23624 14560 23630 14572
rect 17586 14532 17592 14544
rect 15712 14504 16804 14532
rect 16868 14504 17592 14532
rect 15712 14492 15718 14504
rect 16868 14476 16896 14504
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 18601 14535 18659 14541
rect 18601 14501 18613 14535
rect 18647 14532 18659 14535
rect 18647 14504 21312 14532
rect 18647 14501 18659 14504
rect 18601 14495 18659 14501
rect 15473 14467 15531 14473
rect 13504 14436 15424 14464
rect 13504 14424 13510 14436
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 12299 14368 12434 14396
rect 13372 14368 13737 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 8754 14328 8760 14340
rect 1596 14300 8760 14328
rect 1596 14269 1624 14300
rect 8754 14288 8760 14300
rect 8812 14288 8818 14340
rect 12406 14328 12434 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 14182 14356 14188 14408
rect 14240 14396 14246 14408
rect 14826 14396 14832 14408
rect 14240 14368 14832 14396
rect 14240 14356 14246 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15396 14396 15424 14436
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 16850 14464 16856 14476
rect 15473 14427 15531 14433
rect 16316 14436 16856 14464
rect 15838 14396 15844 14408
rect 15396 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16316 14328 16344 14436
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17218 14464 17224 14476
rect 17175 14436 17224 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 17310 14424 17316 14476
rect 17368 14464 17374 14476
rect 17862 14464 17868 14476
rect 17368 14436 17868 14464
rect 17368 14424 17374 14436
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 19300 14436 21189 14464
rect 19300 14424 19306 14436
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21284 14464 21312 14504
rect 22646 14492 22652 14544
rect 22704 14532 22710 14544
rect 22925 14535 22983 14541
rect 22925 14532 22937 14535
rect 22704 14504 22937 14532
rect 22704 14492 22710 14504
rect 22925 14501 22937 14504
rect 22971 14532 22983 14535
rect 23768 14532 23796 14572
rect 26786 14560 26792 14572
rect 26844 14560 26850 14612
rect 28169 14603 28227 14609
rect 28169 14569 28181 14603
rect 28215 14600 28227 14603
rect 28442 14600 28448 14612
rect 28215 14572 28448 14600
rect 28215 14569 28227 14572
rect 28169 14563 28227 14569
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 22971 14504 23796 14532
rect 22971 14501 22983 14504
rect 22925 14495 22983 14501
rect 24946 14464 24952 14476
rect 21284 14436 24952 14464
rect 21177 14427 21235 14433
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 26050 14424 26056 14476
rect 26108 14464 26114 14476
rect 26605 14467 26663 14473
rect 26605 14464 26617 14467
rect 26108 14436 26617 14464
rect 26108 14424 26114 14436
rect 26605 14433 26617 14436
rect 26651 14433 26663 14467
rect 26605 14427 26663 14433
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 17460 14368 17601 14396
rect 17460 14356 17466 14368
rect 17589 14365 17601 14368
rect 17635 14396 17647 14399
rect 17678 14396 17684 14408
rect 17635 14368 17684 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18782 14396 18788 14408
rect 18555 14368 18788 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 19334 14396 19340 14408
rect 18840 14368 19340 14396
rect 18840 14356 18846 14368
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 19610 14396 19616 14408
rect 19475 14368 19616 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 19720 14368 20085 14396
rect 16482 14328 16488 14340
rect 12406 14300 16344 14328
rect 16443 14300 16488 14328
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 16577 14331 16635 14337
rect 16577 14297 16589 14331
rect 16623 14328 16635 14331
rect 19521 14331 19579 14337
rect 19521 14328 19533 14331
rect 16623 14300 19533 14328
rect 16623 14297 16635 14300
rect 16577 14291 16635 14297
rect 19521 14297 19533 14300
rect 19567 14297 19579 14331
rect 19521 14291 19579 14297
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14229 1639 14263
rect 1581 14223 1639 14229
rect 4709 14263 4767 14269
rect 4709 14229 4721 14263
rect 4755 14260 4767 14263
rect 4890 14260 4896 14272
rect 4755 14232 4896 14260
rect 4755 14229 4767 14232
rect 4709 14223 4767 14229
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 10226 14260 10232 14272
rect 10187 14232 10232 14260
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 14274 14260 14280 14272
rect 11747 14232 14280 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 17402 14260 17408 14272
rect 15896 14232 17408 14260
rect 15896 14220 15902 14232
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 19720 14260 19748 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 23474 14396 23480 14408
rect 23435 14368 23480 14396
rect 20073 14359 20131 14365
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 24578 14396 24584 14408
rect 24539 14368 24584 14396
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 28350 14396 28356 14408
rect 28311 14368 28356 14396
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 20346 14288 20352 14340
rect 20404 14328 20410 14340
rect 21174 14328 21180 14340
rect 20404 14300 21180 14328
rect 20404 14288 20410 14300
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 21450 14328 21456 14340
rect 21411 14300 21456 14328
rect 21450 14288 21456 14300
rect 21508 14288 21514 14340
rect 24762 14328 24768 14340
rect 22678 14300 24768 14328
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 24857 14331 24915 14337
rect 24857 14297 24869 14331
rect 24903 14328 24915 14331
rect 25130 14328 25136 14340
rect 24903 14300 25136 14328
rect 24903 14297 24915 14300
rect 24857 14291 24915 14297
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 26142 14328 26148 14340
rect 26082 14300 26148 14328
rect 26142 14288 26148 14300
rect 26200 14288 26206 14340
rect 17920 14232 19748 14260
rect 20165 14263 20223 14269
rect 17920 14220 17926 14232
rect 20165 14229 20177 14263
rect 20211 14260 20223 14263
rect 20530 14260 20536 14272
rect 20211 14232 20536 14260
rect 20211 14229 20223 14232
rect 20165 14223 20223 14229
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 20622 14220 20628 14272
rect 20680 14260 20686 14272
rect 22830 14260 22836 14272
rect 20680 14232 22836 14260
rect 20680 14220 20686 14232
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 3234 14056 3240 14068
rect 1627 14028 3240 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 5810 14056 5816 14068
rect 5771 14028 5816 14056
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 10137 14059 10195 14065
rect 10137 14025 10149 14059
rect 10183 14056 10195 14059
rect 10183 14028 11928 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 8849 13991 8907 13997
rect 8849 13957 8861 13991
rect 8895 13988 8907 13991
rect 10594 13988 10600 14000
rect 8895 13960 10600 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 10965 13991 11023 13997
rect 10965 13957 10977 13991
rect 11011 13988 11023 13991
rect 11790 13988 11796 14000
rect 11011 13960 11796 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 11900 13997 11928 14028
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 13136 14028 13553 14056
rect 13136 14016 13142 14028
rect 13541 14025 13553 14028
rect 13587 14025 13599 14059
rect 13541 14019 13599 14025
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14056 14335 14059
rect 14550 14056 14556 14068
rect 14323 14028 14556 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15344 14028 15945 14056
rect 15344 14016 15350 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 15933 14019 15991 14025
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 16632 14028 17632 14056
rect 16632 14016 16638 14028
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13957 11943 13991
rect 11885 13951 11943 13957
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 12124 13960 13492 13988
rect 12124 13948 12130 13960
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 4890 13920 4896 13932
rect 4851 13892 4896 13920
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6362 13920 6368 13932
rect 6043 13892 6368 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 6546 13920 6552 13932
rect 6507 13892 6552 13920
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 8754 13920 8760 13932
rect 8715 13892 8760 13920
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 10226 13920 10232 13932
rect 9631 13892 10232 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 13464 13929 13492 13960
rect 13630 13948 13636 14000
rect 13688 13988 13694 14000
rect 13688 13960 15148 13988
rect 13688 13948 13694 13960
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 13449 13923 13507 13929
rect 12483 13892 13400 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4709 13855 4767 13861
rect 4709 13852 4721 13855
rect 4212 13824 4721 13852
rect 4212 13812 4218 13824
rect 4709 13821 4721 13824
rect 4755 13821 4767 13855
rect 4709 13815 4767 13821
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 6454 13852 6460 13864
rect 5399 13824 6460 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 8478 13852 8484 13864
rect 6779 13824 8484 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 10336 13852 10364 13883
rect 9548 13824 10364 13852
rect 11793 13855 11851 13861
rect 9548 13812 9554 13824
rect 11793 13821 11805 13855
rect 11839 13852 11851 13855
rect 12802 13852 12808 13864
rect 11839 13824 12808 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13372 13852 13400 13892
rect 13449 13889 13461 13923
rect 13495 13889 13507 13923
rect 14182 13920 14188 13932
rect 14143 13892 14188 13920
rect 13449 13883 13507 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14332 13892 15025 13920
rect 14332 13880 14338 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 14550 13852 14556 13864
rect 13372 13824 14556 13852
rect 14550 13812 14556 13824
rect 14608 13812 14614 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15120 13852 15148 13960
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 17604 13997 17632 14028
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18690 14056 18696 14068
rect 18012 14028 18696 14056
rect 18012 14016 18018 14028
rect 18690 14016 18696 14028
rect 18748 14056 18754 14068
rect 19889 14059 19947 14065
rect 18748 14028 19840 14056
rect 18748 14016 18754 14028
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 15252 13960 17049 13988
rect 15252 13948 15258 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13957 17647 13991
rect 18322 13988 18328 14000
rect 17589 13951 17647 13957
rect 18156 13960 18328 13988
rect 18156 13929 18184 13960
rect 18322 13948 18328 13960
rect 18380 13948 18386 14000
rect 19426 13948 19432 14000
rect 19484 13948 19490 14000
rect 19812 13988 19840 14028
rect 19889 14025 19901 14059
rect 19935 14056 19947 14059
rect 20622 14056 20628 14068
rect 19935 14028 20628 14056
rect 19935 14025 19947 14028
rect 19889 14019 19947 14025
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 23753 14059 23811 14065
rect 23753 14056 23765 14059
rect 22066 14028 23765 14056
rect 19812 13960 20392 13988
rect 20364 13929 20392 13960
rect 20898 13948 20904 14000
rect 20956 13988 20962 14000
rect 22066 13988 22094 14028
rect 23753 14025 23765 14028
rect 23799 14025 23811 14059
rect 23753 14019 23811 14025
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 24084 14028 24992 14056
rect 24084 14016 24090 14028
rect 24486 13988 24492 14000
rect 20956 13960 21220 13988
rect 20956 13948 20962 13960
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13920 20407 13923
rect 21082 13920 21088 13932
rect 20395 13892 21088 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 21192 13929 21220 13960
rect 21468 13960 22094 13988
rect 23506 13960 24492 13988
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 21266 13920 21272 13932
rect 21223 13892 21272 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 14875 13824 15148 13852
rect 15473 13855 15531 13861
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15473 13821 15485 13855
rect 15519 13852 15531 13855
rect 16942 13852 16948 13864
rect 15519 13824 16804 13852
rect 16903 13824 16948 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 13170 13744 13176 13796
rect 13228 13784 13234 13796
rect 13630 13784 13636 13796
rect 13228 13756 13636 13784
rect 13228 13744 13234 13756
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 16776 13784 16804 13824
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 18506 13852 18512 13864
rect 18248 13824 18512 13852
rect 17034 13784 17040 13796
rect 16776 13756 17040 13784
rect 17034 13744 17040 13756
rect 17092 13744 17098 13796
rect 17770 13744 17776 13796
rect 17828 13784 17834 13796
rect 18248 13784 18276 13824
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 20441 13855 20499 13861
rect 18840 13824 20392 13852
rect 18840 13812 18846 13824
rect 17828 13756 18276 13784
rect 20364 13784 20392 13824
rect 20441 13821 20453 13855
rect 20487 13852 20499 13855
rect 20714 13852 20720 13864
rect 20487 13824 20720 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 21468 13852 21496 13960
rect 24486 13948 24492 13960
rect 24544 13948 24550 14000
rect 24854 13988 24860 14000
rect 24815 13960 24860 13988
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 24964 13988 24992 14028
rect 25222 14016 25228 14068
rect 25280 14056 25286 14068
rect 25280 14028 26648 14056
rect 25280 14016 25286 14028
rect 26620 13997 26648 14028
rect 26605 13991 26663 13997
rect 24964 13960 25346 13988
rect 26605 13957 26617 13991
rect 26651 13988 26663 13991
rect 26694 13988 26700 14000
rect 26651 13960 26700 13988
rect 26651 13957 26663 13960
rect 26605 13951 26663 13957
rect 26694 13948 26700 13960
rect 26752 13948 26758 14000
rect 22002 13852 22008 13864
rect 20824 13824 21496 13852
rect 21963 13824 22008 13852
rect 20824 13784 20852 13824
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 24578 13852 24584 13864
rect 24539 13824 24584 13852
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 26142 13852 26148 13864
rect 25976 13824 26148 13852
rect 25976 13796 26004 13824
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 20364 13756 20852 13784
rect 17828 13744 17834 13756
rect 25958 13744 25964 13796
rect 26016 13744 26022 13796
rect 7190 13716 7196 13728
rect 7103 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13716 7254 13728
rect 9122 13716 9128 13728
rect 7248 13688 9128 13716
rect 7248 13676 7254 13688
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9398 13716 9404 13728
rect 9359 13688 9404 13716
rect 9398 13676 9404 13688
rect 9456 13676 9462 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 18138 13716 18144 13728
rect 14332 13688 18144 13716
rect 14332 13676 14338 13688
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 18230 13676 18236 13728
rect 18288 13716 18294 13728
rect 18398 13719 18456 13725
rect 18398 13716 18410 13719
rect 18288 13688 18410 13716
rect 18288 13676 18294 13688
rect 18398 13685 18410 13688
rect 18444 13685 18456 13719
rect 18398 13679 18456 13685
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 21082 13716 21088 13728
rect 18564 13688 21088 13716
rect 18564 13676 18570 13688
rect 21082 13676 21088 13688
rect 21140 13676 21146 13728
rect 21174 13676 21180 13728
rect 21232 13716 21238 13728
rect 22262 13719 22320 13725
rect 22262 13716 22274 13719
rect 21232 13688 22274 13716
rect 21232 13676 21238 13688
rect 22262 13685 22274 13688
rect 22308 13685 22320 13719
rect 22262 13679 22320 13685
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 27614 13716 27620 13728
rect 22428 13688 27620 13716
rect 22428 13676 22434 13688
rect 27614 13676 27620 13688
rect 27672 13676 27678 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 3329 13515 3387 13521
rect 3329 13481 3341 13515
rect 3375 13512 3387 13515
rect 4154 13512 4160 13524
rect 3375 13484 4160 13512
rect 3375 13481 3387 13484
rect 3329 13475 3387 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 6454 13472 6460 13524
rect 6512 13512 6518 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 6512 13484 8309 13512
rect 6512 13472 6518 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 13725 13515 13783 13521
rect 8297 13475 8355 13481
rect 8956 13484 12434 13512
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 7009 13447 7067 13453
rect 7009 13444 7021 13447
rect 6696 13416 7021 13444
rect 6696 13404 6702 13416
rect 7009 13413 7021 13416
rect 7055 13413 7067 13447
rect 7009 13407 7067 13413
rect 7190 13376 7196 13388
rect 6656 13348 7196 13376
rect 3234 13308 3240 13320
rect 3195 13280 3240 13308
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13308 4215 13311
rect 4246 13308 4252 13320
rect 4203 13280 4252 13308
rect 4203 13277 4215 13280
rect 4157 13271 4215 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 6656 13317 6684 13348
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 7708 13348 7941 13376
rect 7708 13336 7714 13348
rect 7929 13345 7941 13348
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 5261 13311 5319 13317
rect 4396 13280 4441 13308
rect 4396 13268 4402 13280
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6822 13308 6828 13320
rect 6783 13280 6828 13308
rect 6641 13271 6699 13277
rect 5276 13240 5304 13271
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13308 7803 13311
rect 8294 13308 8300 13320
rect 7791 13280 8300 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 8294 13268 8300 13280
rect 8352 13308 8358 13320
rect 8846 13308 8852 13320
rect 8352 13280 8852 13308
rect 8352 13268 8358 13280
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 5994 13240 6000 13252
rect 5276 13212 6000 13240
rect 5994 13200 6000 13212
rect 6052 13240 6058 13252
rect 8956 13240 8984 13484
rect 9122 13404 9128 13456
rect 9180 13444 9186 13456
rect 11885 13447 11943 13453
rect 11885 13444 11897 13447
rect 9180 13416 11897 13444
rect 9180 13404 9186 13416
rect 11885 13413 11897 13416
rect 11931 13413 11943 13447
rect 12406 13444 12434 13484
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 13814 13512 13820 13524
rect 13771 13484 13820 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 15194 13512 15200 13524
rect 14691 13484 15200 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15841 13515 15899 13521
rect 15841 13481 15853 13515
rect 15887 13512 15899 13515
rect 16942 13512 16948 13524
rect 15887 13484 16948 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 20438 13512 20444 13524
rect 17052 13484 20444 13512
rect 14274 13444 14280 13456
rect 12406 13416 14280 13444
rect 11885 13407 11943 13413
rect 14274 13404 14280 13416
rect 14332 13404 14338 13456
rect 17052 13444 17080 13484
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 24673 13515 24731 13521
rect 24673 13512 24685 13515
rect 21008 13484 24685 13512
rect 14568 13416 17080 13444
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 10367 13348 11713 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 11848 13348 13093 13376
rect 11848 13336 11854 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 10226 13308 10232 13320
rect 10187 13280 10232 13308
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 11054 13308 11060 13320
rect 11015 13280 11060 13308
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 11514 13308 11520 13320
rect 11475 13280 11520 13308
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 14568 13317 14596 13416
rect 17494 13404 17500 13456
rect 17552 13444 17558 13456
rect 18141 13447 18199 13453
rect 18141 13444 18153 13447
rect 17552 13416 18153 13444
rect 17552 13404 17558 13416
rect 18141 13413 18153 13416
rect 18187 13413 18199 13447
rect 18141 13407 18199 13413
rect 20806 13404 20812 13456
rect 20864 13444 20870 13456
rect 21008 13444 21036 13484
rect 24673 13481 24685 13484
rect 24719 13481 24731 13515
rect 24673 13475 24731 13481
rect 24762 13472 24768 13524
rect 24820 13512 24826 13524
rect 25777 13515 25835 13521
rect 25777 13512 25789 13515
rect 24820 13484 25789 13512
rect 24820 13472 24826 13484
rect 25777 13481 25789 13484
rect 25823 13481 25835 13515
rect 25777 13475 25835 13481
rect 26142 13472 26148 13524
rect 26200 13512 26206 13524
rect 27154 13512 27160 13524
rect 26200 13484 27160 13512
rect 26200 13472 26206 13484
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 21174 13444 21180 13456
rect 20864 13416 21036 13444
rect 21135 13416 21180 13444
rect 20864 13404 20870 13416
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 23198 13404 23204 13456
rect 23256 13444 23262 13456
rect 26234 13444 26240 13456
rect 23256 13416 26240 13444
rect 23256 13404 23262 13416
rect 26234 13404 26240 13416
rect 26292 13404 26298 13456
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13376 15255 13379
rect 15746 13376 15752 13388
rect 15243 13348 15752 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 15896 13348 17785 13376
rect 15896 13336 15902 13348
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 19150 13376 19156 13388
rect 17773 13339 17831 13345
rect 17880 13348 19156 13376
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 12406 13280 13277 13308
rect 12406 13240 12434 13280
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 15378 13308 15384 13320
rect 15339 13280 15384 13308
rect 14553 13271 14611 13277
rect 6052 13212 8984 13240
rect 10888 13212 12434 13240
rect 6052 13200 6058 13212
rect 4798 13172 4804 13184
rect 4759 13144 4804 13172
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 5353 13175 5411 13181
rect 5353 13141 5365 13175
rect 5399 13172 5411 13175
rect 6730 13172 6736 13184
rect 5399 13144 6736 13172
rect 5399 13141 5411 13144
rect 5353 13135 5411 13141
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 9582 13172 9588 13184
rect 9543 13144 9588 13172
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10888 13181 10916 13212
rect 12618 13200 12624 13252
rect 12676 13240 12682 13252
rect 14568 13240 14596 13271
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15764 13308 15792 13336
rect 16482 13308 16488 13320
rect 15764 13280 16488 13308
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17880 13308 17908 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 19392 13348 19441 13376
rect 19392 13336 19398 13348
rect 19429 13345 19441 13348
rect 19475 13376 19487 13379
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 19475 13348 21741 13376
rect 19475 13345 19487 13348
rect 19429 13339 19487 13345
rect 21729 13345 21741 13348
rect 21775 13376 21787 13379
rect 22002 13376 22008 13388
rect 21775 13348 22008 13376
rect 21775 13345 21787 13348
rect 21729 13339 21787 13345
rect 22002 13336 22008 13348
rect 22060 13336 22066 13388
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 23477 13379 23535 13385
rect 23477 13376 23489 13379
rect 22152 13348 23489 13376
rect 22152 13336 22158 13348
rect 23477 13345 23489 13348
rect 23523 13345 23535 13379
rect 23477 13339 23535 13345
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 25222 13376 25228 13388
rect 23624 13348 25228 13376
rect 23624 13336 23630 13348
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 25590 13336 25596 13388
rect 25648 13376 25654 13388
rect 26142 13376 26148 13388
rect 25648 13348 26148 13376
rect 25648 13336 25654 13348
rect 17359 13280 17908 13308
rect 17957 13311 18015 13317
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18138 13308 18144 13320
rect 18003 13280 18144 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 23106 13268 23112 13320
rect 23164 13268 23170 13320
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 25685 13311 25743 13317
rect 25685 13277 25697 13311
rect 25731 13308 25743 13311
rect 25792 13308 25820 13348
rect 26142 13336 26148 13348
rect 26200 13336 26206 13388
rect 26326 13376 26332 13388
rect 26287 13348 26332 13376
rect 26326 13336 26332 13348
rect 26384 13336 26390 13388
rect 26605 13379 26663 13385
rect 26605 13345 26617 13379
rect 26651 13376 26663 13379
rect 27614 13376 27620 13388
rect 26651 13348 27620 13376
rect 26651 13345 26663 13348
rect 26605 13339 26663 13345
rect 27614 13336 27620 13348
rect 27672 13336 27678 13388
rect 27890 13336 27896 13388
rect 27948 13376 27954 13388
rect 28353 13379 28411 13385
rect 28353 13376 28365 13379
rect 27948 13348 28365 13376
rect 27948 13336 27954 13348
rect 28353 13345 28365 13348
rect 28399 13345 28411 13379
rect 28353 13339 28411 13345
rect 25731 13280 25820 13308
rect 25731 13277 25743 13280
rect 25685 13271 25743 13277
rect 12676 13212 14596 13240
rect 16669 13243 16727 13249
rect 12676 13200 12682 13212
rect 16669 13209 16681 13243
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 16761 13243 16819 13249
rect 16761 13209 16773 13243
rect 16807 13240 16819 13243
rect 16850 13240 16856 13252
rect 16807 13212 16856 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 12986 13172 12992 13184
rect 12584 13144 12992 13172
rect 12584 13132 12590 13144
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 16684 13172 16712 13203
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 19610 13240 19616 13252
rect 17460 13212 19616 13240
rect 17460 13200 17466 13212
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 19702 13200 19708 13252
rect 19760 13240 19766 13252
rect 19760 13212 19805 13240
rect 20930 13212 21312 13240
rect 19760 13200 19766 13212
rect 17420 13172 17448 13200
rect 16684 13144 17448 13172
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 21174 13172 21180 13184
rect 18932 13144 21180 13172
rect 18932 13132 18938 13144
rect 21174 13132 21180 13144
rect 21232 13132 21238 13184
rect 21284 13172 21312 13212
rect 21542 13200 21548 13252
rect 21600 13240 21606 13252
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21600 13212 22017 13240
rect 21600 13200 21606 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 22186 13172 22192 13184
rect 21284 13144 22192 13172
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 22278 13132 22284 13184
rect 22336 13172 22342 13184
rect 24302 13172 24308 13184
rect 22336 13144 24308 13172
rect 22336 13132 22342 13144
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 24596 13172 24624 13271
rect 24946 13200 24952 13252
rect 25004 13240 25010 13252
rect 25004 13212 27094 13240
rect 25004 13200 25010 13212
rect 27890 13172 27896 13184
rect 24596 13144 27896 13172
rect 27890 13132 27896 13144
rect 27948 13132 27954 13184
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 4246 12968 4252 12980
rect 4207 12940 4252 12968
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4338 12928 4344 12980
rect 4396 12968 4402 12980
rect 5721 12971 5779 12977
rect 5721 12968 5733 12971
rect 4396 12940 5733 12968
rect 4396 12928 4402 12940
rect 5721 12937 5733 12940
rect 5767 12937 5779 12971
rect 5721 12931 5779 12937
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 11977 12971 12035 12977
rect 9272 12940 10640 12968
rect 9272 12928 9278 12940
rect 8849 12903 8907 12909
rect 8849 12869 8861 12903
rect 8895 12900 8907 12903
rect 9398 12900 9404 12912
rect 8895 12872 9404 12900
rect 8895 12869 8907 12872
rect 8849 12863 8907 12869
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 10612 12909 10640 12940
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 15013 12971 15071 12977
rect 12023 12940 13492 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 10505 12903 10563 12909
rect 10505 12900 10517 12903
rect 9640 12872 10517 12900
rect 9640 12860 9646 12872
rect 10505 12869 10517 12872
rect 10551 12869 10563 12903
rect 10505 12863 10563 12869
rect 10597 12903 10655 12909
rect 10597 12869 10609 12903
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 11149 12903 11207 12909
rect 11149 12869 11161 12903
rect 11195 12900 11207 12903
rect 11698 12900 11704 12912
rect 11195 12872 11704 12900
rect 11195 12869 11207 12872
rect 11149 12863 11207 12869
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 11790 12860 11796 12912
rect 11848 12900 11854 12912
rect 12805 12903 12863 12909
rect 12805 12900 12817 12903
rect 11848 12872 12817 12900
rect 11848 12860 11854 12872
rect 12805 12869 12817 12872
rect 12851 12869 12863 12903
rect 12805 12863 12863 12869
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 5902 12832 5908 12844
rect 5863 12804 5908 12832
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6512 12804 6561 12832
rect 6512 12792 6518 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6730 12832 6736 12844
rect 6691 12804 6736 12832
rect 6549 12795 6607 12801
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12526 12832 12532 12844
rect 12207 12804 12532 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 13464 12832 13492 12940
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15378 12968 15384 12980
rect 15059 12940 15384 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 17681 12971 17739 12977
rect 15488 12940 16712 12968
rect 13630 12860 13636 12912
rect 13688 12900 13694 12912
rect 13688 12872 14964 12900
rect 13688 12860 13694 12872
rect 14936 12841 14964 12872
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13464 12804 14013 12832
rect 14001 12801 14013 12804
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12832 14979 12835
rect 15488 12832 15516 12940
rect 15746 12900 15752 12912
rect 15707 12872 15752 12900
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 14967 12804 15516 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8757 12767 8815 12773
rect 8757 12764 8769 12767
rect 8067 12736 8769 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8757 12733 8769 12736
rect 8803 12733 8815 12767
rect 9030 12764 9036 12776
rect 8991 12736 9036 12764
rect 8757 12727 8815 12733
rect 9030 12724 9036 12736
rect 9088 12764 9094 12776
rect 12713 12767 12771 12773
rect 9088 12736 12434 12764
rect 9088 12724 9094 12736
rect 4798 12656 4804 12708
rect 4856 12696 4862 12708
rect 6917 12699 6975 12705
rect 6917 12696 6929 12699
rect 4856 12668 6929 12696
rect 4856 12656 4862 12668
rect 6917 12665 6929 12668
rect 6963 12665 6975 12699
rect 12406 12696 12434 12736
rect 12713 12733 12725 12767
rect 12759 12764 12771 12767
rect 12802 12764 12808 12776
rect 12759 12736 12808 12764
rect 12759 12733 12771 12736
rect 12713 12727 12771 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 12986 12764 12992 12776
rect 12947 12736 12992 12764
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 13136 12736 15669 12764
rect 13136 12724 13142 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16574 12764 16580 12776
rect 16347 12736 16580 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 16684 12764 16712 12940
rect 17681 12937 17693 12971
rect 17727 12968 17739 12971
rect 18138 12968 18144 12980
rect 17727 12940 18144 12968
rect 17727 12937 17739 12940
rect 17681 12931 17739 12937
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 21634 12928 21640 12980
rect 21692 12968 21698 12980
rect 24118 12968 24124 12980
rect 21692 12940 24124 12968
rect 21692 12928 21698 12940
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 24302 12968 24308 12980
rect 24263 12940 24308 12968
rect 24302 12928 24308 12940
rect 24360 12928 24366 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 26326 12968 26332 12980
rect 24820 12940 26332 12968
rect 24820 12928 24826 12940
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 26513 12971 26571 12977
rect 26513 12937 26525 12971
rect 26559 12968 26571 12971
rect 26602 12968 26608 12980
rect 26559 12940 26608 12968
rect 26559 12937 26571 12940
rect 26513 12931 26571 12937
rect 26602 12928 26608 12940
rect 26660 12928 26666 12980
rect 18690 12900 18696 12912
rect 16868 12872 18696 12900
rect 16868 12841 16896 12872
rect 18690 12860 18696 12872
rect 18748 12860 18754 12912
rect 19702 12900 19708 12912
rect 19663 12872 19708 12900
rect 19702 12860 19708 12872
rect 19760 12860 19766 12912
rect 22278 12900 22284 12912
rect 20930 12872 22284 12900
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 22830 12900 22836 12912
rect 22791 12872 22836 12900
rect 22830 12860 22836 12872
rect 22888 12860 22894 12912
rect 24210 12860 24216 12912
rect 24268 12900 24274 12912
rect 24268 12872 25530 12900
rect 24268 12860 24274 12872
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 17770 12832 17776 12844
rect 17635 12804 17776 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18138 12792 18144 12844
rect 18196 12832 18202 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 18196 12804 18429 12832
rect 18196 12792 18202 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 19392 12804 19441 12832
rect 19392 12792 19398 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 24302 12832 24308 12844
rect 23966 12804 24308 12832
rect 19429 12795 19487 12801
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 24578 12792 24584 12844
rect 24636 12832 24642 12844
rect 24762 12832 24768 12844
rect 24636 12804 24768 12832
rect 24636 12792 24642 12804
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 28350 12832 28356 12844
rect 28311 12804 28356 12832
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 18233 12767 18291 12773
rect 16684 12736 17080 12764
rect 13817 12699 13875 12705
rect 12406 12668 13216 12696
rect 6917 12659 6975 12665
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 4062 12628 4068 12640
rect 1627 12600 4068 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11514 12628 11520 12640
rect 11204 12600 11520 12628
rect 11204 12588 11210 12600
rect 11514 12588 11520 12600
rect 11572 12628 11578 12640
rect 13078 12628 13084 12640
rect 11572 12600 13084 12628
rect 11572 12588 11578 12600
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13188 12628 13216 12668
rect 13817 12665 13829 12699
rect 13863 12696 13875 12699
rect 14734 12696 14740 12708
rect 13863 12668 14740 12696
rect 13863 12665 13875 12668
rect 13817 12659 13875 12665
rect 14734 12656 14740 12668
rect 14792 12656 14798 12708
rect 15286 12628 15292 12640
rect 13188 12600 15292 12628
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 16942 12628 16948 12640
rect 16903 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 17052 12628 17080 12736
rect 18233 12733 18245 12767
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12764 18935 12767
rect 19794 12764 19800 12776
rect 18923 12736 19800 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 18248 12696 18276 12727
rect 19794 12724 19800 12736
rect 19852 12724 19858 12776
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 20824 12736 21465 12764
rect 20824 12708 20852 12736
rect 21453 12733 21465 12736
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 22186 12724 22192 12776
rect 22244 12764 22250 12776
rect 22557 12767 22615 12773
rect 22557 12764 22569 12767
rect 22244 12736 22569 12764
rect 22244 12724 22250 12736
rect 22557 12733 22569 12736
rect 22603 12733 22615 12767
rect 22557 12727 22615 12733
rect 18248 12668 19564 12696
rect 19242 12628 19248 12640
rect 17052 12600 19248 12628
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19536 12628 19564 12668
rect 20806 12656 20812 12708
rect 20864 12656 20870 12708
rect 20916 12668 21956 12696
rect 20916 12628 20944 12668
rect 19536 12600 20944 12628
rect 21928 12628 21956 12668
rect 23198 12628 23204 12640
rect 21928 12600 23204 12628
rect 23198 12588 23204 12600
rect 23256 12588 23262 12640
rect 25028 12631 25086 12637
rect 25028 12597 25040 12631
rect 25074 12628 25086 12631
rect 25222 12628 25228 12640
rect 25074 12600 25228 12628
rect 25074 12597 25086 12600
rect 25028 12591 25086 12597
rect 25222 12588 25228 12600
rect 25280 12628 25286 12640
rect 25590 12628 25596 12640
rect 25280 12600 25596 12628
rect 25280 12588 25286 12600
rect 25590 12588 25596 12600
rect 25648 12628 25654 12640
rect 26418 12628 26424 12640
rect 25648 12600 26424 12628
rect 25648 12588 25654 12600
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 28166 12628 28172 12640
rect 28127 12600 28172 12628
rect 28166 12588 28172 12600
rect 28224 12588 28230 12640
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 6822 12424 6828 12436
rect 6779 12396 6828 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7650 12424 7656 12436
rect 7611 12396 7656 12424
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 11054 12424 11060 12436
rect 9907 12396 11060 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11790 12424 11796 12436
rect 11751 12396 11796 12424
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 15841 12427 15899 12433
rect 11940 12396 14228 12424
rect 11940 12384 11946 12396
rect 7742 12316 7748 12368
rect 7800 12356 7806 12368
rect 9306 12356 9312 12368
rect 7800 12328 9312 12356
rect 7800 12316 7806 12328
rect 9306 12316 9312 12328
rect 9364 12316 9370 12368
rect 11241 12359 11299 12365
rect 11241 12325 11253 12359
rect 11287 12356 11299 12359
rect 14090 12356 14096 12368
rect 11287 12328 14096 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 14200 12356 14228 12396
rect 15841 12393 15853 12427
rect 15887 12424 15899 12427
rect 15930 12424 15936 12436
rect 15887 12396 15936 12424
rect 15887 12393 15899 12396
rect 15841 12387 15899 12393
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 18138 12424 18144 12436
rect 18099 12396 18144 12424
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 19306 12396 21036 12424
rect 19306 12356 19334 12396
rect 14200 12328 19334 12356
rect 21008 12356 21036 12396
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 22612 12396 25329 12424
rect 22612 12384 22618 12396
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 21542 12356 21548 12368
rect 21008 12328 21548 12356
rect 21542 12316 21548 12328
rect 21600 12316 21606 12368
rect 23658 12316 23664 12368
rect 23716 12356 23722 12368
rect 24029 12359 24087 12365
rect 24029 12356 24041 12359
rect 23716 12328 24041 12356
rect 23716 12316 23722 12328
rect 24029 12325 24041 12328
rect 24075 12325 24087 12359
rect 24029 12319 24087 12325
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 11882 12288 11888 12300
rect 6420 12260 11888 12288
rect 6420 12248 6426 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 4939 12192 5549 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5718 12220 5724 12232
rect 5679 12192 5724 12220
rect 5537 12183 5595 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7190 12220 7196 12232
rect 6687 12192 7196 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7484 12220 7512 12260
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 13078 12288 13084 12300
rect 13039 12260 13084 12288
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13538 12248 13544 12300
rect 13596 12288 13602 12300
rect 14292 12288 14504 12300
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 13596 12272 14565 12288
rect 13596 12260 14320 12272
rect 14476 12260 14565 12272
rect 13596 12248 13602 12260
rect 14553 12257 14565 12260
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16632 12260 16865 12288
rect 16632 12248 16638 12260
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 16942 12248 16948 12300
rect 17000 12288 17006 12300
rect 17402 12288 17408 12300
rect 17000 12260 17408 12288
rect 17000 12248 17006 12260
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19392 12260 19717 12288
rect 19392 12248 19398 12260
rect 19705 12257 19717 12260
rect 19751 12288 19763 12291
rect 20622 12288 20628 12300
rect 19751 12260 20628 12288
rect 19751 12257 19763 12260
rect 19705 12251 19763 12257
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 20990 12248 20996 12300
rect 21048 12288 21054 12300
rect 24673 12291 24731 12297
rect 24673 12288 24685 12291
rect 21048 12260 24685 12288
rect 21048 12248 21054 12260
rect 24673 12257 24685 12260
rect 24719 12257 24731 12291
rect 24673 12251 24731 12257
rect 25038 12248 25044 12300
rect 25096 12288 25102 12300
rect 27985 12291 28043 12297
rect 27985 12288 27997 12291
rect 25096 12260 27997 12288
rect 25096 12248 25102 12260
rect 27985 12257 27997 12260
rect 28031 12257 28043 12291
rect 27985 12251 28043 12257
rect 7553 12223 7611 12229
rect 7553 12220 7565 12223
rect 7484 12192 7565 12220
rect 7553 12189 7565 12192
rect 7599 12189 7611 12223
rect 7553 12183 7611 12189
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9674 12220 9680 12232
rect 9447 12192 9680 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 8588 12152 8616 12183
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9824 12192 10057 12220
rect 9824 12180 9830 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12220 11207 12223
rect 11790 12220 11796 12232
rect 11195 12192 11796 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 10226 12152 10232 12164
rect 8588 12124 10232 12152
rect 10226 12112 10232 12124
rect 10284 12112 10290 12164
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 6638 12084 6644 12096
rect 6227 12056 6644 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 8389 12087 8447 12093
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 9582 12084 9588 12096
rect 8435 12056 9588 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10505 12087 10563 12093
rect 10505 12053 10517 12087
rect 10551 12084 10563 12087
rect 11698 12084 11704 12096
rect 10551 12056 11704 12084
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 11992 12084 12020 12183
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12492 12192 12537 12220
rect 12492 12180 12498 12192
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12952 12192 13277 12220
rect 12952 12180 12958 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 12529 12155 12587 12161
rect 12529 12121 12541 12155
rect 12575 12152 12587 12155
rect 14645 12155 14703 12161
rect 12575 12124 14504 12152
rect 12575 12121 12587 12124
rect 12529 12115 12587 12121
rect 12802 12084 12808 12096
rect 11992 12056 12808 12084
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13725 12087 13783 12093
rect 13725 12084 13737 12087
rect 13504 12056 13737 12084
rect 13504 12044 13510 12056
rect 13725 12053 13737 12056
rect 13771 12053 13783 12087
rect 14476 12084 14504 12124
rect 14645 12121 14657 12155
rect 14691 12121 14703 12155
rect 14645 12115 14703 12121
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 15930 12152 15936 12164
rect 15243 12124 15936 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 14660 12084 14688 12115
rect 15930 12112 15936 12124
rect 15988 12112 15994 12164
rect 14476 12056 14688 12084
rect 16040 12084 16068 12183
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 18046 12220 18052 12232
rect 17276 12192 17816 12220
rect 18007 12192 18052 12220
rect 17276 12180 17282 12192
rect 17788 12164 17816 12192
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18690 12220 18696 12232
rect 18651 12192 18696 12220
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 22278 12220 22284 12232
rect 22239 12192 22284 12220
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 23658 12180 23664 12232
rect 23716 12180 23722 12232
rect 24394 12180 24400 12232
rect 24452 12220 24458 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24452 12192 24593 12220
rect 24452 12180 24458 12192
rect 24581 12189 24593 12192
rect 24627 12220 24639 12223
rect 24762 12220 24768 12232
rect 24627 12192 24768 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 24762 12180 24768 12192
rect 24820 12220 24826 12232
rect 25225 12223 25283 12229
rect 25225 12220 25237 12223
rect 24820 12192 25237 12220
rect 24820 12180 24826 12192
rect 25225 12189 25237 12192
rect 25271 12189 25283 12223
rect 26234 12220 26240 12232
rect 26195 12192 26240 12220
rect 25225 12183 25283 12189
rect 26234 12180 26240 12192
rect 26292 12180 26298 12232
rect 16574 12152 16580 12164
rect 16535 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 16669 12155 16727 12161
rect 16669 12121 16681 12155
rect 16715 12152 16727 12155
rect 17494 12152 17500 12164
rect 16715 12124 17500 12152
rect 16715 12121 16727 12124
rect 16669 12115 16727 12121
rect 17494 12112 17500 12124
rect 17552 12112 17558 12164
rect 17770 12112 17776 12164
rect 17828 12152 17834 12164
rect 19886 12152 19892 12164
rect 17828 12124 19892 12152
rect 17828 12112 17834 12124
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 19978 12112 19984 12164
rect 20036 12152 20042 12164
rect 20036 12124 20081 12152
rect 20036 12112 20042 12124
rect 20990 12112 20996 12164
rect 21048 12112 21054 12164
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 21600 12124 21741 12152
rect 21600 12112 21606 12124
rect 21729 12121 21741 12124
rect 21775 12121 21787 12155
rect 22557 12155 22615 12161
rect 21729 12115 21787 12121
rect 22066 12124 22508 12152
rect 17218 12084 17224 12096
rect 16040 12056 17224 12084
rect 13725 12047 13783 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 18690 12084 18696 12096
rect 17460 12056 18696 12084
rect 17460 12044 17466 12056
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 22066 12084 22094 12124
rect 18831 12056 22094 12084
rect 22480 12084 22508 12124
rect 22557 12121 22569 12155
rect 22603 12152 22615 12155
rect 22646 12152 22652 12164
rect 22603 12124 22652 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 22646 12112 22652 12124
rect 22704 12112 22710 12164
rect 25866 12152 25872 12164
rect 23860 12124 25872 12152
rect 23474 12084 23480 12096
rect 22480 12056 23480 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23860 12084 23888 12124
rect 25866 12112 25872 12124
rect 25924 12112 25930 12164
rect 26510 12152 26516 12164
rect 26471 12124 26516 12152
rect 26510 12112 26516 12124
rect 26568 12112 26574 12164
rect 26620 12124 27002 12152
rect 23624 12056 23888 12084
rect 23624 12044 23630 12056
rect 24302 12044 24308 12096
rect 24360 12084 24366 12096
rect 26620 12084 26648 12124
rect 24360 12056 26648 12084
rect 24360 12044 24366 12056
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 5902 11880 5908 11892
rect 5767 11852 5908 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 9401 11883 9459 11889
rect 9401 11880 9413 11883
rect 8536 11852 9413 11880
rect 8536 11840 8542 11852
rect 9401 11849 9413 11852
rect 9447 11849 9459 11883
rect 9401 11843 9459 11849
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 13262 11880 13268 11892
rect 10284 11852 13268 11880
rect 10284 11840 10290 11852
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11880 13510 11892
rect 15381 11883 15439 11889
rect 13504 11852 14044 11880
rect 13504 11840 13510 11852
rect 7576 11784 8616 11812
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 5994 11744 6000 11756
rect 5951 11716 6000 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 7190 11744 7196 11756
rect 7103 11716 7196 11744
rect 7190 11704 7196 11716
rect 7248 11744 7254 11756
rect 7576 11744 7604 11784
rect 7248 11716 7604 11744
rect 7653 11747 7711 11753
rect 7248 11704 7254 11716
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 7668 11676 7696 11707
rect 8294 11676 8300 11688
rect 1636 11648 7696 11676
rect 8255 11648 8300 11676
rect 1636 11636 1642 11648
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8478 11676 8484 11688
rect 8439 11648 8484 11676
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 8588 11676 8616 11784
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 10134 11812 10140 11824
rect 8812 11784 10140 11812
rect 8812 11772 8818 11784
rect 10134 11772 10140 11784
rect 10192 11772 10198 11824
rect 10502 11812 10508 11824
rect 10463 11784 10508 11812
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 10597 11815 10655 11821
rect 10597 11781 10609 11815
rect 10643 11812 10655 11815
rect 10686 11812 10692 11824
rect 10643 11784 10692 11812
rect 10643 11781 10655 11784
rect 10597 11775 10655 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 10870 11772 10876 11824
rect 10928 11812 10934 11824
rect 14016 11821 14044 11852
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15746 11880 15752 11892
rect 15427 11852 15752 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16117 11883 16175 11889
rect 16117 11849 16129 11883
rect 16163 11880 16175 11883
rect 16758 11880 16764 11892
rect 16163 11852 16764 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 19702 11880 19708 11892
rect 16868 11852 19708 11880
rect 14001 11815 14059 11821
rect 10928 11784 13860 11812
rect 10928 11772 10934 11784
rect 9582 11744 9588 11756
rect 9543 11716 9588 11744
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 11698 11744 11704 11756
rect 11659 11716 11704 11744
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11882 11676 11888 11688
rect 8588 11648 11192 11676
rect 11843 11648 11888 11676
rect 7466 11568 7472 11620
rect 7524 11608 7530 11620
rect 9674 11608 9680 11620
rect 7524 11580 9680 11608
rect 7524 11568 7530 11580
rect 9674 11568 9680 11580
rect 9732 11608 9738 11620
rect 11057 11611 11115 11617
rect 11057 11608 11069 11611
rect 9732 11580 11069 11608
rect 9732 11568 9738 11580
rect 11057 11577 11069 11580
rect 11103 11577 11115 11611
rect 11164 11608 11192 11648
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12584 11648 12817 11676
rect 12584 11636 12590 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12986 11676 12992 11688
rect 12947 11648 12992 11676
rect 12805 11639 12863 11645
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 13722 11608 13728 11620
rect 11164 11580 13728 11608
rect 11057 11571 11115 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 13832 11608 13860 11784
rect 14001 11781 14013 11815
rect 14047 11781 14059 11815
rect 14001 11775 14059 11781
rect 14090 11772 14096 11824
rect 14148 11812 14154 11824
rect 16868 11812 16896 11852
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 23014 11880 23020 11892
rect 20036 11852 23020 11880
rect 20036 11840 20042 11852
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 23753 11883 23811 11889
rect 23753 11849 23765 11883
rect 23799 11880 23811 11883
rect 23934 11880 23940 11892
rect 23799 11852 23940 11880
rect 23799 11849 23811 11852
rect 23753 11843 23811 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 14148 11784 14193 11812
rect 14752 11784 16896 11812
rect 16945 11815 17003 11821
rect 14148 11772 14154 11784
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 14056 11648 14289 11676
rect 14056 11636 14062 11648
rect 14277 11645 14289 11648
rect 14323 11676 14335 11679
rect 14642 11676 14648 11688
rect 14323 11648 14648 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 14752 11608 14780 11784
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 18966 11812 18972 11824
rect 16991 11784 18972 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 18966 11772 18972 11784
rect 19024 11772 19030 11824
rect 22186 11812 22192 11824
rect 19918 11784 22192 11812
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 22281 11815 22339 11821
rect 22281 11781 22293 11815
rect 22327 11812 22339 11815
rect 22370 11812 22376 11824
rect 22327 11784 22376 11812
rect 22327 11781 22339 11784
rect 22281 11775 22339 11781
rect 22370 11772 22376 11784
rect 22428 11772 22434 11824
rect 23290 11772 23296 11824
rect 23348 11772 23354 11824
rect 23842 11772 23848 11824
rect 23900 11812 23906 11824
rect 23900 11784 25346 11812
rect 23900 11772 23906 11784
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 17310 11744 17316 11756
rect 16899 11716 17316 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 13832 11580 14780 11608
rect 15304 11608 15332 11707
rect 16316 11676 16344 11707
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 18046 11744 18052 11756
rect 17727 11716 18052 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 22002 11744 22008 11756
rect 21963 11716 22008 11744
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 24578 11744 24584 11756
rect 24539 11716 24584 11744
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 18138 11676 18144 11688
rect 16316 11648 18144 11676
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 18288 11648 18429 11676
rect 18288 11636 18294 11648
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 18690 11676 18696 11688
rect 18651 11648 18696 11676
rect 18417 11639 18475 11645
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 18840 11648 20177 11676
rect 18840 11636 18846 11648
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 21082 11636 21088 11688
rect 21140 11676 21146 11688
rect 23934 11676 23940 11688
rect 21140 11648 23940 11676
rect 21140 11636 21146 11648
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 24026 11636 24032 11688
rect 24084 11676 24090 11688
rect 24854 11676 24860 11688
rect 24084 11648 24860 11676
rect 24084 11636 24090 11648
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 24946 11636 24952 11688
rect 25004 11676 25010 11688
rect 26605 11679 26663 11685
rect 26605 11676 26617 11679
rect 25004 11648 26617 11676
rect 25004 11636 25010 11648
rect 26605 11645 26617 11648
rect 26651 11645 26663 11679
rect 26605 11639 26663 11645
rect 16942 11608 16948 11620
rect 15304 11580 16948 11608
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17218 11568 17224 11620
rect 17276 11608 17282 11620
rect 17276 11580 17908 11608
rect 17276 11568 17282 11580
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7190 11540 7196 11552
rect 7055 11512 7196 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 7745 11543 7803 11549
rect 7745 11509 7757 11543
rect 7791 11540 7803 11543
rect 8754 11540 8760 11552
rect 7791 11512 8760 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 8941 11543 8999 11549
rect 8941 11509 8953 11543
rect 8987 11540 8999 11543
rect 9398 11540 9404 11552
rect 8987 11512 9404 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 12066 11540 12072 11552
rect 9640 11512 12072 11540
rect 9640 11500 9646 11512
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12345 11543 12403 11549
rect 12345 11509 12357 11543
rect 12391 11540 12403 11543
rect 12710 11540 12716 11552
rect 12391 11512 12716 11540
rect 12391 11509 12403 11512
rect 12345 11503 12403 11509
rect 12710 11500 12716 11512
rect 12768 11540 12774 11552
rect 13078 11540 13084 11552
rect 12768 11512 13084 11540
rect 12768 11500 12774 11512
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 17402 11540 17408 11552
rect 13320 11512 17408 11540
rect 13320 11500 13326 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 17497 11543 17555 11549
rect 17497 11509 17509 11543
rect 17543 11540 17555 11543
rect 17770 11540 17776 11552
rect 17543 11512 17776 11540
rect 17543 11509 17555 11512
rect 17497 11503 17555 11509
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 17880 11540 17908 11580
rect 19720 11580 22094 11608
rect 19720 11540 19748 11580
rect 17880 11512 19748 11540
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21542 11540 21548 11552
rect 20864 11512 21548 11540
rect 20864 11500 20870 11512
rect 21542 11500 21548 11512
rect 21600 11500 21606 11552
rect 22066 11540 22094 11580
rect 26510 11540 26516 11552
rect 22066 11512 26516 11540
rect 26510 11500 26516 11512
rect 26568 11500 26574 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 7009 11339 7067 11345
rect 7009 11336 7021 11339
rect 5776 11308 7021 11336
rect 5776 11296 5782 11308
rect 7009 11305 7021 11308
rect 7055 11305 7067 11339
rect 7009 11299 7067 11305
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8478 11336 8484 11348
rect 7699 11308 8484 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9582 11336 9588 11348
rect 9364 11308 9588 11336
rect 9364 11296 9370 11308
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 12250 11336 12256 11348
rect 10643 11308 12256 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12529 11339 12587 11345
rect 12360 11308 12480 11336
rect 10686 11268 10692 11280
rect 8496 11240 10692 11268
rect 8496 11209 8524 11240
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 12360 11268 12388 11308
rect 10836 11240 12388 11268
rect 12452 11268 12480 11308
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12986 11336 12992 11348
rect 12575 11308 12992 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 14366 11296 14372 11348
rect 14424 11336 14430 11348
rect 14550 11336 14556 11348
rect 14424 11308 14556 11336
rect 14424 11296 14430 11308
rect 14550 11296 14556 11308
rect 14608 11336 14614 11348
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 14608 11308 14657 11336
rect 14608 11296 14614 11308
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 14645 11299 14703 11305
rect 15381 11339 15439 11345
rect 15381 11305 15393 11339
rect 15427 11336 15439 11339
rect 15470 11336 15476 11348
rect 15427 11308 15476 11336
rect 15427 11305 15439 11308
rect 15381 11299 15439 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16298 11336 16304 11348
rect 15620 11308 16304 11336
rect 15620 11296 15626 11308
rect 16298 11296 16304 11308
rect 16356 11336 16362 11348
rect 16356 11308 18000 11336
rect 16356 11296 16362 11308
rect 12618 11268 12624 11280
rect 12452 11240 12624 11268
rect 10836 11228 10842 11240
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 17218 11268 17224 11280
rect 13556 11240 17224 11268
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9398 11200 9404 11212
rect 9263 11172 9404 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 11330 11200 11336 11212
rect 11291 11172 11336 11200
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 13556 11200 13584 11240
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 17589 11271 17647 11277
rect 17589 11237 17601 11271
rect 17635 11237 17647 11271
rect 17589 11231 17647 11237
rect 12124 11172 13584 11200
rect 12124 11160 12130 11172
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 13688 11172 14473 11200
rect 13688 11160 13694 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17402 11200 17408 11212
rect 17175 11172 17408 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7340 11104 7849 11132
rect 7340 11092 7346 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 10778 11132 10784 11144
rect 10739 11104 10784 11132
rect 8389 11095 8447 11101
rect 8404 11064 8432 11095
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12618 11132 12624 11144
rect 12483 11104 12624 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 12618 11092 12624 11104
rect 12676 11132 12682 11144
rect 12986 11132 12992 11144
rect 12676 11104 12992 11132
rect 12676 11092 12682 11104
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13538 11132 13544 11144
rect 13499 11104 13544 11132
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 8404 11036 9260 11064
rect 9232 10996 9260 11036
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 9364 11036 9409 11064
rect 9364 11024 9370 11036
rect 10410 11024 10416 11076
rect 10468 11064 10474 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 10468 11036 11437 11064
rect 10468 11024 10474 11036
rect 11425 11033 11437 11036
rect 11471 11033 11483 11067
rect 11425 11027 11483 11033
rect 11977 11067 12035 11073
rect 11977 11033 11989 11067
rect 12023 11064 12035 11067
rect 12342 11064 12348 11076
rect 12023 11036 12348 11064
rect 12023 11033 12035 11036
rect 11977 11027 12035 11033
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 14292 11064 14320 11095
rect 14734 11092 14740 11144
rect 14792 11132 14798 11144
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 14792 11104 15577 11132
rect 14792 11092 14798 11104
rect 15565 11101 15577 11104
rect 15611 11132 15623 11135
rect 15746 11132 15752 11144
rect 15611 11104 15752 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 17604 11132 17632 11231
rect 16960 11104 17632 11132
rect 15838 11064 15844 11076
rect 14292 11036 15844 11064
rect 15838 11024 15844 11036
rect 15896 11064 15902 11076
rect 16114 11064 16120 11076
rect 15896 11036 16120 11064
rect 15896 11024 15902 11036
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 16209 11067 16267 11073
rect 16209 11033 16221 11067
rect 16255 11064 16267 11067
rect 16960 11064 16988 11104
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 17972 11132 18000 11308
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 22646 11336 22652 11348
rect 18104 11308 22652 11336
rect 18104 11296 18110 11308
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 23658 11336 23664 11348
rect 23619 11308 23664 11336
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24486 11296 24492 11348
rect 24544 11336 24550 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 24544 11308 25053 11336
rect 24544 11296 24550 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 26418 11296 26424 11348
rect 26476 11336 26482 11348
rect 26476 11308 27660 11336
rect 26476 11296 26482 11308
rect 18138 11228 18144 11280
rect 18196 11268 18202 11280
rect 20073 11271 20131 11277
rect 20073 11268 20085 11271
rect 18196 11240 20085 11268
rect 18196 11228 18202 11240
rect 20073 11237 20085 11240
rect 20119 11237 20131 11271
rect 24394 11268 24400 11280
rect 20073 11231 20131 11237
rect 23124 11240 24400 11268
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 19610 11200 19616 11212
rect 18371 11172 19616 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 20622 11160 20628 11212
rect 20680 11200 20686 11212
rect 21361 11203 21419 11209
rect 21361 11200 21373 11203
rect 20680 11172 21373 11200
rect 20680 11160 20686 11172
rect 21361 11169 21373 11172
rect 21407 11200 21419 11203
rect 22278 11200 22284 11212
rect 21407 11172 22284 11200
rect 21407 11169 21419 11172
rect 21361 11163 21419 11169
rect 22278 11160 22284 11172
rect 22336 11160 22342 11212
rect 23014 11160 23020 11212
rect 23072 11200 23078 11212
rect 23124 11209 23152 11240
rect 24394 11228 24400 11240
rect 24452 11228 24458 11280
rect 23109 11203 23167 11209
rect 23109 11200 23121 11203
rect 23072 11172 23121 11200
rect 23072 11160 23078 11172
rect 23109 11169 23121 11172
rect 23155 11169 23167 11203
rect 26142 11200 26148 11212
rect 23109 11163 23167 11169
rect 23584 11172 26148 11200
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17828 11104 17873 11132
rect 17972 11104 18245 11132
rect 17828 11092 17834 11104
rect 18233 11101 18245 11104
rect 18279 11132 18291 11135
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 18279 11104 19441 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11132 19579 11135
rect 19794 11132 19800 11144
rect 19567 11104 19800 11132
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 19886 11092 19892 11144
rect 19944 11132 19950 11144
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19944 11104 20269 11132
rect 19944 11092 19950 11104
rect 20257 11101 20269 11104
rect 20303 11132 20315 11135
rect 21082 11132 21088 11144
rect 20303 11104 21088 11132
rect 20303 11101 20315 11104
rect 20257 11095 20315 11101
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 23584 11141 23612 11172
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 26234 11160 26240 11212
rect 26292 11200 26298 11212
rect 26329 11203 26387 11209
rect 26329 11200 26341 11203
rect 26292 11172 26341 11200
rect 26292 11160 26298 11172
rect 26329 11169 26341 11172
rect 26375 11169 26387 11203
rect 26602 11200 26608 11212
rect 26563 11172 26608 11200
rect 26329 11163 26387 11169
rect 26602 11160 26608 11172
rect 26660 11160 26666 11212
rect 27632 11200 27660 11308
rect 28353 11203 28411 11209
rect 28353 11200 28365 11203
rect 27632 11172 28365 11200
rect 28353 11169 28365 11172
rect 28399 11169 28411 11203
rect 28353 11163 28411 11169
rect 23569 11135 23627 11141
rect 23569 11101 23581 11135
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 24762 11092 24768 11144
rect 24820 11132 24826 11144
rect 24949 11135 25007 11141
rect 24949 11132 24961 11135
rect 24820 11104 24961 11132
rect 24820 11092 24826 11104
rect 24949 11101 24961 11104
rect 24995 11132 25007 11135
rect 25593 11135 25651 11141
rect 25593 11132 25605 11135
rect 24995 11104 25605 11132
rect 24995 11101 25007 11104
rect 24949 11095 25007 11101
rect 25593 11101 25605 11104
rect 25639 11101 25651 11135
rect 25593 11095 25651 11101
rect 16255 11036 16988 11064
rect 16255 11033 16267 11036
rect 16209 11027 16267 11033
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 21174 11064 21180 11076
rect 17276 11036 21180 11064
rect 17276 11024 17282 11036
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 21692 11036 21737 11064
rect 22020 11036 22126 11064
rect 21692 11024 21698 11036
rect 10870 10996 10876 11008
rect 9232 10968 10876 10996
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 13633 10999 13691 11005
rect 13633 10965 13645 10999
rect 13679 10996 13691 10999
rect 13722 10996 13728 11008
rect 13679 10968 13728 10996
rect 13679 10965 13691 10968
rect 13633 10959 13691 10965
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 17770 10996 17776 11008
rect 13872 10968 17776 10996
rect 13872 10956 13878 10968
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 22020 10996 22048 11036
rect 23934 11024 23940 11076
rect 23992 11064 23998 11076
rect 23992 11036 27094 11064
rect 23992 11024 23998 11036
rect 18012 10968 22048 10996
rect 18012 10956 18018 10968
rect 24210 10956 24216 11008
rect 24268 10996 24274 11008
rect 25685 10999 25743 11005
rect 25685 10996 25697 10999
rect 24268 10968 25697 10996
rect 24268 10956 24274 10968
rect 25685 10965 25697 10968
rect 25731 10965 25743 10999
rect 25685 10959 25743 10965
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 6733 10795 6791 10801
rect 6733 10761 6745 10795
rect 6779 10792 6791 10795
rect 7282 10792 7288 10804
rect 6779 10764 7288 10792
rect 6779 10761 6791 10764
rect 6733 10755 6791 10761
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 9490 10792 9496 10804
rect 9451 10764 9496 10792
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11882 10792 11888 10804
rect 11011 10764 11888 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12802 10792 12808 10804
rect 12763 10764 12808 10792
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13354 10752 13360 10804
rect 13412 10792 13418 10804
rect 16853 10795 16911 10801
rect 13412 10764 14412 10792
rect 13412 10752 13418 10764
rect 13722 10724 13728 10736
rect 13683 10696 13728 10724
rect 13722 10684 13728 10696
rect 13780 10684 13786 10736
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7742 10656 7748 10668
rect 6963 10628 7748 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 11146 10656 11152 10668
rect 11107 10628 11152 10656
rect 9677 10619 9735 10625
rect 9692 10452 9720 10619
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12308 10628 12357 10656
rect 12308 10616 12314 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13446 10656 13452 10668
rect 13035 10628 13452 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 13633 10591 13691 10597
rect 13633 10557 13645 10591
rect 13679 10588 13691 10591
rect 14274 10588 14280 10600
rect 13679 10560 14280 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 14384 10588 14412 10764
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 17218 10792 17224 10804
rect 16899 10764 17224 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 17494 10792 17500 10804
rect 17455 10764 17500 10792
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 21174 10792 21180 10804
rect 17604 10764 21180 10792
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 15565 10727 15623 10733
rect 15565 10724 15577 10727
rect 14875 10696 15577 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 15565 10693 15577 10696
rect 15611 10693 15623 10727
rect 17604 10724 17632 10764
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 21358 10792 21364 10804
rect 21319 10764 21364 10792
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 26602 10792 26608 10804
rect 22388 10764 26608 10792
rect 22388 10736 22416 10764
rect 26602 10752 26608 10764
rect 26660 10752 26666 10804
rect 28261 10795 28319 10801
rect 28261 10761 28273 10795
rect 28307 10792 28319 10795
rect 29914 10792 29920 10804
rect 28307 10764 29920 10792
rect 28307 10761 28319 10764
rect 28261 10755 28319 10761
rect 29914 10752 29920 10764
rect 29972 10752 29978 10804
rect 20254 10724 20260 10736
rect 15565 10687 15623 10693
rect 17144 10696 17632 10724
rect 20215 10696 20260 10724
rect 14734 10656 14740 10668
rect 14695 10628 14740 10656
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 16942 10616 16948 10668
rect 17000 10640 17006 10668
rect 17037 10643 17095 10649
rect 17037 10640 17049 10643
rect 17000 10616 17049 10640
rect 16960 10612 17049 10616
rect 17037 10609 17049 10612
rect 17083 10640 17095 10643
rect 17144 10640 17172 10696
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 22278 10724 22284 10736
rect 22112 10696 22284 10724
rect 17083 10612 17172 10640
rect 17681 10663 17739 10669
rect 17681 10629 17693 10663
rect 17727 10629 17739 10663
rect 17681 10623 17739 10629
rect 17083 10609 17095 10612
rect 17037 10603 17095 10609
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 14384 10560 15485 10588
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17696 10588 17724 10623
rect 19610 10616 19616 10668
rect 19668 10616 19674 10668
rect 21266 10616 21272 10668
rect 21324 10663 21330 10668
rect 22112 10665 22140 10696
rect 22278 10684 22284 10696
rect 22336 10684 22342 10736
rect 22370 10684 22376 10736
rect 22428 10724 22434 10736
rect 22428 10696 22521 10724
rect 22428 10684 22434 10696
rect 24118 10684 24124 10736
rect 24176 10724 24182 10736
rect 24176 10696 25530 10724
rect 24176 10684 24182 10696
rect 21324 10654 21335 10663
rect 22097 10659 22155 10665
rect 21324 10626 21367 10654
rect 21324 10617 21335 10626
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 21324 10616 21330 10617
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 24210 10616 24216 10668
rect 24268 10656 24274 10668
rect 24268 10628 24532 10656
rect 24268 10616 24274 10628
rect 17276 10560 17724 10588
rect 17276 10548 17282 10560
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18230 10588 18236 10600
rect 18104 10560 18236 10588
rect 18104 10548 18110 10560
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 19058 10588 19064 10600
rect 18555 10560 19064 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19242 10548 19248 10600
rect 19300 10588 19306 10600
rect 20530 10588 20536 10600
rect 19300 10560 20536 10588
rect 19300 10548 19306 10560
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 21542 10588 21548 10600
rect 20772 10560 21548 10588
rect 20772 10548 20778 10560
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24504 10597 24532 10628
rect 24578 10616 24584 10668
rect 24636 10656 24642 10668
rect 24765 10659 24823 10665
rect 24765 10656 24777 10659
rect 24636 10628 24777 10656
rect 24636 10616 24642 10628
rect 24765 10625 24777 10628
rect 24811 10625 24823 10659
rect 28074 10656 28080 10668
rect 28035 10628 28080 10656
rect 24765 10619 24823 10625
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 24489 10591 24547 10597
rect 24176 10560 24221 10588
rect 24176 10548 24182 10560
rect 24489 10557 24501 10591
rect 24535 10588 24547 10591
rect 25041 10591 25099 10597
rect 25041 10588 25053 10591
rect 24535 10560 25053 10588
rect 24535 10557 24547 10560
rect 24489 10551 24547 10557
rect 25041 10557 25053 10560
rect 25087 10588 25099 10591
rect 27798 10588 27804 10600
rect 25087 10560 27804 10588
rect 25087 10557 25099 10560
rect 25041 10551 25099 10557
rect 27798 10548 27804 10560
rect 27856 10548 27862 10600
rect 12161 10523 12219 10529
rect 12161 10489 12173 10523
rect 12207 10520 12219 10523
rect 12894 10520 12900 10532
rect 12207 10492 12900 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 14185 10523 14243 10529
rect 14185 10520 14197 10523
rect 13228 10492 14197 10520
rect 13228 10480 13234 10492
rect 14185 10489 14197 10492
rect 14231 10489 14243 10523
rect 16022 10520 16028 10532
rect 15983 10492 16028 10520
rect 14185 10483 14243 10489
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 17954 10520 17960 10532
rect 16540 10492 17960 10520
rect 16540 10480 16546 10492
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 22094 10520 22100 10532
rect 19536 10492 22100 10520
rect 11790 10452 11796 10464
rect 9692 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10452 11854 10464
rect 12710 10452 12716 10464
rect 11848 10424 12716 10452
rect 11848 10412 11854 10424
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 19536 10452 19564 10492
rect 22094 10480 22100 10492
rect 22152 10480 22158 10532
rect 24302 10520 24308 10532
rect 23400 10492 24308 10520
rect 13044 10424 19564 10452
rect 13044 10412 13050 10424
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 23400 10452 23428 10492
rect 24302 10480 24308 10492
rect 24360 10480 24366 10532
rect 20404 10424 23428 10452
rect 20404 10412 20410 10424
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 26510 10452 26516 10464
rect 24268 10424 26516 10452
rect 24268 10412 24274 10424
rect 26510 10412 26516 10424
rect 26568 10412 26574 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 10870 10248 10876 10260
rect 10152 10220 10876 10248
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 3602 10044 3608 10056
rect 1627 10016 3608 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 10152 10044 10180 10220
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 22094 10248 22100 10260
rect 12768 10220 22100 10248
rect 12768 10208 12774 10220
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 24026 10248 24032 10260
rect 23987 10220 24032 10248
rect 24026 10208 24032 10220
rect 24084 10208 24090 10260
rect 25774 10208 25780 10260
rect 25832 10248 25838 10260
rect 26418 10248 26424 10260
rect 25832 10220 26424 10248
rect 25832 10208 25838 10220
rect 26418 10208 26424 10220
rect 26476 10248 26482 10260
rect 26881 10251 26939 10257
rect 26881 10248 26893 10251
rect 26476 10220 26893 10248
rect 26476 10208 26482 10220
rect 26881 10217 26893 10220
rect 26927 10217 26939 10251
rect 26881 10211 26939 10217
rect 10597 10183 10655 10189
rect 10597 10149 10609 10183
rect 10643 10180 10655 10183
rect 17034 10180 17040 10192
rect 10643 10152 17040 10180
rect 10643 10149 10655 10152
rect 10597 10143 10655 10149
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 17129 10183 17187 10189
rect 17129 10149 17141 10183
rect 17175 10180 17187 10183
rect 18138 10180 18144 10192
rect 17175 10152 18144 10180
rect 17175 10149 17187 10152
rect 17129 10143 17187 10149
rect 18138 10140 18144 10152
rect 18196 10140 18202 10192
rect 21376 10152 22232 10180
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10284 10084 11560 10112
rect 10284 10072 10290 10084
rect 10778 10044 10784 10056
rect 9723 10016 10180 10044
rect 10739 10016 10784 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 10928 10016 11253 10044
rect 10928 10004 10934 10016
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11532 10044 11560 10084
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 11756 10084 12725 10112
rect 11756 10072 11762 10084
rect 12713 10081 12725 10084
rect 12759 10081 12771 10115
rect 12713 10075 12771 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 13136 10084 13185 10112
rect 13136 10072 13142 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 16577 10115 16635 10121
rect 16577 10112 16589 10115
rect 15344 10084 16589 10112
rect 15344 10072 15350 10084
rect 16577 10081 16589 10084
rect 16623 10081 16635 10115
rect 17770 10112 17776 10124
rect 17731 10084 17776 10112
rect 16577 10075 16635 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 18104 10084 19809 10112
rect 18104 10072 18110 10084
rect 19797 10081 19809 10084
rect 19843 10112 19855 10115
rect 20622 10112 20628 10124
rect 19843 10084 20628 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 11532 10016 12541 10044
rect 11425 10007 11483 10013
rect 12529 10013 12541 10016
rect 12575 10044 12587 10047
rect 13262 10044 13268 10056
rect 12575 10016 13268 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 11440 9976 11468 10007
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 17218 10004 17224 10056
rect 17276 10044 17282 10056
rect 17402 10044 17408 10056
rect 17276 10016 17408 10044
rect 17276 10004 17282 10016
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 12894 9976 12900 9988
rect 11440 9948 12900 9976
rect 12894 9936 12900 9948
rect 12952 9936 12958 9988
rect 14461 9979 14519 9985
rect 14461 9945 14473 9979
rect 14507 9976 14519 9979
rect 15197 9979 15255 9985
rect 15197 9976 15209 9979
rect 14507 9948 15209 9976
rect 14507 9945 14519 9948
rect 14461 9939 14519 9945
rect 15197 9945 15209 9948
rect 15243 9945 15255 9979
rect 15197 9939 15255 9945
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 15841 9979 15899 9985
rect 15344 9948 15389 9976
rect 15344 9936 15350 9948
rect 15841 9945 15853 9979
rect 15887 9976 15899 9979
rect 15930 9976 15936 9988
rect 15887 9948 15936 9976
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 16669 9979 16727 9985
rect 16669 9945 16681 9979
rect 16715 9945 16727 9979
rect 16669 9939 16727 9945
rect 17865 9979 17923 9985
rect 17865 9945 17877 9979
rect 17911 9945 17923 9979
rect 18414 9976 18420 9988
rect 18375 9948 18420 9976
rect 17865 9939 17923 9945
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 4890 9908 4896 9920
rect 4851 9880 4896 9908
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 9493 9911 9551 9917
rect 9493 9908 9505 9911
rect 9272 9880 9505 9908
rect 9272 9868 9278 9880
rect 9493 9877 9505 9880
rect 9539 9877 9551 9911
rect 9493 9871 9551 9877
rect 11885 9911 11943 9917
rect 11885 9877 11897 9911
rect 11931 9908 11943 9911
rect 14550 9908 14556 9920
rect 11931 9880 14556 9908
rect 11931 9877 11943 9880
rect 11885 9871 11943 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 16684 9908 16712 9939
rect 14792 9880 16712 9908
rect 14792 9868 14798 9880
rect 16942 9868 16948 9920
rect 17000 9908 17006 9920
rect 17880 9908 17908 9939
rect 18414 9936 18420 9948
rect 18472 9936 18478 9988
rect 19334 9976 19340 9988
rect 18892 9948 19340 9976
rect 17000 9880 17908 9908
rect 17000 9868 17006 9880
rect 18322 9868 18328 9920
rect 18380 9908 18386 9920
rect 18892 9908 18920 9948
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 20070 9976 20076 9988
rect 20031 9948 20076 9976
rect 20070 9936 20076 9948
rect 20128 9936 20134 9988
rect 21082 9936 21088 9988
rect 21140 9936 21146 9988
rect 18380 9880 18920 9908
rect 18380 9868 18386 9880
rect 18966 9868 18972 9920
rect 19024 9908 19030 9920
rect 21376 9908 21404 10152
rect 22204 10112 22232 10152
rect 24210 10140 24216 10192
rect 24268 10180 24274 10192
rect 28169 10183 28227 10189
rect 24268 10152 25268 10180
rect 24268 10140 24274 10152
rect 22646 10112 22652 10124
rect 22204 10084 22652 10112
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 24486 10112 24492 10124
rect 23256 10084 24492 10112
rect 23256 10072 23262 10084
rect 24486 10072 24492 10084
rect 24544 10072 24550 10124
rect 24578 10072 24584 10124
rect 24636 10112 24642 10124
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 24636 10084 25145 10112
rect 24636 10072 24642 10084
rect 25133 10081 25145 10084
rect 25179 10081 25191 10115
rect 25240 10112 25268 10152
rect 28169 10149 28181 10183
rect 28215 10149 28227 10183
rect 28169 10143 28227 10149
rect 28184 10112 28212 10143
rect 25240 10084 28212 10112
rect 25133 10075 25191 10081
rect 22278 10044 22284 10056
rect 22239 10016 22284 10044
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 28350 10044 28356 10056
rect 28311 10016 28356 10044
rect 28350 10004 28356 10016
rect 28408 10004 28414 10056
rect 21821 9979 21879 9985
rect 21821 9976 21833 9979
rect 21468 9948 21833 9976
rect 21468 9920 21496 9948
rect 21821 9945 21833 9948
rect 21867 9945 21879 9979
rect 21821 9939 21879 9945
rect 22186 9936 22192 9988
rect 22244 9976 22250 9988
rect 22557 9979 22615 9985
rect 22557 9976 22569 9979
rect 22244 9948 22569 9976
rect 22244 9936 22250 9948
rect 22557 9945 22569 9948
rect 22603 9945 22615 9979
rect 25396 9979 25454 9985
rect 22557 9939 22615 9945
rect 22664 9948 23046 9976
rect 19024 9880 21404 9908
rect 19024 9868 19030 9880
rect 21450 9868 21456 9920
rect 21508 9868 21514 9920
rect 21542 9868 21548 9920
rect 21600 9908 21606 9920
rect 22664 9908 22692 9948
rect 25396 9945 25408 9979
rect 25442 9945 25454 9979
rect 25396 9939 25454 9945
rect 21600 9880 22692 9908
rect 25424 9908 25452 9939
rect 25866 9936 25872 9988
rect 25924 9936 25930 9988
rect 26050 9908 26056 9920
rect 25424 9880 26056 9908
rect 21600 9868 21606 9880
rect 26050 9868 26056 9880
rect 26108 9868 26114 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 3602 9704 3608 9716
rect 3563 9676 3608 9704
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 10965 9707 11023 9713
rect 10965 9704 10977 9707
rect 10836 9676 10977 9704
rect 10836 9664 10842 9676
rect 10965 9673 10977 9676
rect 11011 9673 11023 9707
rect 10965 9667 11023 9673
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 11204 9676 12173 9704
rect 11204 9664 11210 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 12161 9667 12219 9673
rect 13004 9676 14688 9704
rect 12434 9636 12440 9648
rect 9876 9608 12440 9636
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 4890 9568 4896 9580
rect 3835 9540 4896 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 6638 9568 6644 9580
rect 6599 9540 6644 9568
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 8386 9568 8392 9580
rect 8347 9540 8392 9568
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 9214 9568 9220 9580
rect 9175 9540 9220 9568
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9876 9577 9904 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 9861 9531 9919 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 11149 9571 11207 9577
rect 10468 9540 10513 9568
rect 10468 9528 10474 9540
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11164 9500 11192 9531
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 12345 9571 12403 9577
rect 12345 9568 12357 9571
rect 11296 9540 12357 9568
rect 11296 9528 11302 9540
rect 12345 9537 12357 9540
rect 12391 9568 12403 9571
rect 12802 9568 12808 9580
rect 12391 9540 12808 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 13004 9577 13032 9676
rect 14660 9636 14688 9676
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14792 9676 14933 9704
rect 14792 9664 14798 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 18322 9704 18328 9716
rect 14921 9667 14979 9673
rect 15028 9676 18328 9704
rect 15028 9636 15056 9676
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 18472 9676 20024 9704
rect 18472 9664 18478 9676
rect 17218 9636 17224 9648
rect 14660 9608 15056 9636
rect 17053 9608 17224 9636
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13780 9540 13829 9568
rect 13780 9528 13786 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 15102 9568 15108 9580
rect 15063 9540 15108 9568
rect 14461 9531 14519 9537
rect 11974 9500 11980 9512
rect 11164 9472 11980 9500
rect 11974 9460 11980 9472
rect 12032 9500 12038 9512
rect 14476 9500 14504 9531
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15562 9568 15568 9580
rect 15523 9540 15568 9568
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 17053 9577 17081 9608
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 17497 9639 17555 9645
rect 17497 9636 17509 9639
rect 17460 9608 17509 9636
rect 17460 9596 17466 9608
rect 17497 9605 17509 9608
rect 17543 9605 17555 9639
rect 18230 9636 18236 9648
rect 18191 9608 18236 9636
rect 17497 9599 17555 9605
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 19996 9636 20024 9676
rect 20070 9664 20076 9716
rect 20128 9704 20134 9716
rect 20898 9704 20904 9716
rect 20128 9676 20904 9704
rect 20128 9664 20134 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 21266 9704 21272 9716
rect 21008 9676 21272 9704
rect 21008 9636 21036 9676
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 22833 9639 22891 9645
rect 22833 9636 22845 9639
rect 19996 9608 21036 9636
rect 22066 9608 22845 9636
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16724 9540 16865 9568
rect 16724 9528 16730 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17954 9568 17960 9580
rect 17915 9540 17960 9568
rect 17037 9531 17095 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 20254 9568 20260 9580
rect 19366 9540 20260 9568
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20530 9528 20536 9580
rect 20588 9568 20594 9580
rect 22066 9568 22094 9608
rect 22833 9605 22845 9608
rect 22879 9605 22891 9639
rect 25038 9636 25044 9648
rect 24058 9608 25044 9636
rect 22833 9599 22891 9605
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 20588 9540 22094 9568
rect 20588 9528 20594 9540
rect 22278 9528 22284 9580
rect 22336 9568 22342 9580
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22336 9540 22569 9568
rect 22336 9528 22342 9540
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24636 9540 24869 9568
rect 24636 9528 24642 9540
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 24857 9531 24915 9537
rect 26234 9528 26240 9580
rect 26292 9528 26298 9580
rect 27982 9568 27988 9580
rect 26344 9540 27988 9568
rect 17770 9500 17776 9512
rect 12032 9472 12296 9500
rect 14476 9472 17776 9500
rect 12032 9460 12038 9472
rect 9033 9435 9091 9441
rect 9033 9401 9045 9435
rect 9079 9432 9091 9435
rect 9306 9432 9312 9444
rect 9079 9404 9312 9432
rect 9079 9401 9091 9404
rect 9033 9395 9091 9401
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 9677 9435 9735 9441
rect 9677 9401 9689 9435
rect 9723 9401 9735 9435
rect 12268 9432 12296 9472
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 18840 9472 19717 9500
rect 18840 9460 18846 9472
rect 19705 9469 19717 9472
rect 19751 9500 19763 9503
rect 21358 9500 21364 9512
rect 19751 9472 21364 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 22462 9460 22468 9512
rect 22520 9500 22526 9512
rect 25133 9503 25191 9509
rect 22520 9472 24624 9500
rect 22520 9460 22526 9472
rect 13630 9432 13636 9444
rect 12268 9404 13492 9432
rect 13591 9404 13636 9432
rect 9677 9395 9735 9401
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 5960 9336 6745 9364
rect 5960 9324 5966 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9364 8539 9367
rect 8662 9364 8668 9376
rect 8527 9336 8668 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 9692 9364 9720 9395
rect 12618 9364 12624 9376
rect 9692 9336 12624 9364
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 13078 9364 13084 9376
rect 13039 9336 13084 9364
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 13464 9364 13492 9404
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9432 15715 9435
rect 15703 9404 17908 9432
rect 15703 9401 15715 9404
rect 15657 9395 15715 9401
rect 14090 9364 14096 9376
rect 13464 9336 14096 9364
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14277 9367 14335 9373
rect 14277 9333 14289 9367
rect 14323 9364 14335 9367
rect 17126 9364 17132 9376
rect 14323 9336 17132 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17880 9364 17908 9404
rect 20070 9364 20076 9376
rect 17880 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 21450 9364 21456 9376
rect 20680 9336 21456 9364
rect 20680 9324 20686 9336
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 24302 9364 24308 9376
rect 24263 9336 24308 9364
rect 24302 9324 24308 9336
rect 24360 9324 24366 9376
rect 24596 9364 24624 9472
rect 25133 9469 25145 9503
rect 25179 9500 25191 9503
rect 25774 9500 25780 9512
rect 25179 9472 25780 9500
rect 25179 9469 25191 9472
rect 25133 9463 25191 9469
rect 25774 9460 25780 9472
rect 25832 9500 25838 9512
rect 26344 9500 26372 9540
rect 27982 9528 27988 9540
rect 28040 9528 28046 9580
rect 28353 9571 28411 9577
rect 28353 9537 28365 9571
rect 28399 9568 28411 9571
rect 28442 9568 28448 9580
rect 28399 9540 28448 9568
rect 28399 9537 28411 9540
rect 28353 9531 28411 9537
rect 28442 9528 28448 9540
rect 28500 9528 28506 9580
rect 26602 9500 26608 9512
rect 25832 9472 26372 9500
rect 26563 9472 26608 9500
rect 25832 9460 25838 9472
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27890 9392 27896 9444
rect 27948 9432 27954 9444
rect 28169 9435 28227 9441
rect 28169 9432 28181 9435
rect 27948 9404 28181 9432
rect 27948 9392 27954 9404
rect 28169 9401 28181 9404
rect 28215 9401 28227 9435
rect 28169 9395 28227 9401
rect 27614 9364 27620 9376
rect 24596 9336 27620 9364
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 10870 9160 10876 9172
rect 8527 9132 10876 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11698 9160 11704 9172
rect 11379 9132 11704 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 12529 9163 12587 9169
rect 12529 9160 12541 9163
rect 12492 9132 12541 9160
rect 12492 9120 12498 9132
rect 12529 9129 12541 9132
rect 12575 9160 12587 9163
rect 13354 9160 13360 9172
rect 12575 9132 13360 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 15102 9160 15108 9172
rect 13688 9132 15108 9160
rect 13688 9120 13694 9132
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 24302 9160 24308 9172
rect 18104 9132 24308 9160
rect 18104 9120 18110 9132
rect 24302 9120 24308 9132
rect 24360 9120 24366 9172
rect 24673 9163 24731 9169
rect 24673 9129 24685 9163
rect 24719 9129 24731 9163
rect 24673 9123 24731 9129
rect 12158 9092 12164 9104
rect 1596 9064 12164 9092
rect 1596 8965 1624 9064
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 14645 9095 14703 9101
rect 14645 9092 14657 9095
rect 14240 9064 14657 9092
rect 14240 9052 14246 9064
rect 14645 9061 14657 9064
rect 14691 9061 14703 9095
rect 14645 9055 14703 9061
rect 14734 9052 14740 9104
rect 14792 9092 14798 9104
rect 16758 9092 16764 9104
rect 14792 9064 16764 9092
rect 14792 9052 14798 9064
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 19150 9052 19156 9104
rect 19208 9092 19214 9104
rect 19208 9064 21128 9092
rect 19208 9052 19214 9064
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 7837 9027 7895 9033
rect 4120 8996 7788 9024
rect 4120 8984 4126 8996
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 5902 8956 5908 8968
rect 5863 8928 5908 8956
rect 1581 8919 1639 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 7760 8965 7788 8996
rect 7837 8993 7849 9027
rect 7883 9024 7895 9027
rect 9953 9027 10011 9033
rect 9953 9024 9965 9027
rect 7883 8996 9965 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 9953 8993 9965 8996
rect 9999 8993 10011 9027
rect 9953 8987 10011 8993
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 12069 9027 12127 9033
rect 12069 9024 12081 9027
rect 10652 8996 12081 9024
rect 10652 8984 10658 8996
rect 12069 8993 12081 8996
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 14461 9027 14519 9033
rect 14461 9024 14473 9027
rect 13044 8996 14473 9024
rect 13044 8984 13050 8996
rect 14461 8993 14473 8996
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16206 9024 16212 9036
rect 16071 8996 16212 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 9024 17187 9027
rect 17954 9024 17960 9036
rect 17175 8996 17960 9024
rect 17175 8993 17187 8996
rect 17129 8987 17187 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18414 8984 18420 9036
rect 18472 9024 18478 9036
rect 18472 8996 19334 9024
rect 18472 8984 18478 8996
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8478 8956 8484 8968
rect 8435 8928 8484 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 9306 8956 9312 8968
rect 9267 8928 9312 8956
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9416 8928 10149 8956
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9416 8888 9444 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 11238 8956 11244 8968
rect 11199 8928 11244 8956
rect 10137 8919 10195 8925
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 11974 8956 11980 8968
rect 11931 8928 11980 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13504 8928 13553 8956
rect 13504 8916 13510 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 13541 8919 13599 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 19306 8956 19334 8996
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 20993 9027 21051 9033
rect 20993 9024 21005 9027
rect 20772 8996 21005 9024
rect 20772 8984 20778 8996
rect 20993 8993 21005 8996
rect 21039 8993 21051 9027
rect 21100 9024 21128 9064
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 24688 9092 24716 9123
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 28258 9160 28264 9172
rect 24912 9132 28264 9160
rect 24912 9120 24918 9132
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 23164 9064 24716 9092
rect 23164 9052 23170 9064
rect 21358 9024 21364 9036
rect 21100 8996 21364 9024
rect 20993 8987 21051 8993
rect 21358 8984 21364 8996
rect 21416 8984 21422 9036
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 22462 9024 22468 9036
rect 21692 8996 22468 9024
rect 21692 8984 21698 8996
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 22741 9027 22799 9033
rect 22741 8993 22753 9027
rect 22787 9024 22799 9027
rect 23842 9024 23848 9036
rect 22787 8996 23848 9024
rect 22787 8993 22799 8996
rect 22741 8987 22799 8993
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 24670 8984 24676 9036
rect 24728 9024 24734 9036
rect 26053 9027 26111 9033
rect 26053 9024 26065 9027
rect 24728 8996 26065 9024
rect 24728 8984 24734 8996
rect 26053 8993 26065 8996
rect 26099 8993 26111 9027
rect 26053 8987 26111 8993
rect 26329 9027 26387 9033
rect 26329 8993 26341 9027
rect 26375 9024 26387 9027
rect 26418 9024 26424 9036
rect 26375 8996 26424 9024
rect 26375 8993 26387 8996
rect 26329 8987 26387 8993
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 27614 8984 27620 9036
rect 27672 9024 27678 9036
rect 28077 9027 28135 9033
rect 28077 9024 28089 9027
rect 27672 8996 28089 9024
rect 27672 8984 27678 8996
rect 28077 8993 28089 8996
rect 28123 8993 28135 9027
rect 28077 8987 28135 8993
rect 20806 8956 20812 8968
rect 19306 8928 20812 8956
rect 20806 8916 20812 8928
rect 20864 8916 20870 8968
rect 22370 8916 22376 8968
rect 22428 8916 22434 8968
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 23290 8956 23296 8968
rect 22888 8928 23296 8956
rect 22888 8916 22894 8928
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 24762 8956 24768 8968
rect 24627 8928 24768 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 24762 8916 24768 8928
rect 24820 8956 24826 8968
rect 25225 8959 25283 8965
rect 25225 8956 25237 8959
rect 24820 8928 25237 8956
rect 24820 8916 24826 8928
rect 25225 8925 25237 8928
rect 25271 8925 25283 8959
rect 25225 8919 25283 8925
rect 8352 8860 9444 8888
rect 8352 8848 8358 8860
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 12802 8888 12808 8900
rect 9916 8860 12808 8888
rect 9916 8848 9922 8860
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 13633 8891 13691 8897
rect 13633 8857 13645 8891
rect 13679 8888 13691 8891
rect 13679 8860 16068 8888
rect 13679 8857 13691 8860
rect 13633 8851 13691 8857
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 1762 8820 1768 8832
rect 1719 8792 1768 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 5718 8820 5724 8832
rect 5679 8792 5724 8820
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 9401 8823 9459 8829
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 10410 8820 10416 8832
rect 9447 8792 10416 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10597 8823 10655 8829
rect 10597 8789 10609 8823
rect 10643 8820 10655 8823
rect 11238 8820 11244 8832
rect 10643 8792 11244 8820
rect 10643 8789 10655 8792
rect 10597 8783 10655 8789
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 14734 8820 14740 8832
rect 13964 8792 14740 8820
rect 13964 8780 13970 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 16040 8820 16068 8860
rect 16114 8848 16120 8900
rect 16172 8888 16178 8900
rect 16669 8891 16727 8897
rect 16172 8860 16217 8888
rect 16172 8848 16178 8860
rect 16669 8857 16681 8891
rect 16715 8857 16727 8891
rect 17402 8888 17408 8900
rect 17363 8860 17408 8888
rect 16669 8851 16727 8857
rect 16390 8820 16396 8832
rect 16040 8792 16396 8820
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 16684 8820 16712 8851
rect 17402 8848 17408 8860
rect 17460 8848 17466 8900
rect 21174 8888 21180 8900
rect 18630 8860 21180 8888
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 21269 8891 21327 8897
rect 21269 8857 21281 8891
rect 21315 8857 21327 8891
rect 21269 8851 21327 8857
rect 18138 8820 18144 8832
rect 16684 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 18877 8823 18935 8829
rect 18877 8820 18889 8823
rect 18840 8792 18889 8820
rect 18840 8780 18846 8792
rect 18877 8789 18889 8792
rect 18923 8820 18935 8823
rect 20530 8820 20536 8832
rect 18923 8792 20536 8820
rect 18923 8789 18935 8792
rect 18877 8783 18935 8789
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 20622 8780 20628 8832
rect 20680 8820 20686 8832
rect 21284 8820 21312 8851
rect 22554 8848 22560 8900
rect 22612 8888 22618 8900
rect 23385 8891 23443 8897
rect 22612 8860 23336 8888
rect 22612 8848 22618 8860
rect 20680 8792 21312 8820
rect 23308 8820 23336 8860
rect 23385 8857 23397 8891
rect 23431 8888 23443 8891
rect 25130 8888 25136 8900
rect 23431 8860 25136 8888
rect 23431 8857 23443 8860
rect 23385 8851 23443 8857
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 26786 8848 26792 8900
rect 26844 8848 26850 8900
rect 25317 8823 25375 8829
rect 25317 8820 25329 8823
rect 23308 8792 25329 8820
rect 20680 8780 20686 8792
rect 25317 8789 25329 8792
rect 25363 8789 25375 8823
rect 25317 8783 25375 8789
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8294 8616 8300 8628
rect 8251 8588 8300 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 9398 8616 9404 8628
rect 9359 8588 9404 8616
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 13630 8616 13636 8628
rect 9548 8588 13636 8616
rect 9548 8576 9554 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16114 8616 16120 8628
rect 15979 8588 16120 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 20073 8619 20131 8625
rect 17828 8588 20024 8616
rect 17828 8576 17834 8588
rect 11974 8548 11980 8560
rect 9646 8520 11980 8548
rect 1762 8480 1768 8492
rect 1723 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8128 8344 8156 8443
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8755 8483 8813 8489
rect 8755 8480 8767 8483
rect 8720 8452 8767 8480
rect 8720 8440 8726 8452
rect 8755 8449 8767 8452
rect 8801 8480 8813 8483
rect 9646 8480 9674 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 12483 8520 13032 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 9858 8480 9864 8492
rect 8801 8452 9674 8480
rect 9819 8452 9864 8480
rect 8801 8449 8813 8452
rect 8755 8443 8813 8449
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10468 8452 10701 8480
rect 10468 8440 10474 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8480 11207 8483
rect 13004 8480 13032 8520
rect 13078 8508 13084 8560
rect 13136 8548 13142 8560
rect 14553 8551 14611 8557
rect 14553 8548 14565 8551
rect 13136 8520 14565 8548
rect 13136 8508 13142 8520
rect 14553 8517 14565 8520
rect 14599 8517 14611 8551
rect 14553 8511 14611 8517
rect 14826 8508 14832 8560
rect 14884 8548 14890 8560
rect 17402 8548 17408 8560
rect 14884 8520 17408 8548
rect 14884 8508 14890 8520
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 17954 8548 17960 8560
rect 17788 8520 17960 8548
rect 13170 8480 13176 8492
rect 11195 8452 12434 8480
rect 13004 8452 13176 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 8938 8412 8944 8424
rect 8899 8384 8944 8412
rect 8938 8372 8944 8384
rect 8996 8372 9002 8424
rect 10134 8372 10140 8424
rect 10192 8412 10198 8424
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 10192 8384 10517 8412
rect 10192 8372 10198 8384
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 10836 8384 11805 8412
rect 10836 8372 10842 8384
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8381 12035 8415
rect 12406 8412 12434 8452
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13814 8480 13820 8492
rect 13311 8452 13820 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 13906 8440 13912 8492
rect 13964 8480 13970 8492
rect 13964 8452 14009 8480
rect 13964 8440 13970 8452
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 15654 8480 15660 8492
rect 15252 8452 15660 8480
rect 15252 8440 15258 8452
rect 15654 8440 15660 8452
rect 15712 8480 15718 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15712 8452 15853 8480
rect 15712 8440 15718 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 15841 8443 15899 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17788 8489 17816 8520
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 19996 8548 20024 8588
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20346 8616 20352 8628
rect 20119 8588 20352 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 21634 8616 21640 8628
rect 20772 8588 21640 8616
rect 20772 8576 20778 8588
rect 21634 8576 21640 8588
rect 21692 8616 21698 8628
rect 22002 8616 22008 8628
rect 21692 8588 22008 8616
rect 21692 8576 21698 8588
rect 22002 8576 22008 8588
rect 22060 8616 22066 8628
rect 24118 8616 24124 8628
rect 22060 8588 24124 8616
rect 22060 8576 22066 8588
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 28074 8616 28080 8628
rect 28035 8588 28080 8616
rect 28074 8576 28080 8588
rect 28132 8576 28138 8628
rect 19996 8520 21220 8548
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 14182 8412 14188 8424
rect 12406 8384 14188 8412
rect 11977 8375 12035 8381
rect 8754 8344 8760 8356
rect 8128 8316 8760 8344
rect 8754 8304 8760 8316
rect 8812 8344 8818 8356
rect 9306 8344 9312 8356
rect 8812 8316 9312 8344
rect 8812 8304 8818 8316
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9953 8347 10011 8353
rect 9953 8313 9965 8347
rect 9999 8344 10011 8347
rect 11992 8344 12020 8375
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14461 8415 14519 8421
rect 14461 8381 14473 8415
rect 14507 8412 14519 8415
rect 14507 8384 14688 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 9999 8316 12020 8344
rect 13081 8347 13139 8353
rect 9999 8313 10011 8316
rect 9953 8307 10011 8313
rect 13081 8313 13093 8347
rect 13127 8344 13139 8347
rect 13538 8344 13544 8356
rect 13127 8316 13544 8344
rect 13127 8313 13139 8316
rect 13081 8307 13139 8313
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14660 8344 14688 8384
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 14792 8384 14837 8412
rect 14792 8372 14798 8384
rect 17218 8372 17224 8424
rect 17276 8412 17282 8424
rect 18046 8412 18052 8424
rect 17276 8384 18052 8412
rect 17276 8372 17282 8384
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 19168 8412 19196 8466
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19484 8452 19993 8480
rect 19484 8440 19490 8452
rect 19981 8449 19993 8452
rect 20027 8480 20039 8483
rect 20346 8480 20352 8492
rect 20027 8452 20352 8480
rect 20027 8449 20039 8452
rect 19981 8443 20039 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20714 8480 20720 8492
rect 20671 8452 20720 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 20806 8440 20812 8492
rect 20864 8440 20870 8492
rect 21192 8484 21220 8520
rect 21450 8508 21456 8560
rect 21508 8548 21514 8560
rect 22186 8548 22192 8560
rect 21508 8520 22192 8548
rect 21508 8508 21514 8520
rect 22186 8508 22192 8520
rect 22244 8508 22250 8560
rect 22830 8508 22836 8560
rect 22888 8508 22894 8560
rect 25314 8508 25320 8560
rect 25372 8508 25378 8560
rect 26326 8508 26332 8560
rect 26384 8548 26390 8560
rect 26605 8551 26663 8557
rect 26605 8548 26617 8551
rect 26384 8520 26617 8548
rect 26384 8508 26390 8520
rect 26605 8517 26617 8520
rect 26651 8517 26663 8551
rect 26605 8511 26663 8517
rect 21269 8484 21327 8489
rect 21192 8483 21327 8484
rect 21192 8456 21281 8483
rect 21269 8449 21281 8456
rect 21315 8478 21327 8483
rect 21358 8478 21364 8492
rect 21315 8450 21364 8478
rect 21315 8449 21327 8450
rect 21269 8443 21327 8449
rect 21358 8440 21364 8450
rect 21416 8440 21422 8492
rect 22002 8480 22008 8492
rect 21963 8452 22008 8480
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 28258 8480 28264 8492
rect 28219 8452 28264 8480
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 19242 8412 19248 8424
rect 19168 8384 19248 8412
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8412 19579 8415
rect 19702 8412 19708 8424
rect 19567 8384 19708 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 19702 8372 19708 8384
rect 19760 8372 19766 8424
rect 20824 8412 20852 8440
rect 21450 8412 21456 8424
rect 20824 8384 21456 8412
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8412 22339 8415
rect 22646 8412 22652 8424
rect 22327 8384 22652 8412
rect 22327 8381 22339 8384
rect 22281 8375 22339 8381
rect 22646 8372 22652 8384
rect 22704 8372 22710 8424
rect 24578 8372 24584 8424
rect 24636 8412 24642 8424
rect 24857 8415 24915 8421
rect 24636 8384 24681 8412
rect 24636 8372 24642 8384
rect 24857 8381 24869 8415
rect 24903 8412 24915 8415
rect 26510 8412 26516 8424
rect 24903 8384 26516 8412
rect 24903 8381 24915 8384
rect 24857 8375 24915 8381
rect 26510 8372 26516 8384
rect 26568 8372 26574 8424
rect 20162 8344 20168 8356
rect 13780 8316 13825 8344
rect 14660 8316 17908 8344
rect 13780 8304 13786 8316
rect 1578 8276 1584 8288
rect 1539 8248 1584 8276
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7561 8279 7619 8285
rect 7561 8276 7573 8279
rect 6972 8248 7573 8276
rect 6972 8236 6978 8248
rect 7561 8245 7573 8248
rect 7607 8245 7619 8279
rect 7561 8239 7619 8245
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 14366 8276 14372 8288
rect 9824 8248 14372 8276
rect 9824 8236 9830 8248
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 14734 8276 14740 8288
rect 14516 8248 14740 8276
rect 14516 8236 14522 8248
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 17880 8276 17908 8316
rect 19076 8316 20168 8344
rect 19076 8276 19104 8316
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 20714 8344 20720 8356
rect 20675 8316 20720 8344
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 20806 8304 20812 8356
rect 20864 8344 20870 8356
rect 21361 8347 21419 8353
rect 21361 8344 21373 8347
rect 20864 8316 21373 8344
rect 20864 8304 20870 8316
rect 21361 8313 21373 8316
rect 21407 8313 21419 8347
rect 23750 8344 23756 8356
rect 23711 8316 23756 8344
rect 21361 8307 21419 8313
rect 23750 8304 23756 8316
rect 23808 8304 23814 8356
rect 17880 8248 19104 8276
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 21542 8276 21548 8288
rect 19392 8248 21548 8276
rect 19392 8236 19398 8248
rect 21542 8236 21548 8248
rect 21600 8276 21606 8288
rect 23382 8276 23388 8288
rect 21600 8248 23388 8276
rect 21600 8236 21606 8248
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 8938 8072 8944 8084
rect 7883 8044 8944 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 11790 8072 11796 8084
rect 9416 8044 11796 8072
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 8294 8004 8300 8016
rect 1627 7976 8300 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 9416 7936 9444 8044
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 15286 8072 15292 8084
rect 12483 8044 15292 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 17218 8032 17224 8084
rect 17276 8072 17282 8084
rect 23382 8072 23388 8084
rect 17276 8044 23244 8072
rect 23343 8044 23388 8072
rect 17276 8032 17282 8044
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 8004 10011 8007
rect 12710 8004 12716 8016
rect 9999 7976 12716 8004
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 12710 7964 12716 7976
rect 12768 7964 12774 8016
rect 14366 7964 14372 8016
rect 14424 8004 14430 8016
rect 19334 8004 19340 8016
rect 14424 7976 19340 8004
rect 14424 7964 14430 7976
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 21177 8007 21235 8013
rect 21177 7973 21189 8007
rect 21223 8004 21235 8007
rect 21450 8004 21456 8016
rect 21223 7976 21456 8004
rect 21223 7973 21235 7976
rect 21177 7967 21235 7973
rect 21450 7964 21456 7976
rect 21508 8004 21514 8016
rect 23216 8004 23244 8044
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 23750 8032 23756 8084
rect 23808 8072 23814 8084
rect 26050 8072 26056 8084
rect 23808 8044 26056 8072
rect 23808 8032 23814 8044
rect 26050 8032 26056 8044
rect 26108 8032 26114 8084
rect 27798 8032 27804 8084
rect 27856 8072 27862 8084
rect 28261 8075 28319 8081
rect 28261 8072 28273 8075
rect 27856 8044 28273 8072
rect 27856 8032 27862 8044
rect 28261 8041 28273 8044
rect 28307 8041 28319 8075
rect 28261 8035 28319 8041
rect 24854 8004 24860 8016
rect 21508 7976 21772 8004
rect 23216 7976 24860 8004
rect 21508 7964 21514 7976
rect 7116 7908 9444 7936
rect 9600 7908 10732 7936
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6914 7868 6920 7880
rect 6687 7840 6920 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7116 7877 7144 7908
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7742 7868 7748 7880
rect 7703 7840 7748 7868
rect 7101 7831 7159 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 8570 7868 8576 7880
rect 8531 7840 8576 7868
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 9490 7868 9496 7880
rect 9451 7840 9496 7868
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9600 7800 9628 7908
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10192 7840 10237 7868
rect 10192 7828 10198 7840
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 10597 7871 10655 7877
rect 10597 7868 10609 7871
rect 10560 7840 10609 7868
rect 10560 7828 10566 7840
rect 10597 7837 10609 7840
rect 10643 7837 10655 7871
rect 10704 7868 10732 7908
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 13446 7936 13452 7948
rect 11296 7908 11341 7936
rect 12406 7908 13452 7936
rect 11296 7896 11302 7908
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 10704 7840 10793 7868
rect 10597 7831 10655 7837
rect 10781 7837 10793 7840
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 12406 7868 12434 7908
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 14274 7936 14280 7948
rect 13587 7908 14280 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7936 16359 7939
rect 17034 7936 17040 7948
rect 16347 7908 17040 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 17862 7936 17868 7948
rect 17184 7908 17868 7936
rect 17184 7896 17190 7908
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18138 7936 18144 7948
rect 18012 7908 18144 7936
rect 18012 7896 18018 7908
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 19150 7896 19156 7948
rect 19208 7936 19214 7948
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 19208 7908 19441 7936
rect 19208 7896 19214 7908
rect 19429 7905 19441 7908
rect 19475 7936 19487 7939
rect 21634 7936 21640 7948
rect 19475 7908 21640 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 21744 7936 21772 7976
rect 24854 7964 24860 7976
rect 24912 7964 24918 8016
rect 21913 7939 21971 7945
rect 21913 7936 21925 7939
rect 21744 7908 21925 7936
rect 21913 7905 21925 7908
rect 21959 7905 21971 7939
rect 21913 7899 21971 7905
rect 22278 7896 22284 7948
rect 22336 7936 22342 7948
rect 22336 7908 23244 7936
rect 22336 7896 22342 7908
rect 12618 7868 12624 7880
rect 11839 7840 12434 7868
rect 12579 7840 12624 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 8404 7772 9628 7800
rect 10612 7772 13676 7800
rect 6454 7732 6460 7744
rect 6415 7704 6460 7732
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 8404 7741 8432 7772
rect 7193 7735 7251 7741
rect 7193 7732 7205 7735
rect 6604 7704 7205 7732
rect 6604 7692 6610 7704
rect 7193 7701 7205 7704
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 8389 7735 8447 7741
rect 8389 7701 8401 7735
rect 8435 7701 8447 7735
rect 8389 7695 8447 7701
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 10612 7732 10640 7772
rect 9355 7704 10640 7732
rect 11885 7735 11943 7741
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 11885 7701 11897 7735
rect 11931 7732 11943 7735
rect 12158 7732 12164 7744
rect 11931 7704 12164 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 13648 7732 13676 7772
rect 14182 7760 14188 7812
rect 14240 7800 14246 7812
rect 14829 7803 14887 7809
rect 14829 7800 14841 7803
rect 14240 7772 14841 7800
rect 14240 7760 14246 7772
rect 14829 7769 14841 7772
rect 14875 7769 14887 7803
rect 14829 7763 14887 7769
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 15473 7803 15531 7809
rect 15473 7769 15485 7803
rect 15519 7800 15531 7803
rect 16114 7800 16120 7812
rect 15519 7772 16120 7800
rect 15519 7769 15531 7772
rect 15473 7763 15531 7769
rect 14936 7732 14964 7763
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 16390 7760 16396 7812
rect 16448 7800 16454 7812
rect 16448 7772 16493 7800
rect 16448 7760 16454 7772
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 16945 7803 17003 7809
rect 16945 7800 16957 7803
rect 16724 7772 16957 7800
rect 16724 7760 16730 7772
rect 16945 7769 16957 7772
rect 16991 7769 17003 7803
rect 17862 7800 17868 7812
rect 17823 7772 17868 7800
rect 16945 7763 17003 7769
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 17957 7803 18015 7809
rect 17957 7769 17969 7803
rect 18003 7769 18015 7803
rect 19702 7800 19708 7812
rect 19663 7772 19708 7800
rect 17957 7763 18015 7769
rect 13648 7704 14964 7732
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 17972 7732 18000 7763
rect 19702 7760 19708 7772
rect 19760 7760 19766 7812
rect 19794 7760 19800 7812
rect 19852 7800 19858 7812
rect 23216 7800 23244 7908
rect 23290 7896 23296 7948
rect 23348 7936 23354 7948
rect 23348 7908 23980 7936
rect 23348 7896 23354 7908
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 23845 7871 23903 7877
rect 23845 7868 23857 7871
rect 23808 7840 23857 7868
rect 23808 7828 23814 7840
rect 23845 7837 23857 7840
rect 23891 7837 23903 7871
rect 23952 7868 23980 7908
rect 24118 7896 24124 7948
rect 24176 7936 24182 7948
rect 24578 7936 24584 7948
rect 24176 7908 24584 7936
rect 24176 7896 24182 7908
rect 24578 7896 24584 7908
rect 24636 7936 24642 7948
rect 26513 7939 26571 7945
rect 26513 7936 26525 7939
rect 24636 7908 26525 7936
rect 24636 7896 24642 7908
rect 26513 7905 26525 7908
rect 26559 7905 26571 7939
rect 26513 7899 26571 7905
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 23952 7840 24777 7868
rect 23845 7831 23903 7837
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 25958 7800 25964 7812
rect 19852 7772 20194 7800
rect 21008 7772 21312 7800
rect 19852 7760 19858 7772
rect 16632 7704 18000 7732
rect 16632 7692 16638 7704
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 21008 7732 21036 7772
rect 18104 7704 21036 7732
rect 21284 7732 21312 7772
rect 22020 7772 22402 7800
rect 23216 7772 25964 7800
rect 22020 7732 22048 7772
rect 25958 7760 25964 7772
rect 26016 7760 26022 7812
rect 26786 7800 26792 7812
rect 26747 7772 26792 7800
rect 26786 7760 26792 7772
rect 26844 7760 26850 7812
rect 27798 7760 27804 7812
rect 27856 7760 27862 7812
rect 21284 7704 22048 7732
rect 18104 7692 18110 7704
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 23937 7735 23995 7741
rect 23937 7732 23949 7735
rect 22336 7704 23949 7732
rect 22336 7692 22342 7704
rect 23937 7701 23949 7704
rect 23983 7701 23995 7735
rect 23937 7695 23995 7701
rect 24581 7735 24639 7741
rect 24581 7701 24593 7735
rect 24627 7732 24639 7735
rect 26050 7732 26056 7744
rect 24627 7704 26056 7732
rect 24627 7701 24639 7704
rect 24581 7695 24639 7701
rect 26050 7692 26056 7704
rect 26108 7692 26114 7744
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 12345 7531 12403 7537
rect 12345 7497 12357 7531
rect 12391 7528 12403 7531
rect 12434 7528 12440 7540
rect 12391 7500 12440 7528
rect 12391 7497 12403 7500
rect 12345 7491 12403 7497
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 17678 7528 17684 7540
rect 13504 7500 17684 7528
rect 13504 7488 13510 7500
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 18417 7531 18475 7537
rect 18417 7528 18429 7531
rect 17920 7500 18429 7528
rect 17920 7488 17926 7500
rect 18417 7497 18429 7500
rect 18463 7497 18475 7531
rect 20898 7528 20904 7540
rect 18417 7491 18475 7497
rect 18524 7500 20760 7528
rect 20859 7500 20904 7528
rect 8478 7460 8484 7472
rect 8439 7432 8484 7460
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 8662 7420 8668 7472
rect 8720 7460 8726 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 8720 7432 10425 7460
rect 8720 7420 8726 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10413 7423 10471 7429
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 15657 7463 15715 7469
rect 15657 7460 15669 7463
rect 11296 7432 15669 7460
rect 11296 7420 11302 7432
rect 15657 7429 15669 7432
rect 15703 7429 15715 7463
rect 15657 7423 15715 7429
rect 15746 7420 15752 7472
rect 15804 7460 15810 7472
rect 15804 7432 15849 7460
rect 15804 7420 15810 7432
rect 16114 7420 16120 7472
rect 16172 7460 16178 7472
rect 16301 7463 16359 7469
rect 16301 7460 16313 7463
rect 16172 7432 16313 7460
rect 16172 7420 16178 7432
rect 16301 7429 16313 7432
rect 16347 7460 16359 7463
rect 18524 7460 18552 7500
rect 16347 7432 18552 7460
rect 16347 7429 16359 7432
rect 16301 7423 16359 7429
rect 18782 7420 18788 7472
rect 18840 7460 18846 7472
rect 20732 7460 20760 7500
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 21692 7500 22876 7528
rect 21692 7488 21698 7500
rect 22738 7460 22744 7472
rect 18840 7432 19918 7460
rect 20732 7432 22744 7460
rect 18840 7420 18846 7432
rect 22738 7420 22744 7432
rect 22796 7420 22802 7472
rect 22848 7460 22876 7500
rect 22922 7488 22928 7540
rect 22980 7528 22986 7540
rect 23293 7531 23351 7537
rect 23293 7528 23305 7531
rect 22980 7500 23305 7528
rect 22980 7488 22986 7500
rect 23293 7497 23305 7500
rect 23339 7497 23351 7531
rect 25869 7531 25927 7537
rect 25869 7528 25881 7531
rect 23293 7491 23351 7497
rect 23400 7500 25881 7528
rect 23400 7460 23428 7500
rect 25869 7497 25881 7500
rect 25915 7497 25927 7531
rect 25869 7491 25927 7497
rect 27617 7531 27675 7537
rect 27617 7497 27629 7531
rect 27663 7528 27675 7531
rect 28258 7528 28264 7540
rect 27663 7500 28264 7528
rect 27663 7497 27675 7500
rect 27617 7491 27675 7497
rect 28258 7488 28264 7500
rect 28316 7488 28322 7540
rect 22848 7432 23428 7460
rect 24854 7420 24860 7472
rect 24912 7420 24918 7472
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 9766 7392 9772 7404
rect 9727 7364 9772 7392
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11112 7364 11897 7392
rect 11112 7352 11118 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 12216 7364 14473 7392
rect 12216 7352 12222 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 18690 7392 18696 7404
rect 18003 7364 18696 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 21358 7352 21364 7404
rect 21416 7392 21422 7404
rect 22646 7392 22652 7404
rect 21416 7364 22652 7392
rect 21416 7352 21422 7364
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 23198 7392 23204 7404
rect 23159 7364 23204 7392
rect 23198 7352 23204 7364
rect 23256 7392 23262 7404
rect 23474 7392 23480 7404
rect 23256 7364 23480 7392
rect 23256 7352 23262 7364
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 24118 7392 24124 7404
rect 24079 7364 24124 7392
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 27525 7395 27583 7401
rect 27525 7361 27537 7395
rect 27571 7361 27583 7395
rect 28166 7392 28172 7404
rect 28127 7364 28172 7392
rect 27525 7355 27583 7361
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 7699 7296 8401 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7324 10379 7327
rect 11698 7324 11704 7336
rect 10367 7296 11560 7324
rect 11659 7296 11704 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 8680 7256 8708 7287
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 6880 7228 10885 7256
rect 6880 7216 6886 7228
rect 10873 7225 10885 7228
rect 10919 7225 10931 7259
rect 11532 7256 11560 7296
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12032 7296 13001 7324
rect 12032 7284 12038 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 11790 7256 11796 7268
rect 11532 7228 11796 7256
rect 10873 7219 10931 7225
rect 11790 7216 11796 7228
rect 11848 7216 11854 7268
rect 11882 7216 11888 7268
rect 11940 7256 11946 7268
rect 13188 7256 13216 7287
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13320 7296 14289 7324
rect 13320 7284 13326 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 16298 7324 16304 7336
rect 14700 7296 16304 7324
rect 14700 7284 14706 7296
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 16908 7296 17325 7324
rect 16908 7284 16914 7296
rect 17313 7293 17325 7296
rect 17359 7324 17371 7327
rect 17402 7324 17408 7336
rect 17359 7296 17408 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 18230 7324 18236 7336
rect 17543 7296 18236 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18340 7296 19441 7324
rect 18340 7256 18368 7296
rect 19429 7293 19441 7296
rect 19475 7324 19487 7327
rect 21634 7324 21640 7336
rect 19475 7296 21640 7324
rect 19475 7293 19487 7296
rect 19429 7287 19487 7293
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 22097 7327 22155 7333
rect 22097 7293 22109 7327
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 23566 7324 23572 7336
rect 22327 7296 23572 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 22112 7256 22140 7287
rect 23566 7284 23572 7296
rect 23624 7284 23630 7336
rect 24394 7324 24400 7336
rect 24355 7296 24400 7324
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 24854 7284 24860 7336
rect 24912 7324 24918 7336
rect 27540 7324 27568 7355
rect 28166 7352 28172 7364
rect 28224 7352 28230 7404
rect 24912 7296 27568 7324
rect 24912 7284 24918 7296
rect 24118 7256 24124 7268
rect 11940 7228 13216 7256
rect 13280 7228 18368 7256
rect 20456 7228 21036 7256
rect 22112 7228 24124 7256
rect 11940 7216 11946 7228
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7188 9643 7191
rect 10778 7188 10784 7200
rect 9631 7160 10784 7188
rect 9631 7157 9643 7160
rect 9585 7151 9643 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 12434 7188 12440 7200
rect 11296 7160 12440 7188
rect 11296 7148 11302 7160
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12802 7188 12808 7200
rect 12676 7160 12808 7188
rect 12676 7148 12682 7160
rect 12802 7148 12808 7160
rect 12860 7188 12866 7200
rect 13280 7188 13308 7228
rect 13630 7188 13636 7200
rect 12860 7160 13308 7188
rect 13591 7160 13636 7188
rect 12860 7148 12866 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15654 7148 15660 7200
rect 15712 7188 15718 7200
rect 18874 7188 18880 7200
rect 15712 7160 18880 7188
rect 15712 7148 15718 7160
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 20456 7188 20484 7228
rect 19208 7160 20484 7188
rect 21008 7188 21036 7228
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 22465 7191 22523 7197
rect 22465 7188 22477 7191
rect 21008 7160 22477 7188
rect 19208 7148 19214 7160
rect 22465 7157 22477 7160
rect 22511 7157 22523 7191
rect 22465 7151 22523 7157
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 28261 7191 28319 7197
rect 28261 7188 28273 7191
rect 27672 7160 28273 7188
rect 27672 7148 27678 7160
rect 28261 7157 28273 7160
rect 28307 7157 28319 7191
rect 28261 7151 28319 7157
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 8570 6984 8576 6996
rect 8435 6956 8576 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 8570 6944 8576 6956
rect 8628 6944 8634 6996
rect 11238 6984 11244 6996
rect 8772 6956 11244 6984
rect 7650 6876 7656 6928
rect 7708 6916 7714 6928
rect 8772 6916 8800 6956
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11425 6987 11483 6993
rect 11425 6953 11437 6987
rect 11471 6984 11483 6987
rect 11698 6984 11704 6996
rect 11471 6956 11704 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 14458 6984 14464 6996
rect 11848 6956 14464 6984
rect 11848 6944 11854 6956
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 18288 6956 18429 6984
rect 18288 6944 18294 6956
rect 18417 6953 18429 6956
rect 18463 6953 18475 6987
rect 18417 6947 18475 6953
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 20070 6984 20076 6996
rect 18564 6956 20076 6984
rect 18564 6944 18570 6956
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 7708 6888 8800 6916
rect 7708 6876 7714 6888
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 12345 6919 12403 6925
rect 12345 6916 12357 6919
rect 10192 6888 12357 6916
rect 10192 6876 10198 6888
rect 12345 6885 12357 6888
rect 12391 6885 12403 6919
rect 12345 6879 12403 6885
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 15654 6916 15660 6928
rect 12492 6888 15660 6916
rect 12492 6876 12498 6888
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 16390 6876 16396 6928
rect 16448 6916 16454 6928
rect 16448 6888 23888 6916
rect 16448 6876 16454 6888
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 8904 6820 9413 6848
rect 8904 6808 8910 6820
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 10091 6820 16681 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 16669 6817 16681 6820
rect 16715 6848 16727 6851
rect 17402 6848 17408 6860
rect 16715 6820 17408 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 17552 6820 18644 6848
rect 17552 6808 17558 6820
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7800 6752 7941 6780
rect 7800 6740 7806 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 8754 6780 8760 6792
rect 8619 6752 8760 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9582 6780 9588 6792
rect 9543 6752 9588 6780
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6780 11483 6783
rect 11790 6780 11796 6792
rect 11471 6752 11796 6780
rect 11471 6749 11483 6752
rect 11425 6743 11483 6749
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 12618 6780 12624 6792
rect 12575 6752 12624 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6780 13047 6783
rect 13906 6780 13912 6792
rect 13035 6752 13912 6780
rect 13035 6749 13047 6752
rect 12989 6743 13047 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6780 14979 6783
rect 15194 6780 15200 6792
rect 14967 6752 15200 6780
rect 14967 6749 14979 6752
rect 14921 6743 14979 6749
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 15565 6783 15623 6789
rect 15565 6749 15577 6783
rect 15611 6749 15623 6783
rect 15565 6743 15623 6749
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16482 6780 16488 6792
rect 16255 6752 16488 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 8478 6712 8484 6724
rect 7760 6684 8484 6712
rect 7760 6653 7788 6684
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 8772 6712 8800 6740
rect 9490 6712 9496 6724
rect 8772 6684 9496 6712
rect 9490 6672 9496 6684
rect 9548 6672 9554 6724
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13081 6715 13139 6721
rect 13081 6712 13093 6715
rect 12952 6684 13093 6712
rect 12952 6672 12958 6684
rect 13081 6681 13093 6684
rect 13127 6681 13139 6715
rect 15580 6712 15608 6743
rect 13081 6675 13139 6681
rect 14752 6684 15608 6712
rect 16040 6712 16068 6743
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17773 6783 17831 6789
rect 17276 6752 17321 6780
rect 17276 6740 17282 6752
rect 17773 6749 17785 6783
rect 17819 6780 17831 6783
rect 18506 6780 18512 6792
rect 17819 6752 18512 6780
rect 17819 6749 17831 6752
rect 17773 6743 17831 6749
rect 16850 6712 16856 6724
rect 16040 6684 16856 6712
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6613 7803 6647
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 7745 6607 7803 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 14752 6653 14780 6684
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6613 14795 6647
rect 14737 6607 14795 6613
rect 15381 6647 15439 6653
rect 15381 6613 15393 6647
rect 15427 6644 15439 6647
rect 16574 6644 16580 6656
rect 15427 6616 16580 6644
rect 15427 6613 15439 6616
rect 15381 6607 15439 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17788 6644 17816 6743
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18616 6789 18644 6820
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 19334 6848 19340 6860
rect 18748 6820 19340 6848
rect 18748 6808 18754 6820
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6848 19579 6851
rect 20622 6848 20628 6860
rect 19567 6820 20628 6848
rect 19567 6817 19579 6820
rect 19521 6811 19579 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 21266 6848 21272 6860
rect 21227 6820 21272 6848
rect 21266 6808 21272 6820
rect 21324 6808 21330 6860
rect 22186 6848 22192 6860
rect 22147 6820 22192 6848
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 23290 6848 23296 6860
rect 22704 6820 23296 6848
rect 22704 6808 22710 6820
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 23750 6848 23756 6860
rect 23711 6820 23756 6848
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 18601 6783 18659 6789
rect 18601 6749 18613 6783
rect 18647 6749 18659 6783
rect 18601 6743 18659 6749
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19024 6752 19441 6780
rect 19024 6740 19030 6752
rect 19429 6749 19441 6752
rect 19475 6780 19487 6783
rect 20346 6780 20352 6792
rect 19475 6752 20352 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 20346 6740 20352 6752
rect 20404 6740 20410 6792
rect 17865 6715 17923 6721
rect 17865 6681 17877 6715
rect 17911 6712 17923 6715
rect 19978 6712 19984 6724
rect 17911 6684 19984 6712
rect 17911 6681 17923 6684
rect 17865 6675 17923 6681
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 20438 6672 20444 6724
rect 20496 6712 20502 6724
rect 20625 6715 20683 6721
rect 20625 6712 20637 6715
rect 20496 6684 20637 6712
rect 20496 6672 20502 6684
rect 20625 6681 20637 6684
rect 20671 6681 20683 6715
rect 20625 6675 20683 6681
rect 20717 6715 20775 6721
rect 20717 6681 20729 6715
rect 20763 6712 20775 6715
rect 20806 6712 20812 6724
rect 20763 6684 20812 6712
rect 20763 6681 20775 6684
rect 20717 6675 20775 6681
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 21821 6715 21879 6721
rect 21821 6681 21833 6715
rect 21867 6681 21879 6715
rect 21821 6675 21879 6681
rect 21913 6715 21971 6721
rect 21913 6681 21925 6715
rect 21959 6712 21971 6715
rect 22278 6712 22284 6724
rect 21959 6684 22284 6712
rect 21959 6681 21971 6684
rect 21913 6675 21971 6681
rect 17276 6616 17816 6644
rect 17276 6604 17282 6616
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 21358 6644 21364 6656
rect 18196 6616 21364 6644
rect 18196 6604 18202 6616
rect 21358 6604 21364 6616
rect 21416 6604 21422 6656
rect 21836 6644 21864 6675
rect 22278 6672 22284 6684
rect 22336 6672 22342 6724
rect 23106 6712 23112 6724
rect 23067 6684 23112 6712
rect 23106 6672 23112 6684
rect 23164 6672 23170 6724
rect 23201 6715 23259 6721
rect 23201 6681 23213 6715
rect 23247 6712 23259 6715
rect 23382 6712 23388 6724
rect 23247 6684 23388 6712
rect 23247 6681 23259 6684
rect 23201 6675 23259 6681
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 23860 6712 23888 6888
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 24780 6848 24900 6860
rect 27157 6851 27215 6857
rect 27157 6848 27169 6851
rect 24544 6832 27169 6848
rect 24544 6820 24808 6832
rect 24872 6820 27169 6832
rect 24544 6808 24550 6820
rect 27157 6817 27169 6820
rect 27203 6817 27215 6851
rect 27157 6811 27215 6817
rect 24578 6740 24584 6792
rect 24636 6780 24642 6792
rect 24857 6783 24915 6789
rect 24857 6780 24869 6783
rect 24636 6752 24869 6780
rect 24636 6740 24642 6752
rect 24857 6749 24869 6752
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 26234 6740 26240 6792
rect 26292 6740 26298 6792
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6780 27123 6783
rect 28353 6783 28411 6789
rect 27111 6752 28212 6780
rect 27111 6749 27123 6752
rect 27065 6743 27123 6749
rect 25133 6715 25191 6721
rect 25133 6712 25145 6715
rect 23860 6684 25145 6712
rect 25133 6681 25145 6684
rect 25179 6712 25191 6715
rect 25406 6712 25412 6724
rect 25179 6684 25412 6712
rect 25179 6681 25191 6684
rect 25133 6675 25191 6681
rect 25406 6672 25412 6684
rect 25464 6672 25470 6724
rect 27614 6712 27620 6724
rect 26436 6684 27620 6712
rect 26436 6644 26464 6684
rect 27614 6672 27620 6684
rect 27672 6672 27678 6724
rect 21836 6616 26464 6644
rect 26510 6604 26516 6656
rect 26568 6644 26574 6656
rect 28184 6653 28212 6752
rect 28353 6749 28365 6783
rect 28399 6780 28411 6783
rect 29914 6780 29920 6792
rect 28399 6752 29920 6780
rect 28399 6749 28411 6752
rect 28353 6743 28411 6749
rect 29914 6740 29920 6752
rect 29972 6740 29978 6792
rect 26605 6647 26663 6653
rect 26605 6644 26617 6647
rect 26568 6616 26617 6644
rect 26568 6604 26574 6616
rect 26605 6613 26617 6616
rect 26651 6613 26663 6647
rect 26605 6607 26663 6613
rect 28169 6647 28227 6653
rect 28169 6613 28181 6647
rect 28215 6613 28227 6647
rect 28169 6607 28227 6613
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7800 6412 8033 6440
rect 7800 6400 7806 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 11054 6440 11060 6452
rect 10459 6412 11060 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 14550 6440 14556 6452
rect 11900 6412 14556 6440
rect 5718 6372 5724 6384
rect 1596 6344 5724 6372
rect 1596 6313 1624 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 7469 6375 7527 6381
rect 7469 6341 7481 6375
rect 7515 6372 7527 6375
rect 8662 6372 8668 6384
rect 7515 6344 8668 6372
rect 7515 6341 7527 6344
rect 7469 6335 7527 6341
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 9824 6344 10364 6372
rect 9824 6332 9830 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 6822 6304 6828 6316
rect 4387 6276 6828 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 7650 6304 7656 6316
rect 7423 6276 7656 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 7650 6264 7656 6276
rect 7708 6304 7714 6316
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 7708 6276 8217 6304
rect 7708 6264 7714 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 9030 6304 9036 6316
rect 8991 6276 9036 6304
rect 8205 6267 8263 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9858 6304 9864 6316
rect 9819 6276 9864 6304
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10336 6313 10364 6344
rect 11900 6313 11928 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 15010 6440 15016 6452
rect 14792 6412 15016 6440
rect 14792 6400 14798 6412
rect 15010 6400 15016 6412
rect 15068 6440 15074 6452
rect 15381 6443 15439 6449
rect 15381 6440 15393 6443
rect 15068 6412 15393 6440
rect 15068 6400 15074 6412
rect 15381 6409 15393 6412
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 16209 6443 16267 6449
rect 16209 6409 16221 6443
rect 16255 6440 16267 6443
rect 16298 6440 16304 6452
rect 16255 6412 16304 6440
rect 16255 6409 16267 6412
rect 16209 6403 16267 6409
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 18966 6440 18972 6452
rect 17368 6412 18972 6440
rect 17368 6400 17374 6412
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 19150 6440 19156 6452
rect 19111 6412 19156 6440
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 20438 6440 20444 6452
rect 19392 6412 20444 6440
rect 19392 6400 19398 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 20809 6443 20867 6449
rect 20809 6409 20821 6443
rect 20855 6440 20867 6443
rect 27157 6443 27215 6449
rect 20855 6412 26004 6440
rect 20855 6409 20867 6412
rect 20809 6403 20867 6409
rect 12526 6372 12532 6384
rect 11992 6344 12532 6372
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11195 6276 11897 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 11992 6236 12020 6344
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 14366 6332 14372 6384
rect 14424 6372 14430 6384
rect 17497 6375 17555 6381
rect 17497 6372 17509 6375
rect 14424 6344 17509 6372
rect 14424 6332 14430 6344
rect 17497 6341 17509 6344
rect 17543 6341 17555 6375
rect 20257 6375 20315 6381
rect 20257 6372 20269 6375
rect 17497 6335 17555 6341
rect 18064 6344 20269 6372
rect 12710 6304 12716 6316
rect 12671 6276 12716 6304
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 13630 6304 13636 6316
rect 13543 6276 13636 6304
rect 13630 6264 13636 6276
rect 13688 6304 13694 6316
rect 13688 6276 13952 6304
rect 13688 6264 13694 6276
rect 12526 6236 12532 6248
rect 9171 6208 12020 6236
rect 12487 6208 12532 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 13170 6236 13176 6248
rect 13131 6208 13176 6236
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13780 6208 13829 6236
rect 13780 6196 13786 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13924 6236 13952 6276
rect 14182 6264 14188 6316
rect 14240 6304 14246 6316
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14240 6276 14933 6304
rect 14240 6264 14246 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 17126 6304 17132 6316
rect 16163 6276 17132 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 14734 6236 14740 6248
rect 13924 6208 14596 6236
rect 14695 6208 14740 6236
rect 13817 6199 13875 6205
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 9766 6128 9772 6180
rect 9824 6168 9830 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 9824 6140 10977 6168
rect 9824 6128 9830 6140
rect 10965 6137 10977 6140
rect 11011 6137 11023 6171
rect 10965 6131 11023 6137
rect 13078 6128 13084 6180
rect 13136 6168 13142 6180
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 13136 6140 14013 6168
rect 13136 6128 13142 6140
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14568 6168 14596 6208
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 17402 6236 17408 6248
rect 17363 6208 17408 6236
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 18064 6236 18092 6344
rect 20257 6341 20269 6344
rect 20303 6341 20315 6375
rect 20257 6335 20315 6341
rect 20346 6332 20352 6384
rect 20404 6372 20410 6384
rect 22097 6375 22155 6381
rect 22097 6372 22109 6375
rect 20404 6344 20760 6372
rect 20404 6332 20410 6344
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 19797 6307 19855 6313
rect 19300 6276 19748 6304
rect 19300 6264 19306 6276
rect 17512 6208 18092 6236
rect 17512 6168 17540 6208
rect 18230 6196 18236 6248
rect 18288 6236 18294 6248
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 18288 6208 18521 6236
rect 18288 6196 18294 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 18690 6236 18696 6248
rect 18651 6208 18696 6236
rect 18509 6199 18567 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 19610 6236 19616 6248
rect 19571 6208 19616 6236
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 19720 6236 19748 6276
rect 19797 6273 19809 6307
rect 19843 6304 19855 6307
rect 20622 6304 20628 6316
rect 19843 6276 20628 6304
rect 19843 6273 19855 6276
rect 19797 6267 19855 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 20732 6313 20760 6344
rect 20824 6344 22109 6372
rect 20824 6316 20852 6344
rect 22097 6341 22109 6344
rect 22143 6341 22155 6375
rect 22097 6335 22155 6341
rect 22833 6375 22891 6381
rect 22833 6341 22845 6375
rect 22879 6372 22891 6375
rect 23198 6372 23204 6384
rect 22879 6344 23204 6372
rect 22879 6341 22891 6344
rect 22833 6335 22891 6341
rect 23198 6332 23204 6344
rect 23256 6332 23262 6384
rect 23385 6375 23443 6381
rect 23385 6341 23397 6375
rect 23431 6372 23443 6375
rect 23658 6372 23664 6384
rect 23431 6344 23664 6372
rect 23431 6341 23443 6344
rect 23385 6335 23443 6341
rect 23658 6332 23664 6344
rect 23716 6372 23722 6384
rect 24854 6372 24860 6384
rect 23716 6344 24860 6372
rect 23716 6332 23722 6344
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 25130 6332 25136 6384
rect 25188 6372 25194 6384
rect 25409 6375 25467 6381
rect 25409 6372 25421 6375
rect 25188 6344 25421 6372
rect 25188 6332 25194 6344
rect 25409 6341 25421 6344
rect 25455 6341 25467 6375
rect 25409 6335 25467 6341
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 20806 6264 20812 6316
rect 20864 6264 20870 6316
rect 21542 6264 21548 6316
rect 21600 6304 21606 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21600 6276 22017 6304
rect 21600 6264 21606 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 23474 6264 23480 6316
rect 23532 6304 23538 6316
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 23532 6276 24133 6304
rect 23532 6264 23538 6276
rect 24121 6273 24133 6276
rect 24167 6304 24179 6307
rect 24762 6304 24768 6316
rect 24167 6276 24768 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 24762 6264 24768 6276
rect 24820 6264 24826 6316
rect 19720 6208 20668 6236
rect 14568 6140 17540 6168
rect 17957 6171 18015 6177
rect 14001 6131 14059 6137
rect 17957 6137 17969 6171
rect 18003 6168 18015 6171
rect 18138 6168 18144 6180
rect 18003 6140 18144 6168
rect 18003 6137 18015 6140
rect 17957 6131 18015 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 18874 6128 18880 6180
rect 18932 6168 18938 6180
rect 20640 6168 20668 6208
rect 21358 6196 21364 6248
rect 21416 6236 21422 6248
rect 22554 6236 22560 6248
rect 21416 6208 22560 6236
rect 21416 6196 21422 6208
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 22741 6239 22799 6245
rect 22741 6205 22753 6239
rect 22787 6236 22799 6239
rect 22922 6236 22928 6248
rect 22787 6208 22928 6236
rect 22787 6205 22799 6208
rect 22741 6199 22799 6205
rect 22922 6196 22928 6208
rect 22980 6196 22986 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23124 6208 24225 6236
rect 23124 6168 23152 6208
rect 24213 6205 24225 6208
rect 24259 6205 24271 6239
rect 24213 6199 24271 6205
rect 24670 6196 24676 6248
rect 24728 6236 24734 6248
rect 25317 6239 25375 6245
rect 25317 6236 25329 6239
rect 24728 6208 25329 6236
rect 24728 6196 24734 6208
rect 25317 6205 25329 6208
rect 25363 6205 25375 6239
rect 25682 6236 25688 6248
rect 25643 6208 25688 6236
rect 25317 6199 25375 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 25976 6236 26004 6412
rect 27157 6409 27169 6443
rect 27203 6409 27215 6443
rect 27157 6403 27215 6409
rect 27172 6372 27200 6403
rect 27172 6344 28120 6372
rect 26602 6304 26608 6316
rect 26563 6276 26608 6304
rect 26602 6264 26608 6276
rect 26660 6264 26666 6316
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 28092 6313 28120 6344
rect 27341 6307 27399 6313
rect 27341 6304 27353 6307
rect 27304 6276 27353 6304
rect 27304 6264 27310 6276
rect 27341 6273 27353 6276
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 27798 6236 27804 6248
rect 25976 6208 27804 6236
rect 27798 6196 27804 6208
rect 27856 6196 27862 6248
rect 18932 6140 20392 6168
rect 20640 6140 23152 6168
rect 25700 6168 25728 6196
rect 26234 6168 26240 6180
rect 25700 6140 26240 6168
rect 18932 6128 18938 6140
rect 4154 6100 4160 6112
rect 4115 6072 4160 6100
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 11882 6100 11888 6112
rect 9723 6072 11888 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 15746 6100 15752 6112
rect 12023 6072 15752 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 20070 6100 20076 6112
rect 16908 6072 20076 6100
rect 16908 6060 16914 6072
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20364 6100 20392 6140
rect 26234 6128 26240 6140
rect 26292 6128 26298 6180
rect 28258 6168 28264 6180
rect 28219 6140 28264 6168
rect 28258 6128 28264 6140
rect 28316 6128 28322 6180
rect 23658 6100 23664 6112
rect 20364 6072 23664 6100
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 26421 6103 26479 6109
rect 26421 6069 26433 6103
rect 26467 6100 26479 6103
rect 28074 6100 28080 6112
rect 26467 6072 28080 6100
rect 26467 6069 26479 6072
rect 26421 6063 26479 6069
rect 28074 6060 28080 6072
rect 28132 6060 28138 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 5261 5899 5319 5905
rect 5261 5865 5273 5899
rect 5307 5896 5319 5899
rect 8846 5896 8852 5908
rect 5307 5868 8852 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 10689 5899 10747 5905
rect 10689 5865 10701 5899
rect 10735 5896 10747 5899
rect 10962 5896 10968 5908
rect 10735 5868 10968 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 14366 5896 14372 5908
rect 14327 5868 14372 5896
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 19058 5896 19064 5908
rect 14516 5868 19064 5896
rect 14516 5856 14522 5868
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5828 10011 5831
rect 12342 5828 12348 5840
rect 9999 5800 12348 5828
rect 9999 5797 10011 5800
rect 9953 5791 10011 5797
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 13078 5828 13084 5840
rect 13039 5800 13084 5828
rect 13078 5788 13084 5800
rect 13136 5788 13142 5840
rect 13170 5788 13176 5840
rect 13228 5828 13234 5840
rect 15565 5831 15623 5837
rect 13228 5800 15148 5828
rect 13228 5788 13234 5800
rect 6546 5760 6552 5772
rect 4724 5732 6552 5760
rect 4724 5701 4752 5732
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 10502 5760 10508 5772
rect 9447 5732 10508 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 10502 5720 10508 5732
rect 10560 5760 10566 5772
rect 11241 5763 11299 5769
rect 11241 5760 11253 5763
rect 10560 5732 11253 5760
rect 10560 5720 10566 5732
rect 11241 5729 11253 5732
rect 11287 5760 11299 5763
rect 12526 5760 12532 5772
rect 11287 5732 12532 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 15010 5760 15016 5772
rect 14971 5732 15016 5760
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15120 5760 15148 5800
rect 15565 5797 15577 5831
rect 15611 5828 15623 5831
rect 18874 5828 18880 5840
rect 15611 5800 18880 5828
rect 15611 5797 15623 5800
rect 15565 5791 15623 5797
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 18984 5828 19012 5868
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 23017 5899 23075 5905
rect 23017 5896 23029 5899
rect 19668 5868 23029 5896
rect 19668 5856 19674 5868
rect 23017 5865 23029 5868
rect 23063 5865 23075 5899
rect 23017 5859 23075 5865
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 24946 5896 24952 5908
rect 23164 5868 24952 5896
rect 23164 5856 23170 5868
rect 24946 5856 24952 5868
rect 25004 5856 25010 5908
rect 25038 5856 25044 5908
rect 25096 5896 25102 5908
rect 25317 5899 25375 5905
rect 25317 5896 25329 5899
rect 25096 5868 25329 5896
rect 25096 5856 25102 5868
rect 25317 5865 25329 5868
rect 25363 5865 25375 5899
rect 26602 5896 26608 5908
rect 26563 5868 26608 5896
rect 25317 5859 25375 5865
rect 26602 5856 26608 5868
rect 26660 5856 26666 5908
rect 27246 5896 27252 5908
rect 27207 5868 27252 5896
rect 27246 5856 27252 5868
rect 27304 5856 27310 5908
rect 19886 5828 19892 5840
rect 18984 5800 19892 5828
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 20346 5788 20352 5840
rect 20404 5828 20410 5840
rect 20806 5828 20812 5840
rect 20404 5800 20812 5828
rect 20404 5788 20410 5800
rect 20806 5788 20812 5800
rect 20864 5788 20870 5840
rect 21174 5788 21180 5840
rect 21232 5828 21238 5840
rect 22373 5831 22431 5837
rect 22373 5828 22385 5831
rect 21232 5800 22385 5828
rect 21232 5788 21238 5800
rect 22373 5797 22385 5800
rect 22419 5797 22431 5831
rect 24670 5828 24676 5840
rect 24631 5800 24676 5828
rect 22373 5791 22431 5797
rect 24670 5788 24676 5800
rect 24728 5788 24734 5840
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 15120 5732 17509 5760
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 22554 5720 22560 5772
rect 22612 5760 22618 5772
rect 22612 5732 27844 5760
rect 22612 5720 22618 5732
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 9306 5692 9312 5704
rect 9267 5664 9312 5692
rect 7837 5655 7895 5661
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 5184 5624 5212 5655
rect 3936 5596 5212 5624
rect 7852 5624 7880 5655
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9548 5664 10149 5692
rect 9548 5652 9554 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 11146 5692 11152 5704
rect 10643 5664 11152 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11422 5692 11428 5704
rect 11383 5664 11428 5692
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 12158 5692 12164 5704
rect 11931 5664 12164 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 12158 5652 12164 5664
rect 12216 5692 12222 5704
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12216 5664 12725 5692
rect 12216 5652 12222 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12894 5692 12900 5704
rect 12855 5664 12900 5692
rect 12713 5655 12771 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13872 5664 14289 5692
rect 13872 5652 13878 5664
rect 14277 5661 14289 5664
rect 14323 5692 14335 5695
rect 14458 5692 14464 5704
rect 14323 5664 14464 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 16390 5692 16396 5704
rect 16351 5664 16396 5692
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 18693 5695 18751 5701
rect 16540 5664 16585 5692
rect 16540 5652 16546 5664
rect 18693 5661 18705 5695
rect 18739 5692 18751 5695
rect 19518 5692 19524 5704
rect 18739 5664 19524 5692
rect 18739 5661 18751 5664
rect 18693 5655 18751 5661
rect 19518 5652 19524 5664
rect 19576 5692 19582 5704
rect 19981 5695 20039 5701
rect 19576 5664 19932 5692
rect 19576 5652 19582 5664
rect 14642 5624 14648 5636
rect 7852 5596 14648 5624
rect 3936 5584 3942 5596
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 15105 5627 15163 5633
rect 15105 5593 15117 5627
rect 15151 5593 15163 5627
rect 15105 5587 15163 5593
rect 17589 5627 17647 5633
rect 17589 5593 17601 5627
rect 17635 5593 17647 5627
rect 17589 5587 17647 5593
rect 18141 5627 18199 5633
rect 18141 5593 18153 5627
rect 18187 5624 18199 5627
rect 19904 5624 19932 5664
rect 19981 5661 19993 5695
rect 20027 5692 20039 5695
rect 20070 5692 20076 5704
rect 20027 5664 20076 5692
rect 20027 5661 20039 5664
rect 19981 5655 20039 5661
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20346 5692 20352 5704
rect 20211 5664 20352 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 20438 5652 20444 5704
rect 20496 5692 20502 5704
rect 20625 5695 20683 5701
rect 20625 5692 20637 5695
rect 20496 5664 20637 5692
rect 20496 5652 20502 5664
rect 20625 5661 20637 5664
rect 20671 5661 20683 5695
rect 22278 5692 22284 5704
rect 22239 5664 22284 5692
rect 20625 5655 20683 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 22925 5695 22983 5701
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 23106 5692 23112 5704
rect 22971 5664 23112 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 23290 5652 23296 5704
rect 23348 5692 23354 5704
rect 23569 5695 23627 5701
rect 23569 5692 23581 5695
rect 23348 5664 23581 5692
rect 23348 5652 23354 5664
rect 23569 5661 23581 5664
rect 23615 5661 23627 5695
rect 24578 5692 24584 5704
rect 24539 5664 24584 5692
rect 23569 5655 23627 5661
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25225 5695 25283 5701
rect 25225 5692 25237 5695
rect 24820 5664 25237 5692
rect 24820 5652 24826 5664
rect 25225 5661 25237 5664
rect 25271 5661 25283 5695
rect 26050 5692 26056 5704
rect 26011 5664 26056 5692
rect 25225 5655 25283 5661
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 26513 5695 26571 5701
rect 26513 5661 26525 5695
rect 26559 5661 26571 5695
rect 27154 5692 27160 5704
rect 27115 5664 27160 5692
rect 26513 5655 26571 5661
rect 20898 5624 20904 5636
rect 18187 5596 19840 5624
rect 19904 5596 20904 5624
rect 18187 5593 18199 5596
rect 18141 5587 18199 5593
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 4304 5528 4537 5556
rect 4304 5516 4310 5528
rect 4525 5525 4537 5528
rect 4571 5525 4583 5559
rect 4525 5519 4583 5525
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 6972 5528 7941 5556
rect 6972 5516 6978 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 7929 5519 7987 5525
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 15113 5556 15141 5587
rect 14332 5528 15141 5556
rect 17604 5556 17632 5587
rect 18785 5559 18843 5565
rect 18785 5556 18797 5559
rect 17604 5528 18797 5556
rect 14332 5516 14338 5528
rect 18785 5525 18797 5528
rect 18831 5525 18843 5559
rect 19812 5556 19840 5596
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 22738 5584 22744 5636
rect 22796 5624 22802 5636
rect 26528 5624 26556 5655
rect 27154 5652 27160 5664
rect 27212 5652 27218 5704
rect 27816 5701 27844 5732
rect 27801 5695 27859 5701
rect 27801 5661 27813 5695
rect 27847 5661 27859 5695
rect 27801 5655 27859 5661
rect 22796 5596 26556 5624
rect 22796 5584 22802 5596
rect 21174 5556 21180 5568
rect 19812 5528 21180 5556
rect 18785 5519 18843 5525
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 23658 5556 23664 5568
rect 23619 5528 23664 5556
rect 23658 5516 23664 5528
rect 23716 5516 23722 5568
rect 25869 5559 25927 5565
rect 25869 5525 25881 5559
rect 25915 5556 25927 5559
rect 26050 5556 26056 5568
rect 25915 5528 26056 5556
rect 25915 5525 25927 5528
rect 25869 5519 25927 5525
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 27890 5556 27896 5568
rect 27851 5528 27896 5556
rect 27890 5516 27896 5528
rect 27948 5516 27954 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 9309 5355 9367 5361
rect 9309 5321 9321 5355
rect 9355 5352 9367 5355
rect 9858 5352 9864 5364
rect 9355 5324 9864 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 11422 5352 11428 5364
rect 10091 5324 11428 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 12345 5355 12403 5361
rect 12345 5321 12357 5355
rect 12391 5352 12403 5355
rect 13722 5352 13728 5364
rect 12391 5324 13728 5352
rect 12391 5321 12403 5324
rect 12345 5315 12403 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 14185 5355 14243 5361
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 14274 5352 14280 5364
rect 14231 5324 14280 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14792 5324 14841 5352
rect 14792 5312 14798 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 15473 5355 15531 5361
rect 15473 5321 15485 5355
rect 15519 5352 15531 5355
rect 17494 5352 17500 5364
rect 15519 5324 17500 5352
rect 15519 5321 15531 5324
rect 15473 5315 15531 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 21082 5352 21088 5364
rect 17911 5324 21088 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 21266 5312 21272 5364
rect 21324 5352 21330 5364
rect 21324 5324 24992 5352
rect 21324 5312 21330 5324
rect 6454 5284 6460 5296
rect 1596 5256 6460 5284
rect 1596 5225 1624 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 14550 5284 14556 5296
rect 9968 5256 14556 5284
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 4154 5216 4160 5228
rect 4115 5188 4160 5216
rect 1581 5179 1639 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 8864 5080 8892 5179
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9968 5225 9996 5256
rect 14550 5244 14556 5256
rect 14608 5244 14614 5296
rect 16022 5244 16028 5296
rect 16080 5284 16086 5296
rect 16209 5287 16267 5293
rect 16209 5284 16221 5287
rect 16080 5256 16221 5284
rect 16080 5244 16086 5256
rect 16209 5253 16221 5256
rect 16255 5253 16267 5287
rect 16209 5247 16267 5253
rect 17221 5287 17279 5293
rect 17221 5253 17233 5287
rect 17267 5284 17279 5287
rect 18046 5284 18052 5296
rect 17267 5256 18052 5284
rect 17267 5253 17279 5256
rect 17221 5247 17279 5253
rect 18046 5244 18052 5256
rect 18104 5244 18110 5296
rect 19334 5284 19340 5296
rect 19295 5256 19340 5284
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 20901 5287 20959 5293
rect 20901 5253 20913 5287
rect 20947 5284 20959 5287
rect 23014 5284 23020 5296
rect 20947 5256 23020 5284
rect 20947 5253 20959 5256
rect 20901 5247 20959 5253
rect 23014 5244 23020 5256
rect 23072 5244 23078 5296
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 8996 5188 9505 5216
rect 8996 5176 9002 5188
rect 9493 5185 9505 5188
rect 9539 5216 9551 5219
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9539 5188 9965 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 11195 5188 12265 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12268 5148 12296 5179
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12400 5188 13093 5216
rect 12400 5176 12406 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13722 5216 13728 5228
rect 13683 5188 13728 5216
rect 13081 5179 13139 5185
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 14332 5188 14381 5216
rect 14332 5176 14338 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15620 5188 15669 5216
rect 15620 5176 15626 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16850 5216 16856 5228
rect 16163 5188 16856 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17368 5188 17785 5216
rect 17368 5176 17374 5188
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5216 18567 5219
rect 18966 5216 18972 5228
rect 18555 5188 18972 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 22554 5216 22560 5228
rect 22515 5188 22560 5216
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 23658 5176 23664 5228
rect 23716 5216 23722 5228
rect 24964 5225 24992 5324
rect 26050 5284 26056 5296
rect 26011 5256 26056 5284
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 26234 5244 26240 5296
rect 26292 5284 26298 5296
rect 26605 5287 26663 5293
rect 26605 5284 26617 5287
rect 26292 5256 26617 5284
rect 26292 5244 26298 5256
rect 26605 5253 26617 5256
rect 26651 5253 26663 5287
rect 26605 5247 26663 5253
rect 24029 5219 24087 5225
rect 24029 5216 24041 5219
rect 23716 5188 24041 5216
rect 23716 5176 23722 5188
rect 24029 5185 24041 5188
rect 24075 5185 24087 5219
rect 24029 5179 24087 5185
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5185 25007 5219
rect 28074 5216 28080 5228
rect 28035 5188 28080 5216
rect 24949 5179 25007 5185
rect 28074 5176 28080 5188
rect 28132 5176 28138 5228
rect 15378 5148 15384 5160
rect 12268 5120 15384 5148
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 17144 5148 17172 5176
rect 17862 5148 17868 5160
rect 17144 5120 17868 5148
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5117 19303 5151
rect 19245 5111 19303 5117
rect 11974 5080 11980 5092
rect 8864 5052 11980 5080
rect 11974 5040 11980 5052
rect 12032 5040 12038 5092
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 12986 5080 12992 5092
rect 12943 5052 12992 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 19150 5040 19156 5092
rect 19208 5080 19214 5092
rect 19260 5080 19288 5111
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 19521 5151 19579 5157
rect 19521 5148 19533 5151
rect 19484 5120 19533 5148
rect 19484 5108 19490 5120
rect 19521 5117 19533 5120
rect 19567 5117 19579 5151
rect 20806 5148 20812 5160
rect 20767 5120 20812 5148
rect 19521 5111 19579 5117
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5117 21143 5151
rect 22738 5148 22744 5160
rect 22699 5120 22744 5148
rect 21085 5111 21143 5117
rect 19208 5052 19288 5080
rect 19208 5040 19214 5052
rect 20070 5040 20076 5092
rect 20128 5080 20134 5092
rect 20128 5052 20668 5080
rect 20128 5040 20134 5052
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 8662 5012 8668 5024
rect 8623 4984 8668 5012
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 12066 5012 12072 5024
rect 11011 4984 12072 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 13538 5012 13544 5024
rect 13499 4984 13544 5012
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14642 5012 14648 5024
rect 14056 4984 14648 5012
rect 14056 4972 14062 4984
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 18601 5015 18659 5021
rect 18601 4981 18613 5015
rect 18647 5012 18659 5015
rect 20346 5012 20352 5024
rect 18647 4984 20352 5012
rect 18647 4981 18659 4984
rect 18601 4975 18659 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20640 5012 20668 5052
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 21100 5080 21128 5111
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 23845 5151 23903 5157
rect 23845 5117 23857 5151
rect 23891 5148 23903 5151
rect 24670 5148 24676 5160
rect 23891 5120 24676 5148
rect 23891 5117 23903 5120
rect 23845 5111 23903 5117
rect 24670 5108 24676 5120
rect 24728 5108 24734 5160
rect 25961 5151 26019 5157
rect 25961 5117 25973 5151
rect 26007 5148 26019 5151
rect 27614 5148 27620 5160
rect 26007 5120 27620 5148
rect 26007 5117 26019 5120
rect 25961 5111 26019 5117
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 22922 5080 22928 5092
rect 20772 5052 21128 5080
rect 22883 5052 22928 5080
rect 20772 5040 20778 5052
rect 22922 5040 22928 5052
rect 22980 5080 22986 5092
rect 24213 5083 24271 5089
rect 24213 5080 24225 5083
rect 22980 5052 24225 5080
rect 22980 5040 22986 5052
rect 24213 5049 24225 5052
rect 24259 5049 24271 5083
rect 24213 5043 24271 5049
rect 22370 5012 22376 5024
rect 20640 4984 22376 5012
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 25041 5015 25099 5021
rect 25041 4981 25053 5015
rect 25087 5012 25099 5015
rect 25866 5012 25872 5024
rect 25087 4984 25872 5012
rect 25087 4981 25099 4984
rect 25041 4975 25099 4981
rect 25866 4972 25872 4984
rect 25924 4972 25930 5024
rect 28258 5012 28264 5024
rect 28219 4984 28264 5012
rect 28258 4972 28264 4984
rect 28316 4972 28322 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9582 4808 9588 4820
rect 9171 4780 9588 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 12158 4808 12164 4820
rect 12119 4780 12164 4808
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13722 4808 13728 4820
rect 12943 4780 13728 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14274 4808 14280 4820
rect 14235 4780 14280 4808
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 17678 4768 17684 4820
rect 17736 4768 17742 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 20806 4808 20812 4820
rect 20763 4780 20812 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 20806 4768 20812 4780
rect 20864 4768 20870 4820
rect 20990 4768 20996 4820
rect 21048 4808 21054 4820
rect 21361 4811 21419 4817
rect 21361 4808 21373 4811
rect 21048 4780 21373 4808
rect 21048 4768 21054 4780
rect 21361 4777 21373 4780
rect 21407 4777 21419 4811
rect 22370 4808 22376 4820
rect 22331 4780 22376 4808
rect 21361 4771 21419 4777
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 23014 4808 23020 4820
rect 22975 4780 23020 4808
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 23661 4811 23719 4817
rect 23661 4808 23673 4811
rect 23256 4780 23673 4808
rect 23256 4768 23262 4780
rect 23661 4777 23673 4780
rect 23707 4777 23719 4811
rect 23661 4771 23719 4777
rect 25225 4811 25283 4817
rect 25225 4777 25237 4811
rect 25271 4808 25283 4811
rect 26234 4808 26240 4820
rect 25271 4780 26240 4808
rect 25271 4777 25283 4780
rect 25225 4771 25283 4777
rect 26234 4768 26240 4780
rect 26292 4808 26298 4820
rect 27154 4808 27160 4820
rect 26292 4780 27160 4808
rect 26292 4768 26298 4780
rect 27154 4768 27160 4780
rect 27212 4768 27218 4820
rect 27614 4808 27620 4820
rect 27575 4780 27620 4808
rect 27614 4768 27620 4780
rect 27672 4768 27678 4820
rect 13541 4743 13599 4749
rect 13541 4709 13553 4743
rect 13587 4740 13599 4743
rect 14182 4740 14188 4752
rect 13587 4712 14188 4740
rect 13587 4709 13599 4712
rect 13541 4703 13599 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 14734 4700 14740 4752
rect 14792 4740 14798 4752
rect 17589 4743 17647 4749
rect 17589 4740 17601 4743
rect 14792 4712 17601 4740
rect 14792 4700 14798 4712
rect 17589 4709 17601 4712
rect 17635 4709 17647 4743
rect 17696 4740 17724 4768
rect 17696 4712 19472 4740
rect 17589 4703 17647 4709
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 9732 4644 11805 4672
rect 9732 4632 9738 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 14476 4644 16988 4672
rect 14476 4616 14504 4644
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6914 4604 6920 4616
rect 6227 4576 6920 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 8662 4564 8668 4616
rect 8720 4604 8726 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8720 4576 9321 4604
rect 8720 4564 8726 4576
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11011 4576 11621 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 13044 4576 13093 4604
rect 13044 4564 13050 4576
rect 13081 4573 13093 4576
rect 13127 4573 13139 4607
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 13081 4567 13139 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14458 4604 14464 4616
rect 14371 4576 14464 4604
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 15197 4607 15255 4613
rect 15197 4604 15209 4607
rect 14700 4576 15209 4604
rect 14700 4564 14706 4576
rect 15197 4573 15209 4576
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 15289 4539 15347 4545
rect 15289 4536 15301 4539
rect 11112 4508 15301 4536
rect 11112 4496 11118 4508
rect 15289 4505 15301 4508
rect 15335 4505 15347 4539
rect 15289 4499 15347 4505
rect 5994 4468 6000 4480
rect 5955 4440 6000 4468
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 10321 4471 10379 4477
rect 10321 4437 10333 4471
rect 10367 4468 10379 4471
rect 11698 4468 11704 4480
rect 10367 4440 11704 4468
rect 10367 4437 10379 4440
rect 10321 4431 10379 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15841 4471 15899 4477
rect 15841 4468 15853 4471
rect 15252 4440 15853 4468
rect 15252 4428 15258 4440
rect 15841 4437 15853 4440
rect 15887 4437 15899 4471
rect 16960 4468 16988 4644
rect 18230 4632 18236 4684
rect 18288 4672 18294 4684
rect 19444 4681 19472 4712
rect 19702 4700 19708 4752
rect 19760 4740 19766 4752
rect 19797 4743 19855 4749
rect 19797 4740 19809 4743
rect 19760 4712 19809 4740
rect 19760 4700 19766 4712
rect 19797 4709 19809 4712
rect 19843 4709 19855 4743
rect 19797 4703 19855 4709
rect 20346 4700 20352 4752
rect 20404 4740 20410 4752
rect 22830 4740 22836 4752
rect 20404 4712 22836 4740
rect 20404 4700 20410 4712
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 24946 4700 24952 4752
rect 25004 4740 25010 4752
rect 28261 4743 28319 4749
rect 28261 4740 28273 4743
rect 25004 4712 28273 4740
rect 25004 4700 25010 4712
rect 28261 4709 28273 4712
rect 28307 4709 28319 4743
rect 28261 4703 28319 4709
rect 18509 4675 18567 4681
rect 18509 4672 18521 4675
rect 18288 4644 18521 4672
rect 18288 4632 18294 4644
rect 18509 4641 18521 4644
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 20530 4672 20536 4684
rect 19475 4644 20536 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 20530 4632 20536 4644
rect 20588 4632 20594 4684
rect 26786 4672 26792 4684
rect 22940 4644 26792 4672
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 18138 4604 18144 4616
rect 17451 4576 18144 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 17236 4536 17264 4567
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 19610 4604 19616 4616
rect 19571 4576 19616 4604
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 20806 4604 20812 4616
rect 20671 4576 20812 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 21269 4607 21327 4613
rect 21269 4573 21281 4607
rect 21315 4573 21327 4607
rect 22278 4604 22284 4616
rect 22239 4576 22284 4604
rect 21269 4567 21327 4573
rect 19242 4536 19248 4548
rect 17236 4508 19248 4536
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 19978 4496 19984 4548
rect 20036 4536 20042 4548
rect 21284 4536 21312 4567
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 22940 4613 22968 4644
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4573 22983 4607
rect 22925 4567 22983 4573
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 23842 4604 23848 4616
rect 23615 4576 23848 4604
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 22186 4536 22192 4548
rect 20036 4508 22192 4536
rect 20036 4496 20042 4508
rect 22186 4496 22192 4508
rect 22244 4496 22250 4548
rect 23584 4468 23612 4567
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 23934 4564 23940 4616
rect 23992 4604 23998 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 23992 4576 24593 4604
rect 23992 4564 23998 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4604 24823 4607
rect 25130 4604 25136 4616
rect 24811 4576 25136 4604
rect 24811 4573 24823 4576
rect 24765 4567 24823 4573
rect 25130 4564 25136 4576
rect 25188 4564 25194 4616
rect 25866 4604 25872 4616
rect 25827 4576 25872 4604
rect 25866 4564 25872 4576
rect 25924 4564 25930 4616
rect 27522 4604 27528 4616
rect 27483 4576 27528 4604
rect 27522 4564 27528 4576
rect 27580 4564 27586 4616
rect 28169 4607 28227 4613
rect 28169 4573 28181 4607
rect 28215 4573 28227 4607
rect 28169 4567 28227 4573
rect 27246 4496 27252 4548
rect 27304 4536 27310 4548
rect 28184 4536 28212 4567
rect 27304 4508 28212 4536
rect 27304 4496 27310 4508
rect 16960 4440 23612 4468
rect 25685 4471 25743 4477
rect 15841 4431 15899 4437
rect 25685 4437 25697 4471
rect 25731 4468 25743 4471
rect 28074 4468 28080 4480
rect 25731 4440 28080 4468
rect 25731 4437 25743 4440
rect 25685 4431 25743 4437
rect 28074 4428 28080 4440
rect 28132 4428 28138 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 17862 4224 17868 4276
rect 17920 4264 17926 4276
rect 22189 4267 22247 4273
rect 17920 4236 19334 4264
rect 17920 4224 17926 4236
rect 13538 4196 13544 4208
rect 13499 4168 13544 4196
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 17954 4196 17960 4208
rect 17788 4168 17960 4196
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 7432 4100 7573 4128
rect 7432 4088 7438 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8938 4128 8944 4140
rect 8435 4100 8944 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 11054 4128 11060 4140
rect 10551 4100 11060 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 9048 4060 9076 4091
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11238 4128 11244 4140
rect 11195 4100 11244 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11698 4128 11704 4140
rect 11659 4100 11704 4128
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 14182 4128 14188 4140
rect 14139 4100 14188 4128
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4128 14795 4131
rect 14826 4128 14832 4140
rect 14783 4100 14832 4128
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 17037 4131 17095 4137
rect 15519 4100 16988 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 11882 4060 11888 4072
rect 8220 4032 9076 4060
rect 11843 4032 11888 4060
rect 8220 4001 8248 4032
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 14642 4060 14648 4072
rect 13495 4032 14648 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15620 4032 15669 4060
rect 15620 4020 15626 4032
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3961 8263 3995
rect 8205 3955 8263 3961
rect 8849 3995 8907 4001
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 9674 3992 9680 4004
rect 8895 3964 9680 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 10321 3995 10379 4001
rect 10321 3961 10333 3995
rect 10367 3992 10379 3995
rect 12250 3992 12256 4004
rect 10367 3964 12256 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 12250 3952 12256 3964
rect 12308 3952 12314 4004
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 12406 3964 15853 3992
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 7653 3927 7711 3933
rect 7653 3924 7665 3927
rect 5776 3896 7665 3924
rect 5776 3884 5782 3896
rect 7653 3893 7665 3896
rect 7699 3893 7711 3927
rect 7653 3887 7711 3893
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11974 3924 11980 3936
rect 11011 3896 11980 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 12158 3924 12164 3936
rect 12119 3896 12164 3924
rect 12158 3884 12164 3896
rect 12216 3924 12222 3936
rect 12406 3924 12434 3964
rect 15841 3961 15853 3964
rect 15887 3961 15899 3995
rect 16960 3992 16988 4100
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17788 4128 17816 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 17083 4100 17816 4128
rect 17865 4131 17923 4137
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18046 4128 18052 4140
rect 17911 4100 18052 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4097 18567 4131
rect 19306 4128 19334 4236
rect 22189 4233 22201 4267
rect 22235 4264 22247 4267
rect 22738 4264 22744 4276
rect 22235 4236 22744 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 23934 4264 23940 4276
rect 23895 4236 23940 4264
rect 23934 4224 23940 4236
rect 23992 4224 23998 4276
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 27080 4168 27292 4196
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19306 4100 19441 4128
rect 18509 4091 18567 4097
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 19521 4131 19579 4137
rect 19521 4097 19533 4131
rect 19567 4128 19579 4131
rect 19794 4128 19800 4140
rect 19567 4100 19800 4128
rect 19567 4097 19579 4100
rect 19521 4091 19579 4097
rect 18524 4060 18552 4091
rect 19794 4088 19800 4100
rect 19852 4088 19858 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 17696 4032 18552 4060
rect 20088 4060 20116 4091
rect 20162 4088 20168 4140
rect 20220 4128 20226 4140
rect 20898 4128 20904 4140
rect 20220 4100 20265 4128
rect 20859 4100 20904 4128
rect 20220 4088 20226 4100
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 22370 4128 22376 4140
rect 22331 4100 22376 4128
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 23293 4131 23351 4137
rect 23293 4097 23305 4131
rect 23339 4097 23351 4131
rect 23293 4091 23351 4097
rect 22646 4060 22652 4072
rect 20088 4032 22652 4060
rect 17696 4001 17724 4032
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 17681 3995 17739 4001
rect 16960 3964 17632 3992
rect 15841 3955 15899 3961
rect 14550 3924 14556 3936
rect 12216 3896 12434 3924
rect 14511 3896 14556 3924
rect 12216 3884 12222 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17129 3927 17187 3933
rect 17129 3924 17141 3927
rect 17092 3896 17141 3924
rect 17092 3884 17098 3896
rect 17129 3893 17141 3896
rect 17175 3893 17187 3927
rect 17604 3924 17632 3964
rect 17681 3961 17693 3995
rect 17727 3961 17739 3995
rect 17681 3955 17739 3961
rect 18325 3995 18383 4001
rect 18325 3961 18337 3995
rect 18371 3992 18383 3995
rect 19334 3992 19340 4004
rect 18371 3964 19340 3992
rect 18371 3961 18383 3964
rect 18325 3955 18383 3961
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 19794 3952 19800 4004
rect 19852 3992 19858 4004
rect 21634 3992 21640 4004
rect 19852 3964 21640 3992
rect 19852 3952 19858 3964
rect 21634 3952 21640 3964
rect 21692 3952 21698 4004
rect 23308 3992 23336 4091
rect 23382 4088 23388 4140
rect 23440 4128 23446 4140
rect 24581 4131 24639 4137
rect 23440 4100 23485 4128
rect 23440 4088 23446 4100
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 25958 4128 25964 4140
rect 24627 4100 25964 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 25958 4088 25964 4100
rect 26016 4088 26022 4140
rect 27080 4128 27108 4168
rect 26068 4100 27108 4128
rect 27157 4131 27215 4137
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 26068 4060 26096 4100
rect 27157 4097 27169 4131
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27172 4060 27200 4091
rect 24176 4032 26096 4060
rect 27080 4032 27200 4060
rect 27264 4060 27292 4168
rect 27798 4128 27804 4140
rect 27759 4100 27804 4128
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 27893 4063 27951 4069
rect 27893 4060 27905 4063
rect 27264 4032 27905 4060
rect 24176 4020 24182 4032
rect 25590 3992 25596 4004
rect 23308 3964 25596 3992
rect 25590 3952 25596 3964
rect 25648 3952 25654 4004
rect 26418 3992 26424 4004
rect 25700 3964 26424 3992
rect 19702 3924 19708 3936
rect 17604 3896 19708 3924
rect 17129 3887 17187 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 20717 3927 20775 3933
rect 20717 3924 20729 3927
rect 20496 3896 20729 3924
rect 20496 3884 20502 3896
rect 20717 3893 20729 3896
rect 20763 3893 20775 3927
rect 20717 3887 20775 3893
rect 24026 3884 24032 3936
rect 24084 3924 24090 3936
rect 25700 3924 25728 3964
rect 26418 3952 26424 3964
rect 26476 3992 26482 4004
rect 27080 3992 27108 4032
rect 27893 4029 27905 4032
rect 27939 4029 27951 4063
rect 27893 4023 27951 4029
rect 26476 3964 27108 3992
rect 26476 3952 26482 3964
rect 24084 3896 25728 3924
rect 24084 3884 24090 3896
rect 25774 3884 25780 3936
rect 25832 3924 25838 3936
rect 27249 3927 27307 3933
rect 27249 3924 27261 3927
rect 25832 3896 27261 3924
rect 25832 3884 25838 3896
rect 27249 3893 27261 3896
rect 27295 3893 27307 3927
rect 27249 3887 27307 3893
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 12894 3720 12900 3732
rect 12483 3692 12900 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 13449 3723 13507 3729
rect 13449 3689 13461 3723
rect 13495 3720 13507 3723
rect 13722 3720 13728 3732
rect 13495 3692 13728 3720
rect 13495 3689 13507 3692
rect 13449 3683 13507 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14734 3720 14740 3732
rect 14695 3692 14740 3720
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 15562 3720 15568 3732
rect 15523 3692 15568 3720
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19610 3720 19616 3732
rect 18739 3692 19616 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 21450 3720 21456 3732
rect 20548 3692 21456 3720
rect 11793 3655 11851 3661
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 18141 3655 18199 3661
rect 11839 3624 12434 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 12406 3584 12434 3624
rect 18141 3621 18153 3655
rect 18187 3652 18199 3655
rect 18782 3652 18788 3664
rect 18187 3624 18788 3652
rect 18187 3621 18199 3624
rect 18141 3615 18199 3621
rect 18782 3612 18788 3624
rect 18840 3612 18846 3664
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 19392 3624 19441 3652
rect 19392 3612 19398 3624
rect 19429 3621 19441 3624
rect 19475 3621 19487 3655
rect 19429 3615 19487 3621
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 12406 3556 14473 3584
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 20548 3584 20576 3692
rect 21450 3680 21456 3692
rect 21508 3680 21514 3732
rect 21634 3680 21640 3732
rect 21692 3720 21698 3732
rect 22370 3720 22376 3732
rect 21692 3692 22094 3720
rect 22331 3692 22376 3720
rect 21692 3680 21698 3692
rect 21174 3652 21180 3664
rect 21135 3624 21180 3652
rect 21174 3612 21180 3624
rect 21232 3652 21238 3664
rect 21542 3652 21548 3664
rect 21232 3624 21548 3652
rect 21232 3612 21238 3624
rect 21542 3612 21548 3624
rect 21600 3612 21606 3664
rect 22066 3652 22094 3692
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 23624 3692 23765 3720
rect 23624 3680 23630 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 23753 3683 23811 3689
rect 25038 3680 25044 3732
rect 25096 3720 25102 3732
rect 25225 3723 25283 3729
rect 25225 3720 25237 3723
rect 25096 3692 25237 3720
rect 25096 3680 25102 3692
rect 25225 3689 25237 3692
rect 25271 3689 25283 3723
rect 26234 3720 26240 3732
rect 26195 3692 26240 3720
rect 25225 3683 25283 3689
rect 22066 3624 23704 3652
rect 14884 3556 20576 3584
rect 20625 3587 20683 3593
rect 14884 3544 14890 3556
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 3970 3516 3976 3528
rect 1627 3488 3976 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 12124 3488 12633 3516
rect 12124 3476 12130 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13504 3488 13645 3516
rect 13504 3476 13510 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 15194 3516 15200 3528
rect 14323 3488 15200 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15488 3525 15516 3556
rect 20625 3553 20637 3587
rect 20671 3584 20683 3587
rect 21729 3587 21787 3593
rect 21729 3584 21741 3587
rect 20671 3556 21741 3584
rect 20671 3553 20683 3556
rect 20625 3547 20683 3553
rect 21729 3553 21741 3556
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17586 3516 17592 3528
rect 17083 3488 17592 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17920 3488 18061 3516
rect 17920 3476 17926 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 18874 3516 18880 3528
rect 18835 3488 18880 3516
rect 18049 3479 18107 3485
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19576 3488 19625 3516
rect 19576 3476 19582 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 20438 3476 20444 3528
rect 20496 3476 20502 3528
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 23290 3516 23296 3528
rect 22603 3488 23296 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 23676 3525 23704 3624
rect 25240 3584 25268 3683
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 26789 3723 26847 3729
rect 26789 3689 26801 3723
rect 26835 3720 26847 3723
rect 27798 3720 27804 3732
rect 26835 3692 27804 3720
rect 26835 3689 26847 3692
rect 26789 3683 26847 3689
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 25593 3587 25651 3593
rect 25593 3584 25605 3587
rect 25240 3556 25605 3584
rect 25593 3553 25605 3556
rect 25639 3553 25651 3587
rect 25774 3584 25780 3596
rect 25735 3556 25780 3584
rect 25593 3547 25651 3553
rect 25774 3544 25780 3556
rect 25832 3544 25838 3596
rect 23661 3519 23719 3525
rect 23661 3485 23673 3519
rect 23707 3516 23719 3519
rect 25682 3516 25688 3528
rect 23707 3488 25688 3516
rect 23707 3485 23719 3488
rect 23661 3479 23719 3485
rect 25682 3476 25688 3488
rect 25740 3476 25746 3528
rect 26970 3516 26976 3528
rect 26931 3488 26976 3516
rect 26970 3476 26976 3488
rect 27028 3476 27034 3528
rect 27617 3519 27675 3525
rect 27617 3485 27629 3519
rect 27663 3516 27675 3519
rect 27890 3516 27896 3528
rect 27663 3488 27896 3516
rect 27663 3485 27675 3488
rect 27617 3479 27675 3485
rect 27890 3476 27896 3488
rect 27948 3476 27954 3528
rect 28077 3519 28135 3525
rect 28077 3485 28089 3519
rect 28123 3485 28135 3519
rect 28077 3479 28135 3485
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 14182 3448 14188 3460
rect 12492 3420 14188 3448
rect 12492 3408 12498 3420
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 16666 3408 16672 3460
rect 16724 3448 16730 3460
rect 19426 3448 19432 3460
rect 16724 3420 19432 3448
rect 16724 3408 16730 3420
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 20456 3448 20484 3476
rect 20694 3451 20752 3457
rect 20694 3448 20706 3451
rect 20456 3420 20706 3448
rect 20694 3417 20706 3420
rect 20740 3417 20752 3451
rect 28092 3448 28120 3479
rect 20694 3411 20752 3417
rect 27448 3420 28120 3448
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 16853 3383 16911 3389
rect 16853 3349 16865 3383
rect 16899 3380 16911 3383
rect 17494 3380 17500 3392
rect 16899 3352 17500 3380
rect 16899 3349 16911 3352
rect 16853 3343 16911 3349
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 23382 3380 23388 3392
rect 19300 3352 23388 3380
rect 19300 3340 19306 3352
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 27448 3389 27476 3420
rect 27433 3383 27491 3389
rect 27433 3349 27445 3383
rect 27479 3349 27491 3383
rect 27433 3343 27491 3349
rect 28261 3383 28319 3389
rect 28261 3349 28273 3383
rect 28307 3380 28319 3383
rect 29914 3380 29920 3392
rect 28307 3352 29920 3380
rect 28307 3349 28319 3352
rect 28261 3343 28319 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3878 3176 3884 3188
rect 2363 3148 3884 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 5592 3148 9413 3176
rect 5592 3136 5598 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 13633 3179 13691 3185
rect 13633 3176 13645 3179
rect 11940 3148 13645 3176
rect 11940 3136 11946 3148
rect 13633 3145 13645 3148
rect 13679 3145 13691 3179
rect 13633 3139 13691 3145
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 14148 3148 18092 3176
rect 14148 3136 14154 3148
rect 5994 3108 6000 3120
rect 1596 3080 6000 3108
rect 1596 3049 1624 3080
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 12713 3111 12771 3117
rect 12713 3108 12725 3111
rect 10428 3080 12725 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3142 3040 3148 3052
rect 3103 3012 3148 3040
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 5718 3040 5724 3052
rect 5679 3012 5724 3040
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 10428 3049 10456 3080
rect 12713 3077 12725 3080
rect 12759 3077 12771 3111
rect 12713 3071 12771 3077
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 18064 3108 18092 3148
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 18196 3148 18245 3176
rect 18196 3136 18202 3148
rect 18233 3145 18245 3148
rect 18279 3145 18291 3179
rect 18233 3139 18291 3145
rect 18874 3136 18880 3188
rect 18932 3176 18938 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 18932 3148 20637 3176
rect 18932 3136 18938 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 20625 3139 20683 3145
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 22005 3179 22063 3185
rect 22005 3176 22017 3179
rect 20864 3148 22017 3176
rect 20864 3136 20870 3148
rect 22005 3145 22017 3148
rect 22051 3145 22063 3179
rect 22005 3139 22063 3145
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 23382 3176 23388 3188
rect 22244 3148 22692 3176
rect 23343 3148 23388 3176
rect 22244 3136 22250 3148
rect 19794 3108 19800 3120
rect 15988 3080 17540 3108
rect 18064 3080 19800 3108
rect 15988 3068 15994 3080
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 8987 3012 9597 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12158 3040 12164 3052
rect 12023 3012 12164 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 8386 2972 8392 2984
rect 2976 2944 8392 2972
rect 2976 2913 3004 2944
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8864 2972 8892 3003
rect 11164 2972 11192 3003
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 13078 3040 13084 3052
rect 12667 3012 13084 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 14550 3040 14556 3052
rect 13863 3012 14556 3040
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 16666 3040 16672 3052
rect 15795 3012 16672 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 8864 2944 11100 2972
rect 11164 2944 12081 2972
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2873 3019 2907
rect 2961 2867 3019 2873
rect 7650 2864 7656 2916
rect 7708 2904 7714 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 7708 2876 10977 2904
rect 7708 2864 7714 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 10965 2867 11023 2873
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 5718 2836 5724 2848
rect 5583 2808 5724 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10410 2836 10416 2848
rect 10275 2808 10416 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 11072 2836 11100 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 14844 2972 14872 3003
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17512 3049 17540 3080
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 18141 3043 18199 3049
rect 17644 3012 17689 3040
rect 17644 3000 17650 3012
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18230 3040 18236 3052
rect 18187 3012 18236 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 14844 2944 15853 2972
rect 12069 2935 12127 2941
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 11238 2864 11244 2916
rect 11296 2904 11302 2916
rect 18156 2904 18184 3003
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 18984 3049 19012 3080
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 20640 3080 22094 3108
rect 20640 3052 20668 3080
rect 18969 3043 19027 3049
rect 18969 3009 18981 3043
rect 19015 3009 19027 3043
rect 18969 3003 19027 3009
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 20806 3040 20812 3052
rect 20767 3012 20812 3040
rect 20806 3000 20812 3012
rect 20864 3040 20870 3052
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 20864 3012 21281 3040
rect 20864 3000 20870 3012
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 22066 3040 22094 3080
rect 22664 3049 22692 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 25130 3136 25136 3188
rect 25188 3176 25194 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 25188 3148 25513 3176
rect 25188 3136 25194 3148
rect 25501 3145 25513 3148
rect 25547 3145 25559 3179
rect 25501 3139 25559 3145
rect 27433 3179 27491 3185
rect 27433 3145 27445 3179
rect 27479 3176 27491 3179
rect 27522 3176 27528 3188
rect 27479 3148 27528 3176
rect 27479 3145 27491 3148
rect 27433 3139 27491 3145
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 25866 3108 25872 3120
rect 23308 3080 25872 3108
rect 23308 3049 23336 3080
rect 25866 3068 25872 3080
rect 25924 3068 25930 3120
rect 22189 3043 22247 3049
rect 22189 3040 22201 3043
rect 22066 3012 22201 3040
rect 21269 3003 21327 3009
rect 22189 3009 22201 3012
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 23293 3043 23351 3049
rect 23293 3009 23305 3043
rect 23339 3009 23351 3043
rect 23293 3003 23351 3009
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 24305 3043 24363 3049
rect 24305 3009 24317 3043
rect 24351 3040 24363 3043
rect 25041 3043 25099 3049
rect 25041 3040 25053 3043
rect 24351 3012 25053 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 25041 3009 25053 3012
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 25685 3043 25743 3049
rect 25685 3009 25697 3043
rect 25731 3040 25743 3043
rect 26418 3040 26424 3052
rect 25731 3012 26280 3040
rect 26379 3012 26424 3040
rect 25731 3009 25743 3012
rect 25685 3003 25743 3009
rect 19518 2972 19524 2984
rect 19479 2944 19524 2972
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 19705 2975 19763 2981
rect 19705 2941 19717 2975
rect 19751 2972 19763 2975
rect 21361 2975 21419 2981
rect 21361 2972 21373 2975
rect 19751 2944 21373 2972
rect 19751 2941 19763 2944
rect 19705 2935 19763 2941
rect 21361 2941 21373 2944
rect 21407 2941 21419 2975
rect 21361 2935 21419 2941
rect 21542 2932 21548 2984
rect 21600 2972 21606 2984
rect 24228 2972 24256 3003
rect 21600 2944 24256 2972
rect 21600 2932 21606 2944
rect 11296 2876 18184 2904
rect 11296 2864 11302 2876
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 21450 2904 21456 2916
rect 19392 2876 21456 2904
rect 19392 2864 19398 2876
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 26252 2913 26280 3012
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 27617 3043 27675 3049
rect 27617 3009 27629 3043
rect 27663 3009 27675 3043
rect 28074 3040 28080 3052
rect 28035 3012 28080 3040
rect 27617 3003 27675 3009
rect 27632 2972 27660 3003
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 29086 2972 29092 2984
rect 27632 2944 29092 2972
rect 29086 2932 29092 2944
rect 29144 2932 29150 2984
rect 26237 2907 26295 2913
rect 26237 2873 26249 2907
rect 26283 2873 26295 2907
rect 26237 2867 26295 2873
rect 12342 2836 12348 2848
rect 11072 2808 12348 2836
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 14642 2836 14648 2848
rect 14603 2808 14648 2836
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 15804 2808 16865 2836
rect 15804 2796 15810 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 18782 2836 18788 2848
rect 18743 2808 18788 2836
rect 16853 2799 16911 2805
rect 18782 2796 18788 2808
rect 18840 2796 18846 2848
rect 19702 2796 19708 2848
rect 19760 2836 19766 2848
rect 19889 2839 19947 2845
rect 19889 2836 19901 2839
rect 19760 2808 19901 2836
rect 19760 2796 19766 2808
rect 19889 2805 19901 2808
rect 19935 2805 19947 2839
rect 19889 2799 19947 2805
rect 20254 2796 20260 2848
rect 20312 2836 20318 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 20312 2808 22753 2836
rect 20312 2796 20318 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 22741 2799 22799 2805
rect 24857 2839 24915 2845
rect 24857 2805 24869 2839
rect 24903 2836 24915 2839
rect 27798 2836 27804 2848
rect 24903 2808 27804 2836
rect 24903 2805 24915 2808
rect 24857 2799 24915 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28261 2839 28319 2845
rect 28261 2805 28273 2839
rect 28307 2836 28319 2839
rect 28350 2836 28356 2848
rect 28307 2808 28356 2836
rect 28307 2805 28319 2808
rect 28261 2799 28319 2805
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 7837 2635 7895 2641
rect 7837 2601 7849 2635
rect 7883 2632 7895 2635
rect 9030 2632 9036 2644
rect 7883 2604 9036 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9306 2632 9312 2644
rect 9171 2604 9312 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11204 2604 11713 2632
rect 11204 2592 11210 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 11701 2595 11759 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 18233 2635 18291 2641
rect 18233 2601 18245 2635
rect 18279 2632 18291 2635
rect 18690 2632 18696 2644
rect 18279 2604 18696 2632
rect 18279 2601 18291 2604
rect 18233 2595 18291 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 19576 2604 19717 2632
rect 19576 2592 19582 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 20530 2632 20536 2644
rect 20491 2604 20536 2632
rect 19705 2595 19763 2601
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 22646 2632 22652 2644
rect 22607 2604 22652 2632
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 24578 2632 24584 2644
rect 24539 2604 24584 2632
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 25866 2632 25872 2644
rect 25827 2604 25872 2632
rect 25866 2592 25872 2604
rect 25924 2592 25930 2644
rect 25958 2592 25964 2644
rect 26016 2632 26022 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 26016 2604 27169 2632
rect 26016 2592 26022 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 4246 2564 4252 2576
rect 1596 2536 4252 2564
rect 1596 2437 1624 2536
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 21085 2567 21143 2573
rect 21085 2533 21097 2567
rect 21131 2533 21143 2567
rect 21085 2527 21143 2533
rect 14458 2496 14464 2508
rect 3160 2468 14464 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 3160 2437 3188 2468
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 21100 2496 21128 2527
rect 22278 2524 22284 2576
rect 22336 2564 22342 2576
rect 23293 2567 23351 2573
rect 23293 2564 23305 2567
rect 22336 2536 23305 2564
rect 22336 2524 22342 2536
rect 23293 2533 23305 2536
rect 23339 2533 23351 2567
rect 23293 2527 23351 2533
rect 25225 2567 25283 2573
rect 25225 2533 25237 2567
rect 25271 2564 25283 2567
rect 27246 2564 27252 2576
rect 25271 2536 27252 2564
rect 25271 2533 25283 2536
rect 25225 2527 25283 2533
rect 27246 2524 27252 2536
rect 27304 2524 27310 2576
rect 19904 2468 21128 2496
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2004 2400 2513 2428
rect 2004 2388 2010 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 5534 2428 5540 2440
rect 4663 2400 5540 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5718 2428 5724 2440
rect 5679 2400 5724 2428
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 7650 2428 7656 2440
rect 6595 2400 7656 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9088 2400 9321 2428
rect 9088 2388 9094 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 9309 2391 9367 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11664 2400 11897 2428
rect 11664 2388 11670 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12308 2400 12725 2428
rect 12308 2388 12314 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 14642 2428 14648 2440
rect 13495 2400 14648 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15746 2428 15752 2440
rect 14967 2400 15752 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16172 2400 17049 2428
rect 16172 2388 16178 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17037 2391 17095 2397
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2428 18475 2431
rect 18782 2428 18788 2440
rect 18463 2400 18788 2428
rect 18463 2397 18475 2400
rect 18417 2391 18475 2397
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 19904 2437 19932 2468
rect 19889 2431 19947 2437
rect 19889 2397 19901 2431
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 11790 2360 11796 2372
rect 2332 2332 11796 2360
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 2332 2301 2360 2332
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 20456 2360 20484 2391
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 20588 2400 21281 2428
rect 20588 2388 20594 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21508 2400 22201 2428
rect 21508 2388 21514 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22336 2400 22845 2428
rect 22336 2388 22342 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23256 2400 23489 2428
rect 23256 2388 23262 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 25406 2428 25412 2440
rect 25367 2400 25412 2428
rect 24765 2391 24823 2397
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25832 2400 26065 2428
rect 25832 2388 25838 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 26476 2400 27353 2428
rect 26476 2388 26482 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27798 2428 27804 2440
rect 27759 2400 27804 2428
rect 27341 2391 27399 2397
rect 27798 2388 27804 2400
rect 27856 2388 27862 2440
rect 20456 2332 22048 2360
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 72 2264 1777 2292
rect 72 2252 78 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 1765 2255 1823 2261
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2261 2375 2295
rect 2317 2255 2375 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4580 2264 4813 2292
rect 4580 2252 4586 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5868 2264 5917 2292
rect 5868 2252 5874 2264
rect 5905 2261 5917 2264
rect 5951 2261 5963 2295
rect 5905 2255 5963 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 12894 2292 12900 2304
rect 12855 2264 12900 2292
rect 10597 2255 10655 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13596 2264 13645 2292
rect 13596 2252 13602 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14792 2264 15117 2292
rect 14792 2252 14798 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 22020 2301 22048 2332
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 18690 1368 18696 1420
rect 18748 1408 18754 1420
rect 20530 1408 20536 1420
rect 18748 1380 20536 1408
rect 18748 1368 18754 1380
rect 20530 1368 20536 1380
rect 20588 1368 20594 1420
<< via1 >>
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 1032 27548 1084 27600
rect 6092 27548 6144 27600
rect 7288 27480 7340 27532
rect 10324 27548 10376 27600
rect 13544 27548 13596 27600
rect 15108 27591 15160 27600
rect 15108 27557 15117 27591
rect 15117 27557 15151 27591
rect 15151 27557 15160 27591
rect 15108 27548 15160 27557
rect 16120 27548 16172 27600
rect 18052 27548 18104 27600
rect 3240 27412 3292 27464
rect 3424 27455 3476 27464
rect 3424 27421 3433 27455
rect 3433 27421 3467 27455
rect 3467 27421 3476 27455
rect 3424 27412 3476 27421
rect 4160 27455 4212 27464
rect 4160 27421 4169 27455
rect 4169 27421 4203 27455
rect 4203 27421 4212 27455
rect 4160 27412 4212 27421
rect 5448 27455 5500 27464
rect 5448 27421 5457 27455
rect 5457 27421 5491 27455
rect 5491 27421 5500 27455
rect 5448 27412 5500 27421
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 8024 27455 8076 27464
rect 8024 27421 8033 27455
rect 8033 27421 8067 27455
rect 8067 27421 8076 27455
rect 8024 27412 8076 27421
rect 9036 27412 9088 27464
rect 10416 27455 10468 27464
rect 10416 27421 10425 27455
rect 10425 27421 10459 27455
rect 10459 27421 10468 27455
rect 10416 27412 10468 27421
rect 11060 27412 11112 27464
rect 12440 27412 12492 27464
rect 13176 27412 13228 27464
rect 14372 27412 14424 27464
rect 16856 27455 16908 27464
rect 1676 27387 1728 27396
rect 1676 27353 1685 27387
rect 1685 27353 1719 27387
rect 1719 27353 1728 27387
rect 1676 27344 1728 27353
rect 1860 27387 1912 27396
rect 1860 27353 1869 27387
rect 1869 27353 1903 27387
rect 1903 27353 1912 27387
rect 1860 27344 1912 27353
rect 6460 27276 6512 27328
rect 11980 27344 12032 27396
rect 16856 27421 16865 27455
rect 16865 27421 16899 27455
rect 16899 27421 16908 27455
rect 16856 27412 16908 27421
rect 20720 27548 20772 27600
rect 23480 27548 23532 27600
rect 19616 27455 19668 27464
rect 19616 27421 19625 27455
rect 19625 27421 19659 27455
rect 19659 27421 19668 27455
rect 19616 27412 19668 27421
rect 17776 27344 17828 27396
rect 9588 27276 9640 27328
rect 11704 27319 11756 27328
rect 11704 27285 11713 27319
rect 11713 27285 11747 27319
rect 11747 27285 11756 27319
rect 11704 27276 11756 27285
rect 12716 27276 12768 27328
rect 14740 27276 14792 27328
rect 15660 27319 15712 27328
rect 15660 27285 15669 27319
rect 15669 27285 15703 27319
rect 15703 27285 15712 27319
rect 15660 27276 15712 27285
rect 15936 27276 15988 27328
rect 21364 27412 21416 27464
rect 22100 27412 22152 27464
rect 27528 27616 27580 27668
rect 29276 27616 29328 27668
rect 27712 27548 27764 27600
rect 25136 27480 25188 27532
rect 24216 27344 24268 27396
rect 26424 27412 26476 27464
rect 27436 27412 27488 27464
rect 21548 27276 21600 27328
rect 21640 27276 21692 27328
rect 22652 27319 22704 27328
rect 22652 27285 22661 27319
rect 22661 27285 22695 27319
rect 22695 27285 22704 27319
rect 22652 27276 22704 27285
rect 23388 27319 23440 27328
rect 23388 27285 23397 27319
rect 23397 27285 23431 27319
rect 23431 27285 23440 27319
rect 23388 27276 23440 27285
rect 25044 27276 25096 27328
rect 25596 27276 25648 27328
rect 27160 27319 27212 27328
rect 27160 27285 27169 27319
rect 27169 27285 27203 27319
rect 27203 27285 27212 27319
rect 27160 27276 27212 27285
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 2780 27072 2832 27124
rect 3240 27072 3292 27124
rect 13176 27115 13228 27124
rect 13176 27081 13185 27115
rect 13185 27081 13219 27115
rect 13219 27081 13228 27115
rect 13176 27072 13228 27081
rect 1952 26936 2004 26988
rect 3148 26979 3200 26988
rect 3148 26945 3157 26979
rect 3157 26945 3191 26979
rect 3191 26945 3200 26979
rect 3148 26936 3200 26945
rect 4252 26936 4304 26988
rect 13912 26936 13964 26988
rect 15660 27004 15712 27056
rect 4896 26868 4948 26920
rect 11796 26868 11848 26920
rect 14740 26936 14792 26988
rect 19340 27072 19392 27124
rect 27528 27115 27580 27124
rect 27528 27081 27537 27115
rect 27537 27081 27571 27115
rect 27571 27081 27580 27115
rect 27528 27072 27580 27081
rect 29920 27072 29972 27124
rect 16764 27004 16816 27056
rect 17132 26936 17184 26988
rect 17776 26979 17828 26988
rect 17776 26945 17785 26979
rect 17785 26945 17819 26979
rect 17819 26945 17828 26979
rect 17776 26936 17828 26945
rect 18788 27004 18840 27056
rect 22652 27004 22704 27056
rect 19432 26936 19484 26988
rect 19708 26936 19760 26988
rect 21640 26936 21692 26988
rect 23020 26936 23072 26988
rect 27160 27004 27212 27056
rect 16948 26868 17000 26920
rect 17684 26868 17736 26920
rect 8300 26800 8352 26852
rect 10416 26800 10468 26852
rect 14280 26800 14332 26852
rect 16120 26800 16172 26852
rect 10232 26732 10284 26784
rect 13820 26775 13872 26784
rect 13820 26741 13829 26775
rect 13829 26741 13863 26775
rect 13863 26741 13872 26775
rect 13820 26732 13872 26741
rect 14556 26775 14608 26784
rect 14556 26741 14565 26775
rect 14565 26741 14599 26775
rect 14599 26741 14608 26775
rect 14556 26732 14608 26741
rect 15752 26775 15804 26784
rect 15752 26741 15761 26775
rect 15761 26741 15795 26775
rect 15795 26741 15804 26775
rect 15752 26732 15804 26741
rect 16672 26732 16724 26784
rect 18696 26732 18748 26784
rect 19708 26800 19760 26852
rect 20720 26868 20772 26920
rect 22652 26868 22704 26920
rect 26516 26936 26568 26988
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 27344 26936 27396 26945
rect 27528 26936 27580 26988
rect 27896 26868 27948 26920
rect 23388 26800 23440 26852
rect 19892 26732 19944 26784
rect 21180 26775 21232 26784
rect 21180 26741 21189 26775
rect 21189 26741 21223 26775
rect 21223 26741 21232 26775
rect 21180 26732 21232 26741
rect 22560 26775 22612 26784
rect 22560 26741 22569 26775
rect 22569 26741 22603 26775
rect 22603 26741 22612 26775
rect 22560 26732 22612 26741
rect 22744 26732 22796 26784
rect 23848 26775 23900 26784
rect 23848 26741 23857 26775
rect 23857 26741 23891 26775
rect 23891 26741 23900 26775
rect 23848 26732 23900 26741
rect 24492 26775 24544 26784
rect 24492 26741 24501 26775
rect 24501 26741 24535 26775
rect 24535 26741 24544 26775
rect 24492 26732 24544 26741
rect 25964 26732 26016 26784
rect 26056 26775 26108 26784
rect 26056 26741 26065 26775
rect 26065 26741 26099 26775
rect 26099 26741 26108 26775
rect 26056 26732 26108 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 4252 26571 4304 26580
rect 4252 26537 4261 26571
rect 4261 26537 4295 26571
rect 4295 26537 4304 26571
rect 4252 26528 4304 26537
rect 4896 26571 4948 26580
rect 4896 26537 4905 26571
rect 4905 26537 4939 26571
rect 4939 26537 4948 26571
rect 4896 26528 4948 26537
rect 11888 26528 11940 26580
rect 16948 26528 17000 26580
rect 19432 26571 19484 26580
rect 19432 26537 19441 26571
rect 19441 26537 19475 26571
rect 19475 26537 19484 26571
rect 19432 26528 19484 26537
rect 19616 26528 19668 26580
rect 20720 26571 20772 26580
rect 20720 26537 20729 26571
rect 20729 26537 20763 26571
rect 20763 26537 20772 26571
rect 20720 26528 20772 26537
rect 21364 26571 21416 26580
rect 21364 26537 21373 26571
rect 21373 26537 21407 26571
rect 21407 26537 21416 26571
rect 21364 26528 21416 26537
rect 22652 26571 22704 26580
rect 22652 26537 22661 26571
rect 22661 26537 22695 26571
rect 22695 26537 22704 26571
rect 22652 26528 22704 26537
rect 27344 26571 27396 26580
rect 27344 26537 27353 26571
rect 27353 26537 27387 26571
rect 27387 26537 27396 26571
rect 27344 26528 27396 26537
rect 28632 26528 28684 26580
rect 9312 26460 9364 26512
rect 1768 26367 1820 26376
rect 1768 26333 1777 26367
rect 1777 26333 1811 26367
rect 1811 26333 1820 26367
rect 1768 26324 1820 26333
rect 5080 26367 5132 26376
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 5080 26324 5132 26333
rect 15292 26460 15344 26512
rect 18880 26460 18932 26512
rect 11980 26367 12032 26376
rect 11980 26333 11989 26367
rect 11989 26333 12023 26367
rect 12023 26333 12032 26367
rect 11980 26324 12032 26333
rect 12716 26367 12768 26376
rect 12716 26333 12725 26367
rect 12725 26333 12759 26367
rect 12759 26333 12768 26367
rect 12716 26324 12768 26333
rect 13820 26392 13872 26444
rect 16672 26435 16724 26444
rect 16672 26401 16681 26435
rect 16681 26401 16715 26435
rect 16715 26401 16724 26435
rect 16672 26392 16724 26401
rect 14188 26324 14240 26376
rect 15752 26324 15804 26376
rect 18788 26392 18840 26444
rect 12256 26256 12308 26308
rect 18972 26324 19024 26376
rect 19432 26324 19484 26376
rect 19064 26256 19116 26308
rect 20168 26324 20220 26376
rect 21548 26367 21600 26376
rect 21548 26333 21557 26367
rect 21557 26333 21591 26367
rect 21591 26333 21600 26367
rect 21548 26324 21600 26333
rect 22744 26324 22796 26376
rect 25872 26460 25924 26512
rect 25964 26392 26016 26444
rect 21456 26256 21508 26308
rect 23572 26324 23624 26376
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26884 26367 26936 26376
rect 26884 26333 26893 26367
rect 26893 26333 26927 26367
rect 26927 26333 26936 26367
rect 26884 26324 26936 26333
rect 27252 26324 27304 26376
rect 26516 26256 26568 26308
rect 11980 26188 12032 26240
rect 12440 26188 12492 26240
rect 13360 26188 13412 26240
rect 18144 26231 18196 26240
rect 18144 26197 18153 26231
rect 18153 26197 18187 26231
rect 18187 26197 18196 26231
rect 18144 26188 18196 26197
rect 22836 26188 22888 26240
rect 24952 26231 25004 26240
rect 24952 26197 24961 26231
rect 24961 26197 24995 26231
rect 24995 26197 25004 26231
rect 24952 26188 25004 26197
rect 26700 26231 26752 26240
rect 26700 26197 26709 26231
rect 26709 26197 26743 26231
rect 26743 26197 26752 26231
rect 26700 26188 26752 26197
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 5080 25984 5132 26036
rect 13912 25984 13964 26036
rect 27528 26027 27580 26036
rect 27528 25993 27537 26027
rect 27537 25993 27571 26027
rect 27571 25993 27580 26027
rect 27528 25984 27580 25993
rect 11796 25959 11848 25968
rect 11796 25925 11805 25959
rect 11805 25925 11839 25959
rect 11839 25925 11848 25959
rect 11796 25916 11848 25925
rect 11888 25959 11940 25968
rect 11888 25925 11897 25959
rect 11897 25925 11931 25959
rect 11931 25925 11940 25959
rect 13360 25959 13412 25968
rect 11888 25916 11940 25925
rect 13360 25925 13369 25959
rect 13369 25925 13403 25959
rect 13403 25925 13412 25959
rect 13360 25916 13412 25925
rect 6460 25848 6512 25900
rect 9772 25848 9824 25900
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 15292 25848 15344 25900
rect 17224 25848 17276 25900
rect 19432 25916 19484 25968
rect 20996 25891 21048 25900
rect 20996 25857 21005 25891
rect 21005 25857 21039 25891
rect 21039 25857 21048 25891
rect 20996 25848 21048 25857
rect 21088 25848 21140 25900
rect 24952 25848 25004 25900
rect 26700 25848 26752 25900
rect 27712 25891 27764 25900
rect 27712 25857 27721 25891
rect 27721 25857 27755 25891
rect 27755 25857 27764 25891
rect 27712 25848 27764 25857
rect 13268 25823 13320 25832
rect 13268 25789 13277 25823
rect 13277 25789 13311 25823
rect 13311 25789 13320 25823
rect 13268 25780 13320 25789
rect 18236 25780 18288 25832
rect 18696 25823 18748 25832
rect 18696 25789 18705 25823
rect 18705 25789 18739 25823
rect 18739 25789 18748 25823
rect 18696 25780 18748 25789
rect 22652 25823 22704 25832
rect 22652 25789 22661 25823
rect 22661 25789 22695 25823
rect 22695 25789 22704 25823
rect 22652 25780 22704 25789
rect 24124 25780 24176 25832
rect 27528 25780 27580 25832
rect 11244 25644 11296 25696
rect 11888 25644 11940 25696
rect 14280 25644 14332 25696
rect 15108 25644 15160 25696
rect 21548 25712 21600 25764
rect 24768 25712 24820 25764
rect 17132 25687 17184 25696
rect 17132 25653 17141 25687
rect 17141 25653 17175 25687
rect 17175 25653 17184 25687
rect 17132 25644 17184 25653
rect 17960 25687 18012 25696
rect 17960 25653 17969 25687
rect 17969 25653 18003 25687
rect 18003 25653 18012 25687
rect 17960 25644 18012 25653
rect 18880 25687 18932 25696
rect 18880 25653 18889 25687
rect 18889 25653 18923 25687
rect 18923 25653 18932 25687
rect 18880 25644 18932 25653
rect 21364 25644 21416 25696
rect 22100 25687 22152 25696
rect 22100 25653 22109 25687
rect 22109 25653 22143 25687
rect 22143 25653 22152 25687
rect 22100 25644 22152 25653
rect 23388 25644 23440 25696
rect 25688 25687 25740 25696
rect 25688 25653 25697 25687
rect 25697 25653 25731 25687
rect 25731 25653 25740 25687
rect 25688 25644 25740 25653
rect 27344 25644 27396 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 13912 25440 13964 25492
rect 14372 25483 14424 25492
rect 14372 25449 14381 25483
rect 14381 25449 14415 25483
rect 14415 25449 14424 25483
rect 14372 25440 14424 25449
rect 16856 25440 16908 25492
rect 18236 25440 18288 25492
rect 21548 25483 21600 25492
rect 21548 25449 21557 25483
rect 21557 25449 21591 25483
rect 21591 25449 21600 25483
rect 21548 25440 21600 25449
rect 27436 25440 27488 25492
rect 27896 25483 27948 25492
rect 27896 25449 27905 25483
rect 27905 25449 27939 25483
rect 27939 25449 27948 25483
rect 27896 25440 27948 25449
rect 13176 25372 13228 25424
rect 13268 25372 13320 25424
rect 11152 25279 11204 25288
rect 11152 25245 11161 25279
rect 11161 25245 11195 25279
rect 11195 25245 11204 25279
rect 11152 25236 11204 25245
rect 11704 25236 11756 25288
rect 13084 25279 13136 25288
rect 11060 25168 11112 25220
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 13728 25236 13780 25288
rect 17132 25304 17184 25356
rect 16488 25279 16540 25288
rect 16488 25245 16497 25279
rect 16497 25245 16531 25279
rect 16531 25245 16540 25279
rect 16488 25236 16540 25245
rect 15108 25211 15160 25220
rect 15108 25177 15117 25211
rect 15117 25177 15151 25211
rect 15151 25177 15160 25211
rect 15108 25168 15160 25177
rect 15752 25211 15804 25220
rect 10324 25143 10376 25152
rect 10324 25109 10333 25143
rect 10333 25109 10367 25143
rect 10367 25109 10376 25143
rect 10324 25100 10376 25109
rect 11796 25100 11848 25152
rect 12624 25100 12676 25152
rect 14096 25100 14148 25152
rect 14372 25100 14424 25152
rect 15752 25177 15761 25211
rect 15761 25177 15795 25211
rect 15795 25177 15804 25211
rect 15752 25168 15804 25177
rect 18144 25236 18196 25288
rect 18972 25236 19024 25288
rect 19984 25236 20036 25288
rect 20260 25236 20312 25288
rect 25688 25372 25740 25424
rect 21364 25347 21416 25356
rect 21364 25313 21373 25347
rect 21373 25313 21407 25347
rect 21407 25313 21416 25347
rect 21364 25304 21416 25313
rect 23756 25304 23808 25356
rect 22744 25279 22796 25288
rect 19248 25168 19300 25220
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 24492 25236 24544 25288
rect 25044 25236 25096 25288
rect 25412 25279 25464 25288
rect 25412 25245 25421 25279
rect 25421 25245 25455 25279
rect 25455 25245 25464 25279
rect 25412 25236 25464 25245
rect 25504 25236 25556 25288
rect 26792 25236 26844 25288
rect 27804 25279 27856 25288
rect 27804 25245 27813 25279
rect 27813 25245 27847 25279
rect 27847 25245 27856 25279
rect 27804 25236 27856 25245
rect 20168 25100 20220 25152
rect 28172 25168 28224 25220
rect 23204 25100 23256 25152
rect 25136 25100 25188 25152
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 11980 24896 12032 24948
rect 15752 24896 15804 24948
rect 1768 24803 1820 24812
rect 1768 24769 1777 24803
rect 1777 24769 1811 24803
rect 1811 24769 1820 24803
rect 1768 24760 1820 24769
rect 8392 24760 8444 24812
rect 9864 24803 9916 24812
rect 9864 24769 9873 24803
rect 9873 24769 9907 24803
rect 9907 24769 9916 24803
rect 9864 24760 9916 24769
rect 10692 24760 10744 24812
rect 11796 24760 11848 24812
rect 13176 24760 13228 24812
rect 14096 24803 14148 24812
rect 14096 24769 14105 24803
rect 14105 24769 14139 24803
rect 14139 24769 14148 24803
rect 14096 24760 14148 24769
rect 14556 24760 14608 24812
rect 20904 24896 20956 24948
rect 10876 24692 10928 24744
rect 16488 24692 16540 24744
rect 20168 24760 20220 24812
rect 18788 24692 18840 24744
rect 19248 24692 19300 24744
rect 19800 24692 19852 24744
rect 21088 24760 21140 24812
rect 22744 24828 22796 24880
rect 23940 24828 23992 24880
rect 23848 24760 23900 24812
rect 25412 24871 25464 24880
rect 25412 24837 25421 24871
rect 25421 24837 25455 24871
rect 25455 24837 25464 24871
rect 25412 24828 25464 24837
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 27344 24760 27396 24812
rect 28172 24803 28224 24812
rect 28172 24769 28181 24803
rect 28181 24769 28215 24803
rect 28215 24769 28224 24803
rect 28172 24760 28224 24769
rect 21272 24692 21324 24744
rect 22192 24735 22244 24744
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 9772 24624 9824 24676
rect 11152 24624 11204 24676
rect 23296 24692 23348 24744
rect 26056 24692 26108 24744
rect 22928 24624 22980 24676
rect 25504 24624 25556 24676
rect 4068 24556 4120 24608
rect 11060 24556 11112 24608
rect 12992 24556 13044 24608
rect 14648 24556 14700 24608
rect 19340 24556 19392 24608
rect 19524 24599 19576 24608
rect 19524 24565 19533 24599
rect 19533 24565 19567 24599
rect 19567 24565 19576 24599
rect 19524 24556 19576 24565
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 20812 24599 20864 24608
rect 20812 24565 20821 24599
rect 20821 24565 20855 24599
rect 20855 24565 20864 24599
rect 20812 24556 20864 24565
rect 22560 24556 22612 24608
rect 24584 24556 24636 24608
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 26056 24556 26108 24608
rect 28540 24556 28592 24608
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 13084 24352 13136 24404
rect 14372 24352 14424 24404
rect 17684 24352 17736 24404
rect 9864 24284 9916 24336
rect 10324 24216 10376 24268
rect 11980 24216 12032 24268
rect 8392 24191 8444 24200
rect 8392 24157 8401 24191
rect 8401 24157 8435 24191
rect 8435 24157 8444 24191
rect 8392 24148 8444 24157
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 16304 24284 16356 24336
rect 19156 24284 19208 24336
rect 20996 24352 21048 24404
rect 22192 24352 22244 24404
rect 24768 24352 24820 24404
rect 27252 24395 27304 24404
rect 19616 24284 19668 24336
rect 19800 24284 19852 24336
rect 22928 24327 22980 24336
rect 22928 24293 22937 24327
rect 22937 24293 22971 24327
rect 22971 24293 22980 24327
rect 22928 24284 22980 24293
rect 23112 24284 23164 24336
rect 27252 24361 27261 24395
rect 27261 24361 27295 24395
rect 27295 24361 27304 24395
rect 27252 24352 27304 24361
rect 27712 24352 27764 24404
rect 19708 24216 19760 24268
rect 20076 24216 20128 24268
rect 12808 24191 12860 24200
rect 12808 24157 12817 24191
rect 12817 24157 12851 24191
rect 12851 24157 12860 24191
rect 12808 24148 12860 24157
rect 13176 24148 13228 24200
rect 15292 24148 15344 24200
rect 16120 24191 16172 24200
rect 16120 24157 16129 24191
rect 16129 24157 16163 24191
rect 16163 24157 16172 24191
rect 16120 24148 16172 24157
rect 10600 24012 10652 24064
rect 12624 24012 12676 24064
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 15200 24012 15252 24064
rect 18144 24148 18196 24200
rect 18788 24148 18840 24200
rect 19616 24148 19668 24200
rect 19984 24148 20036 24200
rect 21456 24148 21508 24200
rect 23388 24216 23440 24268
rect 24584 24259 24636 24268
rect 24584 24225 24593 24259
rect 24593 24225 24627 24259
rect 24627 24225 24636 24259
rect 24584 24216 24636 24225
rect 26056 24259 26108 24268
rect 23112 24148 23164 24200
rect 23572 24148 23624 24200
rect 23848 24148 23900 24200
rect 25688 24148 25740 24200
rect 18604 24012 18656 24064
rect 19156 24012 19208 24064
rect 25504 24080 25556 24132
rect 26056 24225 26065 24259
rect 26065 24225 26099 24259
rect 26099 24225 26108 24259
rect 26056 24216 26108 24225
rect 26424 24148 26476 24200
rect 19616 24012 19668 24064
rect 20444 24012 20496 24064
rect 22192 24012 22244 24064
rect 25228 24012 25280 24064
rect 25320 24012 25372 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 9220 23808 9272 23860
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 9312 23715 9364 23724
rect 9312 23681 9321 23715
rect 9321 23681 9355 23715
rect 9355 23681 9364 23715
rect 9312 23672 9364 23681
rect 11060 23672 11112 23724
rect 8392 23604 8444 23656
rect 12900 23672 12952 23724
rect 10692 23536 10744 23588
rect 10416 23468 10468 23520
rect 12992 23604 13044 23656
rect 15936 23740 15988 23792
rect 18880 23740 18932 23792
rect 19156 23783 19208 23792
rect 19156 23749 19165 23783
rect 19165 23749 19199 23783
rect 19199 23749 19208 23783
rect 19156 23740 19208 23749
rect 19708 23808 19760 23860
rect 22652 23808 22704 23860
rect 24124 23808 24176 23860
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 22468 23740 22520 23792
rect 23296 23783 23348 23792
rect 23296 23749 23305 23783
rect 23305 23749 23339 23783
rect 23339 23749 23348 23783
rect 23296 23740 23348 23749
rect 24676 23740 24728 23792
rect 15476 23672 15528 23724
rect 16948 23672 17000 23724
rect 17684 23672 17736 23724
rect 17960 23672 18012 23724
rect 20168 23715 20220 23724
rect 20168 23681 20177 23715
rect 20177 23681 20211 23715
rect 20211 23681 20220 23715
rect 20168 23672 20220 23681
rect 21088 23672 21140 23724
rect 25596 23740 25648 23792
rect 25044 23715 25096 23724
rect 14648 23647 14700 23656
rect 14648 23613 14657 23647
rect 14657 23613 14691 23647
rect 14691 23613 14700 23647
rect 14648 23604 14700 23613
rect 15384 23604 15436 23656
rect 16212 23604 16264 23656
rect 19432 23604 19484 23656
rect 19524 23647 19576 23656
rect 19524 23613 19533 23647
rect 19533 23613 19567 23647
rect 19567 23613 19576 23647
rect 19524 23604 19576 23613
rect 19708 23604 19760 23656
rect 11796 23468 11848 23520
rect 14924 23468 14976 23520
rect 18788 23536 18840 23588
rect 20536 23604 20588 23656
rect 22192 23604 22244 23656
rect 25044 23681 25053 23715
rect 25053 23681 25087 23715
rect 25087 23681 25096 23715
rect 25044 23672 25096 23681
rect 25136 23672 25188 23724
rect 26056 23672 26108 23724
rect 28356 23715 28408 23724
rect 28356 23681 28365 23715
rect 28365 23681 28399 23715
rect 28399 23681 28408 23715
rect 28356 23672 28408 23681
rect 24952 23604 25004 23656
rect 23480 23536 23532 23588
rect 24032 23536 24084 23588
rect 27804 23536 27856 23588
rect 17500 23468 17552 23520
rect 17776 23468 17828 23520
rect 21272 23468 21324 23520
rect 21364 23468 21416 23520
rect 22928 23468 22980 23520
rect 26240 23468 26292 23520
rect 26608 23468 26660 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 10600 23307 10652 23316
rect 10600 23273 10609 23307
rect 10609 23273 10643 23307
rect 10643 23273 10652 23307
rect 10600 23264 10652 23273
rect 14004 23264 14056 23316
rect 14924 23307 14976 23316
rect 14924 23273 14933 23307
rect 14933 23273 14967 23307
rect 14967 23273 14976 23307
rect 14924 23264 14976 23273
rect 18144 23264 18196 23316
rect 10416 23171 10468 23180
rect 10416 23137 10425 23171
rect 10425 23137 10459 23171
rect 10459 23137 10468 23171
rect 10416 23128 10468 23137
rect 11060 23128 11112 23180
rect 12440 23171 12492 23180
rect 12440 23137 12449 23171
rect 12449 23137 12483 23171
rect 12483 23137 12492 23171
rect 12440 23128 12492 23137
rect 8300 23060 8352 23112
rect 11244 23060 11296 23112
rect 11888 23060 11940 23112
rect 13912 23128 13964 23180
rect 15292 23128 15344 23180
rect 19892 23264 19944 23316
rect 21272 23264 21324 23316
rect 24676 23307 24728 23316
rect 24676 23273 24685 23307
rect 24685 23273 24719 23307
rect 24719 23273 24728 23307
rect 24676 23264 24728 23273
rect 26424 23307 26476 23316
rect 26424 23273 26433 23307
rect 26433 23273 26467 23307
rect 26467 23273 26476 23307
rect 26424 23264 26476 23273
rect 13820 23060 13872 23112
rect 14372 23060 14424 23112
rect 17500 23103 17552 23112
rect 17500 23069 17509 23103
rect 17509 23069 17543 23103
rect 17543 23069 17552 23103
rect 17500 23060 17552 23069
rect 17684 23060 17736 23112
rect 19156 23060 19208 23112
rect 16304 23035 16356 23044
rect 16304 23001 16313 23035
rect 16313 23001 16347 23035
rect 16347 23001 16356 23035
rect 16856 23035 16908 23044
rect 16304 22992 16356 23001
rect 16856 23001 16865 23035
rect 16865 23001 16899 23035
rect 16899 23001 16908 23035
rect 16856 22992 16908 23001
rect 21088 23128 21140 23180
rect 21456 23128 21508 23180
rect 21180 23060 21232 23112
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 21640 23060 21692 23112
rect 24952 23128 25004 23180
rect 19524 23035 19576 23044
rect 12072 22924 12124 22976
rect 14740 22924 14792 22976
rect 15752 22924 15804 22976
rect 16488 22924 16540 22976
rect 19524 23001 19533 23035
rect 19533 23001 19567 23035
rect 19567 23001 19576 23035
rect 19524 22992 19576 23001
rect 17868 22924 17920 22976
rect 18880 22924 18932 22976
rect 19340 22924 19392 22976
rect 19800 22992 19852 23044
rect 21088 22992 21140 23044
rect 23756 23060 23808 23112
rect 24492 23060 24544 23112
rect 26240 23060 26292 23112
rect 23664 23035 23716 23044
rect 23664 23001 23673 23035
rect 23673 23001 23707 23035
rect 23707 23001 23716 23035
rect 23664 22992 23716 23001
rect 28448 23060 28500 23112
rect 20812 22924 20864 22976
rect 23296 22924 23348 22976
rect 25688 22967 25740 22976
rect 25688 22933 25697 22967
rect 25697 22933 25731 22967
rect 25731 22933 25740 22967
rect 25688 22924 25740 22933
rect 25872 22924 25924 22976
rect 27804 22924 27856 22976
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 11888 22763 11940 22772
rect 11888 22729 11897 22763
rect 11897 22729 11931 22763
rect 11931 22729 11940 22763
rect 11888 22720 11940 22729
rect 1860 22652 1912 22704
rect 18696 22720 18748 22772
rect 19432 22720 19484 22772
rect 19800 22720 19852 22772
rect 19892 22720 19944 22772
rect 9128 22516 9180 22568
rect 9772 22584 9824 22636
rect 10968 22584 11020 22636
rect 11796 22627 11848 22636
rect 11796 22593 11805 22627
rect 11805 22593 11839 22627
rect 11839 22593 11848 22627
rect 11796 22584 11848 22593
rect 12348 22584 12400 22636
rect 13084 22627 13136 22636
rect 13084 22593 13093 22627
rect 13093 22593 13127 22627
rect 13127 22593 13136 22627
rect 15476 22652 15528 22704
rect 15752 22695 15804 22704
rect 15752 22661 15761 22695
rect 15761 22661 15795 22695
rect 15795 22661 15804 22695
rect 15752 22652 15804 22661
rect 16856 22652 16908 22704
rect 22744 22652 22796 22704
rect 13084 22584 13136 22593
rect 13728 22584 13780 22636
rect 14740 22584 14792 22636
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17500 22627 17552 22636
rect 17500 22593 17509 22627
rect 17509 22593 17543 22627
rect 17543 22593 17552 22627
rect 17500 22584 17552 22593
rect 17868 22584 17920 22636
rect 11060 22516 11112 22568
rect 12532 22516 12584 22568
rect 14004 22516 14056 22568
rect 11704 22448 11756 22500
rect 13636 22448 13688 22500
rect 14372 22448 14424 22500
rect 18788 22516 18840 22568
rect 19432 22516 19484 22568
rect 20260 22516 20312 22568
rect 20996 22584 21048 22636
rect 22560 22584 22612 22636
rect 22928 22627 22980 22636
rect 22928 22593 22937 22627
rect 22937 22593 22971 22627
rect 22971 22593 22980 22627
rect 22928 22584 22980 22593
rect 21272 22516 21324 22568
rect 25688 22720 25740 22772
rect 23848 22652 23900 22704
rect 25596 22652 25648 22704
rect 23572 22516 23624 22568
rect 19892 22448 19944 22500
rect 20076 22448 20128 22500
rect 21180 22448 21232 22500
rect 8760 22380 8812 22432
rect 10324 22380 10376 22432
rect 10508 22380 10560 22432
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 14740 22380 14792 22432
rect 16764 22380 16816 22432
rect 18880 22380 18932 22432
rect 19524 22380 19576 22432
rect 19616 22380 19668 22432
rect 20904 22380 20956 22432
rect 22192 22380 22244 22432
rect 22744 22380 22796 22432
rect 27896 22584 27948 22636
rect 28264 22491 28316 22500
rect 28264 22457 28273 22491
rect 28273 22457 28307 22491
rect 28307 22457 28316 22491
rect 28264 22448 28316 22457
rect 24676 22380 24728 22432
rect 25688 22380 25740 22432
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 10876 22176 10928 22228
rect 13728 22176 13780 22228
rect 14188 22176 14240 22228
rect 18788 22176 18840 22228
rect 18880 22176 18932 22228
rect 19156 22176 19208 22228
rect 19432 22219 19484 22228
rect 19432 22185 19441 22219
rect 19441 22185 19475 22219
rect 19475 22185 19484 22219
rect 19432 22176 19484 22185
rect 19892 22176 19944 22228
rect 9128 22108 9180 22160
rect 13820 22108 13872 22160
rect 10324 22040 10376 22092
rect 14280 22040 14332 22092
rect 1768 22015 1820 22024
rect 1768 21981 1777 22015
rect 1777 21981 1811 22015
rect 1811 21981 1820 22015
rect 1768 21972 1820 21981
rect 8760 21972 8812 22024
rect 10508 21972 10560 22024
rect 7380 21904 7432 21956
rect 11244 21972 11296 22024
rect 11980 22015 12032 22024
rect 11980 21981 11989 22015
rect 11989 21981 12023 22015
rect 12023 21981 12032 22015
rect 11980 21972 12032 21981
rect 12164 22015 12216 22024
rect 12164 21981 12173 22015
rect 12173 21981 12207 22015
rect 12207 21981 12216 22015
rect 12164 21972 12216 21981
rect 12440 21972 12492 22024
rect 15200 22108 15252 22160
rect 16856 22108 16908 22160
rect 20076 22108 20128 22160
rect 20260 22108 20312 22160
rect 20720 22108 20772 22160
rect 21180 22108 21232 22160
rect 22744 22108 22796 22160
rect 23572 22176 23624 22228
rect 24400 22176 24452 22228
rect 27620 22176 27672 22228
rect 15016 22040 15068 22092
rect 15936 22083 15988 22092
rect 15936 22049 15945 22083
rect 15945 22049 15979 22083
rect 15979 22049 15988 22083
rect 15936 22040 15988 22049
rect 18052 22040 18104 22092
rect 20996 22083 21048 22092
rect 20996 22049 21005 22083
rect 21005 22049 21039 22083
rect 21039 22049 21048 22083
rect 20996 22040 21048 22049
rect 22928 22083 22980 22092
rect 22928 22049 22937 22083
rect 22937 22049 22971 22083
rect 22971 22049 22980 22083
rect 22928 22040 22980 22049
rect 11152 21904 11204 21956
rect 14372 21904 14424 21956
rect 8760 21836 8812 21888
rect 10048 21836 10100 21888
rect 11060 21836 11112 21888
rect 12624 21879 12676 21888
rect 12624 21845 12633 21879
rect 12633 21845 12667 21879
rect 12667 21845 12676 21879
rect 12624 21836 12676 21845
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 15016 21904 15068 21956
rect 13728 21836 13780 21845
rect 14648 21836 14700 21888
rect 16028 21972 16080 22024
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 19524 21972 19576 22024
rect 22560 21972 22612 22024
rect 15384 21947 15436 21956
rect 15384 21913 15393 21947
rect 15393 21913 15427 21947
rect 15427 21913 15436 21947
rect 15384 21904 15436 21913
rect 15568 21904 15620 21956
rect 16488 21836 16540 21888
rect 16580 21836 16632 21888
rect 17776 21904 17828 21956
rect 20812 21904 20864 21956
rect 21364 21904 21416 21956
rect 22376 21947 22428 21956
rect 21088 21836 21140 21888
rect 22376 21913 22385 21947
rect 22385 21913 22419 21947
rect 22419 21913 22428 21947
rect 22376 21904 22428 21913
rect 23388 21904 23440 21956
rect 24124 21972 24176 22024
rect 27712 22040 27764 22092
rect 25596 21972 25648 22024
rect 26240 22015 26292 22024
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 24216 21904 24268 21956
rect 25320 21947 25372 21956
rect 25320 21913 25329 21947
rect 25329 21913 25363 21947
rect 25363 21913 25372 21947
rect 25320 21904 25372 21913
rect 26516 21947 26568 21956
rect 26516 21913 26525 21947
rect 26525 21913 26559 21947
rect 26559 21913 26568 21947
rect 26516 21904 26568 21913
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 25044 21836 25096 21888
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 7380 21675 7432 21684
rect 7380 21641 7389 21675
rect 7389 21641 7423 21675
rect 7423 21641 7432 21675
rect 7380 21632 7432 21641
rect 7288 21539 7340 21548
rect 7288 21505 7297 21539
rect 7297 21505 7331 21539
rect 7331 21505 7340 21539
rect 7288 21496 7340 21505
rect 9956 21496 10008 21548
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 12716 21632 12768 21684
rect 14372 21632 14424 21684
rect 20260 21632 20312 21684
rect 20720 21632 20772 21684
rect 12624 21564 12676 21616
rect 15752 21607 15804 21616
rect 13544 21496 13596 21548
rect 13820 21539 13872 21548
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 14464 21496 14516 21548
rect 15016 21496 15068 21548
rect 12440 21471 12492 21480
rect 12440 21437 12449 21471
rect 12449 21437 12483 21471
rect 12483 21437 12492 21471
rect 12440 21428 12492 21437
rect 15108 21471 15160 21480
rect 15108 21437 15117 21471
rect 15117 21437 15151 21471
rect 15151 21437 15160 21471
rect 15108 21428 15160 21437
rect 15752 21573 15761 21607
rect 15761 21573 15795 21607
rect 15795 21573 15804 21607
rect 15752 21564 15804 21573
rect 17776 21564 17828 21616
rect 18512 21564 18564 21616
rect 22192 21564 22244 21616
rect 24676 21632 24728 21684
rect 24860 21632 24912 21684
rect 23020 21607 23072 21616
rect 20076 21496 20128 21548
rect 22560 21496 22612 21548
rect 23020 21573 23029 21607
rect 23029 21573 23063 21607
rect 23063 21573 23072 21607
rect 23020 21564 23072 21573
rect 23480 21564 23532 21616
rect 24492 21564 24544 21616
rect 24584 21564 24636 21616
rect 17684 21428 17736 21480
rect 17776 21428 17828 21480
rect 17960 21471 18012 21480
rect 17960 21437 17969 21471
rect 17969 21437 18003 21471
rect 18003 21437 18012 21471
rect 17960 21428 18012 21437
rect 18236 21471 18288 21480
rect 18236 21437 18245 21471
rect 18245 21437 18279 21471
rect 18279 21437 18288 21471
rect 18236 21428 18288 21437
rect 18972 21428 19024 21480
rect 19248 21428 19300 21480
rect 23388 21428 23440 21480
rect 23572 21428 23624 21480
rect 24492 21471 24544 21480
rect 24492 21437 24501 21471
rect 24501 21437 24535 21471
rect 24535 21437 24544 21471
rect 24492 21428 24544 21437
rect 24676 21496 24728 21548
rect 26240 21496 26292 21548
rect 27160 21539 27212 21548
rect 24768 21428 24820 21480
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 28172 21428 28224 21480
rect 19616 21360 19668 21412
rect 10324 21335 10376 21344
rect 10324 21301 10333 21335
rect 10333 21301 10367 21335
rect 10367 21301 10376 21335
rect 10324 21292 10376 21301
rect 11888 21292 11940 21344
rect 12256 21292 12308 21344
rect 12440 21292 12492 21344
rect 15660 21292 15712 21344
rect 17868 21292 17920 21344
rect 19708 21335 19760 21344
rect 19708 21301 19717 21335
rect 19717 21301 19751 21335
rect 19751 21301 19760 21335
rect 19708 21292 19760 21301
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 22284 21292 22336 21344
rect 24216 21360 24268 21412
rect 25780 21360 25832 21412
rect 24032 21292 24084 21344
rect 28080 21292 28132 21344
rect 28264 21335 28316 21344
rect 28264 21301 28273 21335
rect 28273 21301 28307 21335
rect 28307 21301 28316 21335
rect 28264 21292 28316 21301
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 12164 21088 12216 21140
rect 15752 21088 15804 21140
rect 16580 21088 16632 21140
rect 17040 21088 17092 21140
rect 13360 21020 13412 21072
rect 10324 20952 10376 21004
rect 15200 21020 15252 21072
rect 19616 21088 19668 21140
rect 20168 21088 20220 21140
rect 20628 21088 20680 21140
rect 23112 21131 23164 21140
rect 23112 21097 23121 21131
rect 23121 21097 23155 21131
rect 23155 21097 23164 21131
rect 23112 21088 23164 21097
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 6092 20927 6144 20936
rect 6092 20893 6101 20927
rect 6101 20893 6135 20927
rect 6135 20893 6144 20927
rect 6092 20884 6144 20893
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 11152 20884 11204 20936
rect 11888 20884 11940 20936
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 12532 20884 12584 20936
rect 14648 20884 14700 20936
rect 19248 20952 19300 21004
rect 24124 21088 24176 21140
rect 18696 20884 18748 20936
rect 19340 20884 19392 20936
rect 19524 20884 19576 20936
rect 21824 20952 21876 21004
rect 22836 20952 22888 21004
rect 24768 20952 24820 21004
rect 26240 20952 26292 21004
rect 24032 20884 24084 20936
rect 3976 20748 4028 20800
rect 6184 20791 6236 20800
rect 6184 20757 6193 20791
rect 6193 20757 6227 20791
rect 6227 20757 6236 20791
rect 6184 20748 6236 20757
rect 9864 20748 9916 20800
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 10508 20748 10560 20800
rect 15568 20816 15620 20868
rect 16672 20859 16724 20868
rect 16672 20825 16681 20859
rect 16681 20825 16715 20859
rect 16715 20825 16724 20859
rect 16672 20816 16724 20825
rect 16764 20859 16816 20868
rect 16764 20825 16773 20859
rect 16773 20825 16807 20859
rect 16807 20825 16816 20859
rect 16764 20816 16816 20825
rect 12808 20748 12860 20800
rect 15200 20748 15252 20800
rect 15384 20748 15436 20800
rect 19156 20748 19208 20800
rect 21088 20816 21140 20868
rect 22836 20748 22888 20800
rect 27620 20816 27672 20868
rect 28264 20816 28316 20868
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 10508 20587 10560 20596
rect 10508 20553 10517 20587
rect 10517 20553 10551 20587
rect 10551 20553 10560 20587
rect 10508 20544 10560 20553
rect 10968 20544 11020 20596
rect 12992 20544 13044 20596
rect 18144 20544 18196 20596
rect 18236 20544 18288 20596
rect 21364 20544 21416 20596
rect 21640 20544 21692 20596
rect 22468 20544 22520 20596
rect 26424 20544 26476 20596
rect 27896 20587 27948 20596
rect 27896 20553 27905 20587
rect 27905 20553 27939 20587
rect 27939 20553 27948 20587
rect 27896 20544 27948 20553
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 10048 20451 10100 20460
rect 10048 20417 10057 20451
rect 10057 20417 10091 20451
rect 10091 20417 10100 20451
rect 10048 20408 10100 20417
rect 10968 20408 11020 20460
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 15660 20408 15712 20460
rect 17132 20408 17184 20460
rect 17500 20408 17552 20460
rect 6092 20340 6144 20392
rect 11060 20340 11112 20392
rect 13452 20383 13504 20392
rect 13452 20349 13461 20383
rect 13461 20349 13495 20383
rect 13495 20349 13504 20383
rect 13452 20340 13504 20349
rect 13544 20340 13596 20392
rect 14740 20383 14792 20392
rect 14740 20349 14749 20383
rect 14749 20349 14783 20383
rect 14783 20349 14792 20383
rect 14740 20340 14792 20349
rect 19708 20476 19760 20528
rect 17960 20408 18012 20460
rect 19432 20408 19484 20460
rect 19616 20408 19668 20460
rect 5080 20272 5132 20324
rect 15200 20272 15252 20324
rect 19432 20272 19484 20324
rect 20076 20272 20128 20324
rect 5724 20204 5776 20256
rect 7748 20204 7800 20256
rect 11704 20204 11756 20256
rect 12440 20204 12492 20256
rect 14372 20204 14424 20256
rect 16764 20204 16816 20256
rect 19064 20204 19116 20256
rect 19340 20204 19392 20256
rect 20444 20383 20496 20392
rect 20444 20349 20453 20383
rect 20453 20349 20487 20383
rect 20487 20349 20496 20383
rect 20444 20340 20496 20349
rect 23480 20476 23532 20528
rect 21640 20408 21692 20460
rect 28080 20451 28132 20460
rect 22008 20340 22060 20392
rect 28080 20417 28089 20451
rect 28089 20417 28123 20451
rect 28123 20417 28132 20451
rect 28080 20408 28132 20417
rect 23112 20272 23164 20324
rect 20720 20204 20772 20256
rect 21364 20204 21416 20256
rect 23020 20204 23072 20256
rect 23572 20340 23624 20392
rect 25044 20340 25096 20392
rect 24676 20204 24728 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 5080 20043 5132 20052
rect 5080 20009 5089 20043
rect 5089 20009 5123 20043
rect 5123 20009 5132 20043
rect 5080 20000 5132 20009
rect 6092 20000 6144 20052
rect 12164 20000 12216 20052
rect 14740 20000 14792 20052
rect 16120 20000 16172 20052
rect 17776 20000 17828 20052
rect 17960 20000 18012 20052
rect 18420 20000 18472 20052
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 4068 19796 4120 19848
rect 6736 19796 6788 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 10784 19796 10836 19848
rect 11980 19796 12032 19848
rect 14096 19796 14148 19848
rect 18236 19932 18288 19984
rect 22192 20000 22244 20052
rect 16856 19864 16908 19916
rect 21548 19932 21600 19984
rect 23112 20000 23164 20052
rect 25964 20000 26016 20052
rect 28172 20043 28224 20052
rect 28172 20009 28181 20043
rect 28181 20009 28215 20043
rect 28215 20009 28224 20043
rect 28172 20000 28224 20009
rect 16028 19796 16080 19848
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 18144 19796 18196 19848
rect 18604 19864 18656 19916
rect 19248 19864 19300 19916
rect 21640 19864 21692 19916
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 24676 19907 24728 19916
rect 24676 19873 24685 19907
rect 24685 19873 24719 19907
rect 24719 19873 24728 19907
rect 24676 19864 24728 19873
rect 26056 19932 26108 19984
rect 18696 19796 18748 19848
rect 19432 19796 19484 19848
rect 21272 19796 21324 19848
rect 28356 19839 28408 19848
rect 28356 19805 28365 19839
rect 28365 19805 28399 19839
rect 28399 19805 28408 19839
rect 28356 19796 28408 19805
rect 13268 19728 13320 19780
rect 3700 19660 3752 19712
rect 9220 19703 9272 19712
rect 9220 19669 9229 19703
rect 9229 19669 9263 19703
rect 9263 19669 9272 19703
rect 9220 19660 9272 19669
rect 10508 19660 10560 19712
rect 11152 19660 11204 19712
rect 12624 19660 12676 19712
rect 13544 19703 13596 19712
rect 13544 19669 13553 19703
rect 13553 19669 13587 19703
rect 13587 19669 13596 19703
rect 13544 19660 13596 19669
rect 15660 19660 15712 19712
rect 16764 19771 16816 19780
rect 16764 19737 16773 19771
rect 16773 19737 16807 19771
rect 16807 19737 16816 19771
rect 16764 19728 16816 19737
rect 17500 19660 17552 19712
rect 18052 19660 18104 19712
rect 18696 19660 18748 19712
rect 19616 19660 19668 19712
rect 19892 19728 19944 19780
rect 21916 19728 21968 19780
rect 22468 19728 22520 19780
rect 23296 19728 23348 19780
rect 21364 19660 21416 19712
rect 24492 19728 24544 19780
rect 26700 19771 26752 19780
rect 26700 19737 26709 19771
rect 26709 19737 26743 19771
rect 26743 19737 26752 19771
rect 26700 19728 26752 19737
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 10968 19499 11020 19508
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 11980 19499 12032 19508
rect 11980 19465 11989 19499
rect 11989 19465 12023 19499
rect 12023 19465 12032 19499
rect 11980 19456 12032 19465
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 14556 19456 14608 19508
rect 16028 19499 16080 19508
rect 16028 19465 16037 19499
rect 16037 19465 16071 19499
rect 16071 19465 16080 19499
rect 16028 19456 16080 19465
rect 22468 19456 22520 19508
rect 23020 19456 23072 19508
rect 26424 19456 26476 19508
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 11060 19388 11112 19440
rect 9956 19320 10008 19372
rect 10508 19363 10560 19372
rect 10508 19329 10517 19363
rect 10517 19329 10551 19363
rect 10551 19329 10560 19363
rect 10508 19320 10560 19329
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 13360 19388 13412 19440
rect 18696 19388 18748 19440
rect 20996 19388 21048 19440
rect 21548 19388 21600 19440
rect 25136 19388 25188 19440
rect 12164 19184 12216 19236
rect 7380 19159 7432 19168
rect 7380 19125 7389 19159
rect 7389 19125 7423 19159
rect 7423 19125 7432 19159
rect 7380 19116 7432 19125
rect 9864 19116 9916 19168
rect 11704 19116 11756 19168
rect 13544 19320 13596 19372
rect 13636 19252 13688 19304
rect 13912 19295 13964 19304
rect 13912 19261 13921 19295
rect 13921 19261 13955 19295
rect 13955 19261 13964 19295
rect 13912 19252 13964 19261
rect 17408 19320 17460 19372
rect 17592 19320 17644 19372
rect 17960 19320 18012 19372
rect 20812 19320 20864 19372
rect 21456 19320 21508 19372
rect 21640 19320 21692 19372
rect 23756 19320 23808 19372
rect 24676 19320 24728 19372
rect 16948 19252 17000 19304
rect 19984 19252 20036 19304
rect 23204 19252 23256 19304
rect 23296 19252 23348 19304
rect 25044 19295 25096 19304
rect 25044 19261 25053 19295
rect 25053 19261 25087 19295
rect 25087 19261 25096 19295
rect 25044 19252 25096 19261
rect 16304 19116 16356 19168
rect 19892 19159 19944 19168
rect 19892 19125 19901 19159
rect 19901 19125 19935 19159
rect 19935 19125 19944 19159
rect 19892 19116 19944 19125
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 20720 19116 20772 19168
rect 22836 19116 22888 19168
rect 23204 19116 23256 19168
rect 27620 19184 27672 19236
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 10416 18912 10468 18964
rect 22836 18955 22888 18964
rect 6736 18844 6788 18896
rect 6828 18708 6880 18760
rect 17960 18844 18012 18896
rect 19064 18844 19116 18896
rect 22836 18921 22845 18955
rect 22845 18921 22879 18955
rect 22879 18921 22888 18955
rect 22836 18912 22888 18921
rect 26240 18912 26292 18964
rect 27988 18912 28040 18964
rect 9220 18776 9272 18828
rect 10324 18776 10376 18828
rect 13268 18776 13320 18828
rect 14372 18776 14424 18828
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 11888 18708 11940 18760
rect 14556 18708 14608 18760
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 18972 18776 19024 18828
rect 19248 18776 19300 18828
rect 23388 18844 23440 18896
rect 24584 18819 24636 18828
rect 15476 18708 15528 18717
rect 7104 18640 7156 18692
rect 13636 18640 13688 18692
rect 15568 18640 15620 18692
rect 16212 18708 16264 18760
rect 1768 18615 1820 18624
rect 1768 18581 1777 18615
rect 1777 18581 1811 18615
rect 1811 18581 1820 18615
rect 1768 18572 1820 18581
rect 8300 18572 8352 18624
rect 12256 18572 12308 18624
rect 14464 18572 14516 18624
rect 16212 18572 16264 18624
rect 17408 18572 17460 18624
rect 18144 18708 18196 18760
rect 18420 18708 18472 18760
rect 20904 18708 20956 18760
rect 17868 18640 17920 18692
rect 19892 18640 19944 18692
rect 21272 18640 21324 18692
rect 22836 18640 22888 18692
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 26516 18844 26568 18896
rect 27068 18844 27120 18896
rect 29920 18708 29972 18760
rect 18328 18572 18380 18624
rect 23112 18572 23164 18624
rect 24216 18640 24268 18692
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 8300 18411 8352 18420
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 12164 18368 12216 18420
rect 6736 18300 6788 18352
rect 7380 18232 7432 18284
rect 8392 18232 8444 18284
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 10876 18232 10928 18284
rect 11888 18232 11940 18284
rect 12256 18275 12308 18284
rect 12256 18241 12265 18275
rect 12265 18241 12299 18275
rect 12299 18241 12308 18275
rect 12256 18232 12308 18241
rect 13912 18368 13964 18420
rect 15568 18368 15620 18420
rect 14464 18343 14516 18352
rect 14464 18309 14473 18343
rect 14473 18309 14507 18343
rect 14507 18309 14516 18343
rect 14464 18300 14516 18309
rect 14556 18300 14608 18352
rect 19524 18368 19576 18420
rect 19984 18411 20036 18420
rect 19984 18377 19993 18411
rect 19993 18377 20027 18411
rect 20027 18377 20036 18411
rect 19984 18368 20036 18377
rect 20444 18368 20496 18420
rect 23204 18368 23256 18420
rect 23572 18368 23624 18420
rect 25136 18368 25188 18420
rect 16948 18343 17000 18352
rect 16948 18309 16957 18343
rect 16957 18309 16991 18343
rect 16991 18309 17000 18343
rect 16948 18300 17000 18309
rect 17040 18343 17092 18352
rect 17040 18309 17049 18343
rect 17049 18309 17083 18343
rect 17083 18309 17092 18343
rect 17040 18300 17092 18309
rect 17408 18300 17460 18352
rect 19892 18300 19944 18352
rect 25872 18300 25924 18352
rect 7472 18164 7524 18216
rect 8576 18164 8628 18216
rect 11060 18164 11112 18216
rect 9864 18096 9916 18148
rect 11888 18096 11940 18148
rect 13912 18232 13964 18284
rect 15476 18232 15528 18284
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 15936 18232 15988 18284
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16304 18232 16356 18284
rect 14372 18207 14424 18216
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 17224 18207 17276 18216
rect 5540 18028 5592 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 11980 18028 12032 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 18052 18164 18104 18216
rect 18880 18164 18932 18216
rect 23296 18096 23348 18148
rect 19616 18028 19668 18080
rect 23572 18028 23624 18080
rect 23940 18164 23992 18216
rect 24584 18028 24636 18080
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 6828 17824 6880 17876
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 9312 17867 9364 17876
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 9404 17824 9456 17876
rect 5356 17484 5408 17536
rect 8392 17620 8444 17672
rect 9404 17688 9456 17740
rect 9680 17688 9732 17740
rect 13636 17824 13688 17876
rect 24308 17824 24360 17876
rect 24400 17824 24452 17876
rect 15200 17799 15252 17808
rect 15200 17765 15209 17799
rect 15209 17765 15243 17799
rect 15243 17765 15252 17799
rect 15200 17756 15252 17765
rect 17040 17756 17092 17808
rect 17960 17756 18012 17808
rect 15844 17688 15896 17740
rect 9220 17663 9272 17672
rect 9220 17629 9229 17663
rect 9229 17629 9263 17663
rect 9263 17629 9272 17663
rect 9220 17620 9272 17629
rect 11244 17620 11296 17672
rect 11980 17663 12032 17672
rect 11060 17552 11112 17604
rect 10968 17484 11020 17536
rect 11152 17527 11204 17536
rect 11152 17493 11161 17527
rect 11161 17493 11195 17527
rect 11195 17493 11204 17527
rect 11152 17484 11204 17493
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 12348 17620 12400 17672
rect 12900 17620 12952 17672
rect 13728 17663 13780 17672
rect 12992 17552 13044 17604
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14280 17620 14332 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 17592 17620 17644 17672
rect 18052 17688 18104 17740
rect 18696 17688 18748 17740
rect 21640 17731 21692 17740
rect 21640 17697 21649 17731
rect 21649 17697 21683 17731
rect 21683 17697 21692 17731
rect 21640 17688 21692 17697
rect 24952 17756 25004 17808
rect 24492 17688 24544 17740
rect 24584 17688 24636 17740
rect 27896 17688 27948 17740
rect 11980 17484 12032 17536
rect 17960 17552 18012 17604
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 18236 17620 18288 17672
rect 18788 17484 18840 17536
rect 19892 17484 19944 17536
rect 20628 17484 20680 17536
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 21548 17552 21600 17604
rect 22008 17552 22060 17604
rect 22376 17552 22428 17604
rect 23572 17552 23624 17604
rect 26240 17552 26292 17604
rect 23388 17527 23440 17536
rect 23388 17493 23397 17527
rect 23397 17493 23431 17527
rect 23431 17493 23440 17527
rect 23388 17484 23440 17493
rect 24308 17484 24360 17536
rect 28172 17484 28224 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 6920 17280 6972 17332
rect 8300 17212 8352 17264
rect 11796 17280 11848 17332
rect 12348 17323 12400 17332
rect 12348 17289 12357 17323
rect 12357 17289 12391 17323
rect 12391 17289 12400 17323
rect 12348 17280 12400 17289
rect 13360 17280 13412 17332
rect 5172 17144 5224 17196
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 7196 17144 7248 17196
rect 11152 17187 11204 17196
rect 11152 17153 11161 17187
rect 11161 17153 11195 17187
rect 11195 17153 11204 17187
rect 11152 17144 11204 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 13452 17212 13504 17264
rect 14188 17212 14240 17264
rect 16028 17280 16080 17332
rect 17132 17212 17184 17264
rect 17592 17280 17644 17332
rect 18604 17212 18656 17264
rect 20168 17280 20220 17332
rect 20628 17280 20680 17332
rect 20720 17280 20772 17332
rect 21364 17280 21416 17332
rect 21456 17280 21508 17332
rect 21824 17280 21876 17332
rect 25136 17212 25188 17264
rect 7472 17076 7524 17128
rect 1768 17051 1820 17060
rect 1768 17017 1777 17051
rect 1777 17017 1811 17051
rect 1811 17017 1820 17051
rect 1768 17008 1820 17017
rect 5724 17051 5776 17060
rect 5724 17017 5733 17051
rect 5733 17017 5767 17051
rect 5767 17017 5776 17051
rect 5724 17008 5776 17017
rect 8024 17076 8076 17128
rect 12624 17076 12676 17128
rect 16580 17144 16632 17196
rect 17408 17144 17460 17196
rect 18052 17187 18104 17196
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 13360 17119 13412 17128
rect 11244 17008 11296 17060
rect 12992 17008 13044 17060
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 14556 17008 14608 17060
rect 14740 17008 14792 17060
rect 17868 17076 17920 17128
rect 20812 17144 20864 17196
rect 21088 17144 21140 17196
rect 21640 17144 21692 17196
rect 24584 17144 24636 17196
rect 28356 17187 28408 17196
rect 28356 17153 28365 17187
rect 28365 17153 28399 17187
rect 28399 17153 28408 17187
rect 28356 17144 28408 17153
rect 22284 17076 22336 17128
rect 22468 17076 22520 17128
rect 24124 17076 24176 17128
rect 24492 17076 24544 17128
rect 26700 17076 26752 17128
rect 21916 17008 21968 17060
rect 22008 17008 22060 17060
rect 19708 16940 19760 16992
rect 19892 16940 19944 16992
rect 22560 16940 22612 16992
rect 24032 16940 24084 16992
rect 27988 16940 28040 16992
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 5172 16736 5224 16788
rect 7196 16736 7248 16788
rect 3976 16668 4028 16720
rect 7012 16668 7064 16720
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 8024 16532 8076 16584
rect 12532 16736 12584 16788
rect 12624 16736 12676 16788
rect 21456 16736 21508 16788
rect 8576 16668 8628 16720
rect 11704 16668 11756 16720
rect 9864 16643 9916 16652
rect 9864 16609 9873 16643
rect 9873 16609 9907 16643
rect 9907 16609 9916 16643
rect 9864 16600 9916 16609
rect 12440 16600 12492 16652
rect 14556 16668 14608 16720
rect 18972 16668 19024 16720
rect 19340 16668 19392 16720
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 15384 16600 15436 16652
rect 15844 16600 15896 16652
rect 15936 16600 15988 16652
rect 16304 16600 16356 16652
rect 11244 16532 11296 16584
rect 12072 16464 12124 16516
rect 6920 16396 6972 16448
rect 10968 16396 11020 16448
rect 12440 16396 12492 16448
rect 17132 16532 17184 16584
rect 17592 16532 17644 16584
rect 17960 16532 18012 16584
rect 18144 16532 18196 16584
rect 19248 16600 19300 16652
rect 20720 16668 20772 16720
rect 23388 16736 23440 16788
rect 20076 16600 20128 16652
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 21916 16600 21968 16652
rect 22468 16600 22520 16652
rect 22560 16600 22612 16652
rect 23756 16600 23808 16652
rect 24584 16600 24636 16652
rect 26608 16643 26660 16652
rect 26608 16609 26617 16643
rect 26617 16609 26651 16643
rect 26651 16609 26660 16643
rect 26608 16600 26660 16609
rect 19616 16464 19668 16516
rect 21272 16464 21324 16516
rect 21640 16464 21692 16516
rect 21824 16464 21876 16516
rect 22376 16464 22428 16516
rect 23204 16464 23256 16516
rect 25136 16464 25188 16516
rect 27620 16464 27672 16516
rect 28080 16464 28132 16516
rect 16120 16396 16172 16448
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 17132 16439 17184 16448
rect 16212 16396 16264 16405
rect 17132 16405 17141 16439
rect 17141 16405 17175 16439
rect 17175 16405 17184 16439
rect 17132 16396 17184 16405
rect 17776 16439 17828 16448
rect 17776 16405 17785 16439
rect 17785 16405 17819 16439
rect 17819 16405 17828 16439
rect 17776 16396 17828 16405
rect 20352 16396 20404 16448
rect 20444 16396 20496 16448
rect 21548 16396 21600 16448
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 7104 16192 7156 16244
rect 9772 16192 9824 16244
rect 12072 16192 12124 16244
rect 12440 16192 12492 16244
rect 13452 16192 13504 16244
rect 14188 16235 14240 16244
rect 14188 16201 14197 16235
rect 14197 16201 14231 16235
rect 14231 16201 14240 16235
rect 14188 16192 14240 16201
rect 14740 16192 14792 16244
rect 10600 16124 10652 16176
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 3700 16056 3752 16108
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 9036 16099 9088 16108
rect 9036 16065 9045 16099
rect 9045 16065 9079 16099
rect 9079 16065 9088 16099
rect 9036 16056 9088 16065
rect 9312 16056 9364 16108
rect 11244 16056 11296 16108
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 9220 15988 9272 16040
rect 9772 15988 9824 16040
rect 10232 15920 10284 15972
rect 10508 16031 10560 16040
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 13636 16124 13688 16176
rect 17132 16192 17184 16244
rect 21916 16192 21968 16244
rect 17500 16167 17552 16176
rect 12716 16056 12768 16108
rect 13176 16056 13228 16108
rect 15476 16056 15528 16108
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 10508 15988 10560 15997
rect 6552 15852 6604 15904
rect 11060 15920 11112 15972
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 17500 16133 17509 16167
rect 17509 16133 17543 16167
rect 17543 16133 17552 16167
rect 17500 16124 17552 16133
rect 17868 16056 17920 16108
rect 19248 16124 19300 16176
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 20996 16056 21048 16108
rect 21088 16056 21140 16108
rect 22468 16124 22520 16176
rect 24492 16192 24544 16244
rect 24584 16124 24636 16176
rect 25136 16124 25188 16176
rect 18972 16031 19024 16040
rect 15660 15920 15712 15972
rect 10968 15895 11020 15904
rect 10968 15861 10977 15895
rect 10977 15861 11011 15895
rect 11011 15861 11020 15895
rect 13544 15895 13596 15904
rect 10968 15852 11020 15861
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 19524 15988 19576 16040
rect 20260 15988 20312 16040
rect 21732 15920 21784 15972
rect 22100 15988 22152 16040
rect 28540 16056 28592 16108
rect 22468 16031 22520 16040
rect 22468 15997 22477 16031
rect 22477 15997 22511 16031
rect 22511 15997 22520 16031
rect 22468 15988 22520 15997
rect 22560 15988 22612 16040
rect 24032 15988 24084 16040
rect 26424 16031 26476 16040
rect 26424 15997 26433 16031
rect 26433 15997 26467 16031
rect 26467 15997 26476 16031
rect 26424 15988 26476 15997
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 21640 15852 21692 15904
rect 22192 15852 22244 15904
rect 23940 15895 23992 15904
rect 23940 15861 23949 15895
rect 23949 15861 23983 15895
rect 23983 15861 23992 15895
rect 23940 15852 23992 15861
rect 24768 15852 24820 15904
rect 26700 15852 26752 15904
rect 28264 15895 28316 15904
rect 28264 15861 28273 15895
rect 28273 15861 28307 15895
rect 28307 15861 28316 15895
rect 28264 15852 28316 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 9956 15648 10008 15700
rect 11152 15648 11204 15700
rect 11244 15648 11296 15700
rect 21548 15648 21600 15700
rect 7748 15580 7800 15632
rect 6184 15512 6236 15564
rect 7748 15444 7800 15496
rect 9312 15444 9364 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 8392 15376 8444 15428
rect 9036 15376 9088 15428
rect 8300 15308 8352 15360
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 16948 15580 17000 15632
rect 22100 15648 22152 15700
rect 22284 15648 22336 15700
rect 24216 15648 24268 15700
rect 26332 15648 26384 15700
rect 13544 15512 13596 15564
rect 18236 15512 18288 15564
rect 18696 15512 18748 15564
rect 19248 15512 19300 15564
rect 23020 15580 23072 15632
rect 24584 15580 24636 15632
rect 22928 15512 22980 15564
rect 11152 15444 11204 15496
rect 12716 15444 12768 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 15844 15444 15896 15496
rect 12164 15308 12216 15360
rect 13360 15376 13412 15428
rect 13268 15308 13320 15360
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 14740 15419 14792 15428
rect 14740 15385 14749 15419
rect 14749 15385 14783 15419
rect 14783 15385 14792 15419
rect 14740 15376 14792 15385
rect 15200 15308 15252 15360
rect 15384 15376 15436 15428
rect 17592 15444 17644 15496
rect 17868 15444 17920 15496
rect 18144 15444 18196 15496
rect 18788 15444 18840 15496
rect 16304 15376 16356 15428
rect 16396 15376 16448 15428
rect 19340 15376 19392 15428
rect 19616 15376 19668 15428
rect 20720 15376 20772 15428
rect 16580 15308 16632 15360
rect 18604 15308 18656 15360
rect 21824 15376 21876 15428
rect 21916 15419 21968 15428
rect 21916 15385 21925 15419
rect 21925 15385 21959 15419
rect 21959 15385 21968 15419
rect 21916 15376 21968 15385
rect 22376 15376 22428 15428
rect 27712 15512 27764 15564
rect 21548 15308 21600 15360
rect 21732 15308 21784 15360
rect 25872 15376 25924 15428
rect 27804 15376 27856 15428
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 7748 15104 7800 15156
rect 10876 15147 10928 15156
rect 10876 15113 10885 15147
rect 10885 15113 10919 15147
rect 10919 15113 10928 15147
rect 10876 15104 10928 15113
rect 11152 15104 11204 15156
rect 9312 14968 9364 15020
rect 12256 15036 12308 15088
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 12992 14968 13044 15020
rect 13452 15104 13504 15156
rect 17040 15104 17092 15156
rect 16488 15036 16540 15088
rect 18604 15036 18656 15088
rect 20444 15104 20496 15156
rect 20352 15036 20404 15088
rect 22376 15104 22428 15156
rect 22836 15104 22888 15156
rect 23480 15104 23532 15156
rect 25044 15104 25096 15156
rect 23112 15036 23164 15088
rect 15936 15011 15988 15020
rect 9680 14832 9732 14884
rect 12440 14900 12492 14952
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 18236 15011 18288 15020
rect 14464 14900 14516 14952
rect 14832 14900 14884 14952
rect 16856 14900 16908 14952
rect 13452 14832 13504 14884
rect 10140 14764 10192 14816
rect 12440 14764 12492 14816
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 14556 14832 14608 14884
rect 16488 14764 16540 14816
rect 16672 14764 16724 14816
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 20076 14968 20128 15020
rect 20628 14968 20680 15020
rect 21364 14968 21416 15020
rect 18144 14900 18196 14952
rect 19064 14900 19116 14952
rect 22192 14968 22244 15020
rect 24952 15036 25004 15088
rect 27160 15011 27212 15020
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 27988 15011 28040 15020
rect 27988 14977 27997 15011
rect 27997 14977 28031 15011
rect 28031 14977 28040 15011
rect 27988 14968 28040 14977
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24860 14943 24912 14952
rect 24860 14909 24869 14943
rect 24869 14909 24903 14943
rect 24903 14909 24912 14943
rect 24860 14900 24912 14909
rect 26608 14943 26660 14952
rect 26608 14909 26617 14943
rect 26617 14909 26651 14943
rect 26651 14909 26660 14943
rect 26608 14900 26660 14909
rect 19616 14832 19668 14884
rect 22284 14832 22336 14884
rect 20168 14764 20220 14816
rect 20536 14764 20588 14816
rect 24860 14764 24912 14816
rect 26240 14764 26292 14816
rect 27620 14764 27672 14816
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 8392 14560 8444 14612
rect 9956 14560 10008 14612
rect 10508 14560 10560 14612
rect 10140 14424 10192 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 5816 14356 5868 14408
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 11980 14356 12032 14408
rect 13452 14424 13504 14476
rect 16672 14560 16724 14612
rect 15660 14492 15712 14544
rect 21180 14560 21232 14612
rect 23572 14603 23624 14612
rect 23572 14569 23581 14603
rect 23581 14569 23615 14603
rect 23615 14569 23624 14603
rect 23572 14560 23624 14569
rect 17592 14492 17644 14544
rect 8760 14288 8812 14340
rect 14188 14356 14240 14408
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 14832 14356 14884 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 15844 14356 15896 14408
rect 16856 14424 16908 14476
rect 17224 14424 17276 14476
rect 17316 14424 17368 14476
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 19248 14424 19300 14476
rect 22652 14492 22704 14544
rect 26792 14560 26844 14612
rect 28448 14560 28500 14612
rect 24952 14424 25004 14476
rect 26056 14424 26108 14476
rect 17408 14356 17460 14408
rect 17684 14356 17736 14408
rect 18788 14356 18840 14408
rect 19340 14356 19392 14408
rect 19616 14356 19668 14408
rect 16488 14331 16540 14340
rect 16488 14297 16497 14331
rect 16497 14297 16531 14331
rect 16531 14297 16540 14331
rect 16488 14288 16540 14297
rect 4896 14220 4948 14272
rect 10232 14263 10284 14272
rect 10232 14229 10241 14263
rect 10241 14229 10275 14263
rect 10275 14229 10284 14263
rect 10232 14220 10284 14229
rect 14280 14220 14332 14272
rect 15844 14220 15896 14272
rect 17408 14220 17460 14272
rect 17868 14220 17920 14272
rect 23480 14399 23532 14408
rect 23480 14365 23489 14399
rect 23489 14365 23523 14399
rect 23523 14365 23532 14399
rect 23480 14356 23532 14365
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 28356 14399 28408 14408
rect 28356 14365 28365 14399
rect 28365 14365 28399 14399
rect 28399 14365 28408 14399
rect 28356 14356 28408 14365
rect 20352 14288 20404 14340
rect 21180 14288 21232 14340
rect 21456 14331 21508 14340
rect 21456 14297 21465 14331
rect 21465 14297 21499 14331
rect 21499 14297 21508 14331
rect 21456 14288 21508 14297
rect 24768 14288 24820 14340
rect 25136 14288 25188 14340
rect 26148 14288 26200 14340
rect 20536 14220 20588 14272
rect 20628 14220 20680 14272
rect 22836 14220 22888 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 3240 14016 3292 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 10600 13948 10652 14000
rect 11796 13948 11848 14000
rect 13084 14016 13136 14068
rect 14556 14016 14608 14068
rect 15292 14016 15344 14068
rect 16580 14016 16632 14068
rect 12072 13948 12124 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 4896 13923 4948 13932
rect 4896 13889 4905 13923
rect 4905 13889 4939 13923
rect 4939 13889 4948 13923
rect 4896 13880 4948 13889
rect 6368 13880 6420 13932
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 10232 13880 10284 13932
rect 13636 13948 13688 14000
rect 4160 13812 4212 13864
rect 6460 13812 6512 13864
rect 8484 13812 8536 13864
rect 9496 13812 9548 13864
rect 12808 13812 12860 13864
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 14280 13880 14332 13932
rect 14556 13812 14608 13864
rect 15200 13948 15252 14000
rect 17960 14016 18012 14068
rect 18696 14016 18748 14068
rect 18328 13948 18380 14000
rect 19432 13948 19484 14000
rect 20628 14016 20680 14068
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 20904 13948 20956 14000
rect 24032 14016 24084 14068
rect 21088 13880 21140 13932
rect 21272 13880 21324 13932
rect 16948 13855 17000 13864
rect 13176 13744 13228 13796
rect 13636 13744 13688 13796
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17040 13744 17092 13796
rect 17776 13744 17828 13796
rect 18512 13812 18564 13864
rect 18788 13812 18840 13864
rect 20720 13812 20772 13864
rect 24492 13948 24544 14000
rect 24860 13991 24912 14000
rect 24860 13957 24869 13991
rect 24869 13957 24903 13991
rect 24903 13957 24912 13991
rect 24860 13948 24912 13957
rect 25228 14016 25280 14068
rect 26700 13948 26752 14000
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 24584 13855 24636 13864
rect 24584 13821 24593 13855
rect 24593 13821 24627 13855
rect 24627 13821 24636 13855
rect 24584 13812 24636 13821
rect 26148 13812 26200 13864
rect 25964 13744 26016 13796
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 9128 13676 9180 13728
rect 9404 13719 9456 13728
rect 9404 13685 9413 13719
rect 9413 13685 9447 13719
rect 9447 13685 9456 13719
rect 9404 13676 9456 13685
rect 14280 13676 14332 13728
rect 18144 13676 18196 13728
rect 18236 13676 18288 13728
rect 18512 13676 18564 13728
rect 21088 13676 21140 13728
rect 21180 13676 21232 13728
rect 22376 13676 22428 13728
rect 27620 13676 27672 13728
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 4160 13472 4212 13524
rect 6460 13472 6512 13524
rect 6644 13404 6696 13456
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 4252 13268 4304 13320
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 7196 13336 7248 13388
rect 7656 13336 7708 13388
rect 4344 13268 4396 13277
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8300 13268 8352 13320
rect 8852 13268 8904 13320
rect 6000 13200 6052 13252
rect 9128 13404 9180 13456
rect 13820 13472 13872 13524
rect 15200 13472 15252 13524
rect 16948 13472 17000 13524
rect 14280 13404 14332 13456
rect 20444 13472 20496 13524
rect 11796 13336 11848 13388
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 17500 13404 17552 13456
rect 20812 13404 20864 13456
rect 24768 13472 24820 13524
rect 26148 13472 26200 13524
rect 27160 13472 27212 13524
rect 21180 13447 21232 13456
rect 21180 13413 21189 13447
rect 21189 13413 21223 13447
rect 21223 13413 21232 13447
rect 21180 13404 21232 13413
rect 23204 13404 23256 13456
rect 26240 13404 26292 13456
rect 15752 13336 15804 13388
rect 15844 13336 15896 13388
rect 15384 13311 15436 13320
rect 4804 13175 4856 13184
rect 4804 13141 4813 13175
rect 4813 13141 4847 13175
rect 4847 13141 4856 13175
rect 4804 13132 4856 13141
rect 6736 13132 6788 13184
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 12624 13200 12676 13252
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 16488 13268 16540 13320
rect 19156 13336 19208 13388
rect 19340 13336 19392 13388
rect 22008 13336 22060 13388
rect 22100 13336 22152 13388
rect 23572 13336 23624 13388
rect 25228 13336 25280 13388
rect 25596 13336 25648 13388
rect 18144 13268 18196 13320
rect 23112 13268 23164 13320
rect 26148 13336 26200 13388
rect 26332 13379 26384 13388
rect 26332 13345 26341 13379
rect 26341 13345 26375 13379
rect 26375 13345 26384 13379
rect 26332 13336 26384 13345
rect 27620 13336 27672 13388
rect 27896 13336 27948 13388
rect 12532 13132 12584 13184
rect 12992 13132 13044 13184
rect 16856 13200 16908 13252
rect 17408 13200 17460 13252
rect 19616 13200 19668 13252
rect 19708 13243 19760 13252
rect 19708 13209 19717 13243
rect 19717 13209 19751 13243
rect 19751 13209 19760 13243
rect 19708 13200 19760 13209
rect 18880 13132 18932 13184
rect 21180 13132 21232 13184
rect 21548 13200 21600 13252
rect 22192 13132 22244 13184
rect 22284 13132 22336 13184
rect 24308 13132 24360 13184
rect 24952 13200 25004 13252
rect 27896 13132 27948 13184
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 4344 12928 4396 12980
rect 9220 12928 9272 12980
rect 9404 12860 9456 12912
rect 9588 12860 9640 12912
rect 11704 12860 11756 12912
rect 11796 12860 11848 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 6460 12792 6512 12844
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 12532 12792 12584 12844
rect 15384 12928 15436 12980
rect 13636 12860 13688 12912
rect 15752 12903 15804 12912
rect 15752 12869 15761 12903
rect 15761 12869 15795 12903
rect 15795 12869 15804 12903
rect 15752 12860 15804 12869
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 4804 12656 4856 12708
rect 12808 12724 12860 12776
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 13084 12724 13136 12776
rect 16580 12724 16632 12776
rect 18144 12928 18196 12980
rect 21640 12928 21692 12980
rect 24124 12928 24176 12980
rect 24308 12971 24360 12980
rect 24308 12937 24317 12971
rect 24317 12937 24351 12971
rect 24351 12937 24360 12971
rect 24308 12928 24360 12937
rect 24768 12928 24820 12980
rect 26332 12928 26384 12980
rect 26608 12928 26660 12980
rect 18696 12860 18748 12912
rect 19708 12903 19760 12912
rect 19708 12869 19717 12903
rect 19717 12869 19751 12903
rect 19751 12869 19760 12903
rect 19708 12860 19760 12869
rect 22284 12860 22336 12912
rect 22836 12903 22888 12912
rect 22836 12869 22845 12903
rect 22845 12869 22879 12903
rect 22879 12869 22888 12903
rect 22836 12860 22888 12869
rect 24216 12860 24268 12912
rect 17776 12792 17828 12844
rect 18144 12792 18196 12844
rect 19340 12792 19392 12844
rect 24308 12792 24360 12844
rect 24584 12792 24636 12844
rect 24768 12835 24820 12844
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 28356 12835 28408 12844
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 4068 12588 4120 12640
rect 11152 12588 11204 12640
rect 11520 12588 11572 12640
rect 13084 12588 13136 12640
rect 14740 12656 14792 12708
rect 15292 12588 15344 12640
rect 16948 12631 17000 12640
rect 16948 12597 16957 12631
rect 16957 12597 16991 12631
rect 16991 12597 17000 12631
rect 16948 12588 17000 12597
rect 19800 12724 19852 12776
rect 22192 12724 22244 12776
rect 19248 12588 19300 12640
rect 20812 12656 20864 12708
rect 23204 12588 23256 12640
rect 25228 12588 25280 12640
rect 25596 12588 25648 12640
rect 26424 12588 26476 12640
rect 28172 12631 28224 12640
rect 28172 12597 28181 12631
rect 28181 12597 28215 12631
rect 28215 12597 28224 12631
rect 28172 12588 28224 12597
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 6828 12384 6880 12436
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 11060 12384 11112 12436
rect 11796 12427 11848 12436
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 11888 12384 11940 12436
rect 7748 12316 7800 12368
rect 9312 12316 9364 12368
rect 14096 12316 14148 12368
rect 15936 12384 15988 12436
rect 18144 12427 18196 12436
rect 18144 12393 18153 12427
rect 18153 12393 18187 12427
rect 18187 12393 18196 12427
rect 18144 12384 18196 12393
rect 22560 12384 22612 12436
rect 21548 12316 21600 12368
rect 23664 12316 23716 12368
rect 6368 12248 6420 12300
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 7196 12180 7248 12232
rect 11888 12248 11940 12300
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 13544 12248 13596 12300
rect 16580 12248 16632 12300
rect 16948 12248 17000 12300
rect 17408 12248 17460 12300
rect 19340 12248 19392 12300
rect 20628 12248 20680 12300
rect 20996 12248 21048 12300
rect 25044 12248 25096 12300
rect 9680 12180 9732 12232
rect 9772 12180 9824 12232
rect 11796 12180 11848 12232
rect 10232 12112 10284 12164
rect 6644 12044 6696 12096
rect 9588 12044 9640 12096
rect 11704 12044 11756 12096
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 12900 12180 12952 12232
rect 12808 12044 12860 12096
rect 13452 12044 13504 12096
rect 15936 12112 15988 12164
rect 17224 12180 17276 12232
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 22284 12223 22336 12232
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 23664 12180 23716 12232
rect 24400 12180 24452 12232
rect 24768 12180 24820 12232
rect 26240 12223 26292 12232
rect 26240 12189 26249 12223
rect 26249 12189 26283 12223
rect 26283 12189 26292 12223
rect 26240 12180 26292 12189
rect 16580 12155 16632 12164
rect 16580 12121 16589 12155
rect 16589 12121 16623 12155
rect 16623 12121 16632 12155
rect 16580 12112 16632 12121
rect 17500 12112 17552 12164
rect 17776 12112 17828 12164
rect 19892 12112 19944 12164
rect 19984 12155 20036 12164
rect 19984 12121 19993 12155
rect 19993 12121 20027 12155
rect 20027 12121 20036 12155
rect 19984 12112 20036 12121
rect 20996 12112 21048 12164
rect 21548 12112 21600 12164
rect 17224 12044 17276 12096
rect 17408 12044 17460 12096
rect 18696 12044 18748 12096
rect 22652 12112 22704 12164
rect 23480 12044 23532 12096
rect 23572 12044 23624 12096
rect 25872 12112 25924 12164
rect 26516 12155 26568 12164
rect 26516 12121 26525 12155
rect 26525 12121 26559 12155
rect 26559 12121 26568 12155
rect 26516 12112 26568 12121
rect 24308 12044 24360 12096
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 5908 11840 5960 11892
rect 8484 11840 8536 11892
rect 10232 11840 10284 11892
rect 13268 11840 13320 11892
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 6000 11704 6052 11756
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 1584 11636 1636 11688
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 8484 11679 8536 11688
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 8760 11772 8812 11824
rect 10140 11772 10192 11824
rect 10508 11815 10560 11824
rect 10508 11781 10517 11815
rect 10517 11781 10551 11815
rect 10551 11781 10560 11815
rect 10508 11772 10560 11781
rect 10692 11772 10744 11824
rect 10876 11772 10928 11824
rect 15752 11840 15804 11892
rect 16764 11840 16816 11892
rect 9588 11747 9640 11756
rect 9588 11713 9597 11747
rect 9597 11713 9631 11747
rect 9631 11713 9640 11747
rect 9588 11704 9640 11713
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 11888 11679 11940 11688
rect 7472 11568 7524 11620
rect 9680 11568 9732 11620
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 12532 11636 12584 11688
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 13728 11568 13780 11620
rect 14096 11815 14148 11824
rect 14096 11781 14105 11815
rect 14105 11781 14139 11815
rect 14139 11781 14148 11815
rect 19708 11840 19760 11892
rect 19984 11840 20036 11892
rect 23020 11840 23072 11892
rect 23940 11840 23992 11892
rect 14096 11772 14148 11781
rect 14004 11636 14056 11688
rect 14648 11636 14700 11688
rect 18972 11772 19024 11824
rect 22192 11772 22244 11824
rect 22376 11772 22428 11824
rect 23296 11772 23348 11824
rect 23848 11772 23900 11824
rect 17316 11704 17368 11756
rect 18052 11704 18104 11756
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 24584 11704 24636 11713
rect 18144 11636 18196 11688
rect 18236 11636 18288 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 18788 11636 18840 11688
rect 21088 11636 21140 11688
rect 23940 11636 23992 11688
rect 24032 11636 24084 11688
rect 24860 11679 24912 11688
rect 24860 11645 24869 11679
rect 24869 11645 24903 11679
rect 24903 11645 24912 11679
rect 24860 11636 24912 11645
rect 24952 11636 25004 11688
rect 16948 11568 17000 11620
rect 17224 11568 17276 11620
rect 7196 11500 7248 11552
rect 8760 11500 8812 11552
rect 9404 11500 9456 11552
rect 9588 11500 9640 11552
rect 12072 11500 12124 11552
rect 12716 11500 12768 11552
rect 13084 11500 13136 11552
rect 13268 11500 13320 11552
rect 17408 11500 17460 11552
rect 17776 11500 17828 11552
rect 20812 11500 20864 11552
rect 21548 11500 21600 11552
rect 26516 11500 26568 11552
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 5724 11296 5776 11348
rect 8484 11296 8536 11348
rect 9312 11296 9364 11348
rect 9588 11296 9640 11348
rect 12256 11296 12308 11348
rect 10692 11228 10744 11280
rect 10784 11228 10836 11280
rect 12992 11296 13044 11348
rect 14372 11296 14424 11348
rect 14556 11296 14608 11348
rect 15476 11296 15528 11348
rect 15568 11296 15620 11348
rect 16304 11296 16356 11348
rect 12624 11228 12676 11280
rect 9404 11160 9456 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 12072 11160 12124 11212
rect 17224 11228 17276 11280
rect 13636 11160 13688 11212
rect 17408 11160 17460 11212
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7288 11092 7340 11144
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 12624 11092 12676 11144
rect 12992 11092 13044 11144
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 10416 11024 10468 11076
rect 12348 11024 12400 11076
rect 14740 11092 14792 11144
rect 15752 11092 15804 11144
rect 15844 11024 15896 11076
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 18052 11296 18104 11348
rect 22652 11296 22704 11348
rect 23664 11339 23716 11348
rect 23664 11305 23673 11339
rect 23673 11305 23707 11339
rect 23707 11305 23716 11339
rect 23664 11296 23716 11305
rect 24492 11296 24544 11348
rect 26424 11296 26476 11348
rect 18144 11228 18196 11280
rect 19616 11160 19668 11212
rect 20628 11160 20680 11212
rect 22284 11160 22336 11212
rect 23020 11160 23072 11212
rect 24400 11228 24452 11280
rect 17776 11092 17828 11101
rect 19800 11092 19852 11144
rect 19892 11092 19944 11144
rect 21088 11092 21140 11144
rect 26148 11160 26200 11212
rect 26240 11160 26292 11212
rect 26608 11203 26660 11212
rect 26608 11169 26617 11203
rect 26617 11169 26651 11203
rect 26651 11169 26660 11203
rect 26608 11160 26660 11169
rect 24768 11092 24820 11144
rect 17224 11024 17276 11076
rect 21180 11024 21232 11076
rect 21640 11067 21692 11076
rect 21640 11033 21649 11067
rect 21649 11033 21683 11067
rect 21683 11033 21692 11067
rect 21640 11024 21692 11033
rect 10876 10956 10928 11008
rect 13728 10956 13780 11008
rect 13820 10956 13872 11008
rect 17776 10956 17828 11008
rect 17960 10956 18012 11008
rect 23940 11024 23992 11076
rect 24216 10956 24268 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 7288 10752 7340 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 9496 10795 9548 10804
rect 9496 10761 9505 10795
rect 9505 10761 9539 10795
rect 9539 10761 9548 10795
rect 9496 10752 9548 10761
rect 11888 10752 11940 10804
rect 12808 10795 12860 10804
rect 12808 10761 12817 10795
rect 12817 10761 12851 10795
rect 12851 10761 12860 10795
rect 12808 10752 12860 10761
rect 13360 10752 13412 10804
rect 13728 10727 13780 10736
rect 13728 10693 13737 10727
rect 13737 10693 13771 10727
rect 13771 10693 13780 10727
rect 13728 10684 13780 10693
rect 7748 10616 7800 10668
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 12256 10616 12308 10668
rect 13452 10616 13504 10668
rect 14280 10548 14332 10600
rect 17224 10752 17276 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 21180 10752 21232 10804
rect 21364 10795 21416 10804
rect 21364 10761 21373 10795
rect 21373 10761 21407 10795
rect 21407 10761 21416 10795
rect 21364 10752 21416 10761
rect 26608 10752 26660 10804
rect 29920 10752 29972 10804
rect 20260 10727 20312 10736
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 16948 10616 17000 10668
rect 20260 10693 20269 10727
rect 20269 10693 20303 10727
rect 20303 10693 20312 10727
rect 20260 10684 20312 10693
rect 17224 10548 17276 10600
rect 19616 10616 19668 10668
rect 21272 10657 21324 10668
rect 22284 10684 22336 10736
rect 22376 10727 22428 10736
rect 22376 10693 22385 10727
rect 22385 10693 22419 10727
rect 22419 10693 22428 10727
rect 22376 10684 22428 10693
rect 24124 10684 24176 10736
rect 21272 10623 21289 10657
rect 21289 10623 21323 10657
rect 21323 10623 21324 10657
rect 21272 10616 21324 10623
rect 23480 10616 23532 10668
rect 24216 10616 24268 10668
rect 18052 10548 18104 10600
rect 18236 10591 18288 10600
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 19064 10548 19116 10600
rect 19248 10548 19300 10600
rect 20536 10548 20588 10600
rect 20720 10548 20772 10600
rect 21548 10548 21600 10600
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24584 10616 24636 10668
rect 28080 10659 28132 10668
rect 28080 10625 28089 10659
rect 28089 10625 28123 10659
rect 28123 10625 28132 10659
rect 28080 10616 28132 10625
rect 24124 10548 24176 10557
rect 27804 10548 27856 10600
rect 12900 10480 12952 10532
rect 13176 10480 13228 10532
rect 16028 10523 16080 10532
rect 16028 10489 16037 10523
rect 16037 10489 16071 10523
rect 16071 10489 16080 10523
rect 16028 10480 16080 10489
rect 16488 10480 16540 10532
rect 17960 10480 18012 10532
rect 11796 10412 11848 10464
rect 12716 10412 12768 10464
rect 12992 10412 13044 10464
rect 22100 10480 22152 10532
rect 20352 10412 20404 10464
rect 24308 10480 24360 10532
rect 24216 10412 24268 10464
rect 26516 10455 26568 10464
rect 26516 10421 26525 10455
rect 26525 10421 26559 10455
rect 26559 10421 26568 10455
rect 26516 10412 26568 10421
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 3608 10004 3660 10056
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 10876 10208 10928 10260
rect 12716 10208 12768 10260
rect 22100 10208 22152 10260
rect 24032 10251 24084 10260
rect 24032 10217 24041 10251
rect 24041 10217 24075 10251
rect 24075 10217 24084 10251
rect 24032 10208 24084 10217
rect 25780 10208 25832 10260
rect 26424 10208 26476 10260
rect 17040 10140 17092 10192
rect 18144 10140 18196 10192
rect 10232 10072 10284 10124
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 10876 10004 10928 10056
rect 11704 10072 11756 10124
rect 13084 10072 13136 10124
rect 15292 10072 15344 10124
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 18052 10072 18104 10124
rect 20628 10072 20680 10124
rect 13268 10004 13320 10056
rect 17224 10004 17276 10056
rect 17408 10004 17460 10056
rect 12900 9936 12952 9988
rect 15292 9979 15344 9988
rect 15292 9945 15301 9979
rect 15301 9945 15335 9979
rect 15335 9945 15344 9979
rect 15292 9936 15344 9945
rect 15936 9936 15988 9988
rect 18420 9979 18472 9988
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 4896 9911 4948 9920
rect 4896 9877 4905 9911
rect 4905 9877 4939 9911
rect 4939 9877 4948 9911
rect 4896 9868 4948 9877
rect 9220 9868 9272 9920
rect 14556 9868 14608 9920
rect 14740 9868 14792 9920
rect 16948 9868 17000 9920
rect 18420 9945 18429 9979
rect 18429 9945 18463 9979
rect 18463 9945 18472 9979
rect 18420 9936 18472 9945
rect 18328 9868 18380 9920
rect 19340 9936 19392 9988
rect 20076 9979 20128 9988
rect 20076 9945 20085 9979
rect 20085 9945 20119 9979
rect 20119 9945 20128 9979
rect 20076 9936 20128 9945
rect 21088 9936 21140 9988
rect 18972 9868 19024 9920
rect 24216 10140 24268 10192
rect 22652 10072 22704 10124
rect 23204 10072 23256 10124
rect 24492 10072 24544 10124
rect 24584 10072 24636 10124
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 28356 10047 28408 10056
rect 28356 10013 28365 10047
rect 28365 10013 28399 10047
rect 28399 10013 28408 10047
rect 28356 10004 28408 10013
rect 22192 9936 22244 9988
rect 21456 9868 21508 9920
rect 21548 9868 21600 9920
rect 25872 9936 25924 9988
rect 26056 9868 26108 9920
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 3608 9707 3660 9716
rect 3608 9673 3617 9707
rect 3617 9673 3651 9707
rect 3651 9673 3660 9707
rect 3608 9664 3660 9673
rect 10784 9664 10836 9716
rect 11152 9664 11204 9716
rect 4896 9528 4948 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 12440 9596 12492 9648
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 11244 9528 11296 9580
rect 12808 9528 12860 9580
rect 14740 9664 14792 9716
rect 18328 9664 18380 9716
rect 18420 9664 18472 9716
rect 13728 9528 13780 9580
rect 15108 9571 15160 9580
rect 11980 9460 12032 9512
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 16672 9528 16724 9580
rect 17224 9596 17276 9648
rect 17408 9596 17460 9648
rect 18236 9639 18288 9648
rect 18236 9605 18245 9639
rect 18245 9605 18279 9639
rect 18279 9605 18288 9639
rect 18236 9596 18288 9605
rect 20076 9664 20128 9716
rect 20904 9664 20956 9716
rect 21272 9664 21324 9716
rect 17960 9571 18012 9580
rect 17960 9537 17969 9571
rect 17969 9537 18003 9571
rect 18003 9537 18012 9571
rect 17960 9528 18012 9537
rect 20260 9528 20312 9580
rect 20536 9528 20588 9580
rect 25044 9596 25096 9648
rect 22284 9528 22336 9580
rect 24584 9528 24636 9580
rect 26240 9528 26292 9580
rect 9312 9392 9364 9444
rect 17776 9460 17828 9512
rect 18788 9460 18840 9512
rect 21364 9460 21416 9512
rect 22468 9460 22520 9512
rect 13636 9435 13688 9444
rect 5908 9324 5960 9376
rect 8668 9324 8720 9376
rect 12624 9324 12676 9376
rect 13084 9367 13136 9376
rect 13084 9333 13093 9367
rect 13093 9333 13127 9367
rect 13127 9333 13136 9367
rect 13084 9324 13136 9333
rect 13636 9401 13645 9435
rect 13645 9401 13679 9435
rect 13679 9401 13688 9435
rect 13636 9392 13688 9401
rect 14096 9324 14148 9376
rect 17132 9324 17184 9376
rect 20076 9324 20128 9376
rect 20628 9324 20680 9376
rect 21456 9324 21508 9376
rect 24308 9367 24360 9376
rect 24308 9333 24317 9367
rect 24317 9333 24351 9367
rect 24351 9333 24360 9367
rect 24308 9324 24360 9333
rect 25780 9460 25832 9512
rect 27988 9528 28040 9580
rect 28448 9528 28500 9580
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 27896 9392 27948 9444
rect 27620 9324 27672 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 10876 9120 10928 9172
rect 11704 9120 11756 9172
rect 12440 9120 12492 9172
rect 13360 9120 13412 9172
rect 13636 9120 13688 9172
rect 15108 9120 15160 9172
rect 18052 9120 18104 9172
rect 24308 9120 24360 9172
rect 12164 9052 12216 9104
rect 14188 9052 14240 9104
rect 14740 9052 14792 9104
rect 16764 9052 16816 9104
rect 19156 9052 19208 9104
rect 4068 8984 4120 9036
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 10600 8984 10652 9036
rect 12992 8984 13044 9036
rect 16212 8984 16264 9036
rect 17960 8984 18012 9036
rect 18420 8984 18472 9036
rect 8484 8916 8536 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 8300 8848 8352 8900
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 11980 8916 12032 8968
rect 13452 8916 13504 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 20720 8984 20772 9036
rect 23112 9052 23164 9104
rect 24860 9120 24912 9172
rect 28264 9120 28316 9172
rect 21364 8984 21416 9036
rect 21640 8984 21692 9036
rect 22468 8984 22520 9036
rect 23848 8984 23900 9036
rect 24676 8984 24728 9036
rect 26424 8984 26476 9036
rect 27620 8984 27672 9036
rect 20812 8916 20864 8968
rect 22376 8916 22428 8968
rect 22836 8916 22888 8968
rect 23296 8959 23348 8968
rect 23296 8925 23305 8959
rect 23305 8925 23339 8959
rect 23339 8925 23348 8959
rect 23296 8916 23348 8925
rect 24768 8916 24820 8968
rect 9864 8848 9916 8900
rect 12808 8848 12860 8900
rect 1768 8780 1820 8832
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 10416 8780 10468 8832
rect 11244 8780 11296 8832
rect 13912 8780 13964 8832
rect 14740 8780 14792 8832
rect 16120 8891 16172 8900
rect 16120 8857 16129 8891
rect 16129 8857 16163 8891
rect 16163 8857 16172 8891
rect 16120 8848 16172 8857
rect 17408 8891 17460 8900
rect 16396 8780 16448 8832
rect 17408 8857 17417 8891
rect 17417 8857 17451 8891
rect 17451 8857 17460 8891
rect 17408 8848 17460 8857
rect 21180 8848 21232 8900
rect 18144 8780 18196 8832
rect 18788 8780 18840 8832
rect 20536 8780 20588 8832
rect 20628 8780 20680 8832
rect 22560 8848 22612 8900
rect 25136 8848 25188 8900
rect 26792 8848 26844 8900
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 8300 8576 8352 8628
rect 9404 8619 9456 8628
rect 9404 8585 9413 8619
rect 9413 8585 9447 8619
rect 9447 8585 9456 8619
rect 9404 8576 9456 8585
rect 9496 8576 9548 8628
rect 13636 8576 13688 8628
rect 16120 8576 16172 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17776 8576 17828 8628
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8668 8440 8720 8492
rect 11980 8508 12032 8560
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10416 8440 10468 8492
rect 13084 8508 13136 8560
rect 14832 8508 14884 8560
rect 17408 8508 17460 8560
rect 8944 8415 8996 8424
rect 8944 8381 8953 8415
rect 8953 8381 8987 8415
rect 8987 8381 8996 8415
rect 8944 8372 8996 8381
rect 10140 8372 10192 8424
rect 10784 8372 10836 8424
rect 13176 8440 13228 8492
rect 13820 8440 13872 8492
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 15200 8440 15252 8492
rect 15660 8440 15712 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17960 8508 18012 8560
rect 20352 8576 20404 8628
rect 20720 8576 20772 8628
rect 21640 8576 21692 8628
rect 22008 8576 22060 8628
rect 24124 8576 24176 8628
rect 28080 8619 28132 8628
rect 28080 8585 28089 8619
rect 28089 8585 28123 8619
rect 28123 8585 28132 8619
rect 28080 8576 28132 8585
rect 8760 8304 8812 8356
rect 9312 8304 9364 8356
rect 14188 8372 14240 8424
rect 13544 8304 13596 8356
rect 13728 8347 13780 8356
rect 13728 8313 13737 8347
rect 13737 8313 13771 8347
rect 13771 8313 13780 8347
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 17224 8372 17276 8424
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 19432 8440 19484 8492
rect 20352 8440 20404 8492
rect 20720 8440 20772 8492
rect 20812 8440 20864 8492
rect 21456 8508 21508 8560
rect 22192 8508 22244 8560
rect 22836 8508 22888 8560
rect 25320 8508 25372 8560
rect 26332 8508 26384 8560
rect 21364 8440 21416 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 19248 8372 19300 8424
rect 19708 8372 19760 8424
rect 21456 8372 21508 8424
rect 22652 8372 22704 8424
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 26516 8372 26568 8424
rect 13728 8304 13780 8313
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 6920 8236 6972 8288
rect 9772 8236 9824 8288
rect 14372 8236 14424 8288
rect 14464 8236 14516 8288
rect 14740 8236 14792 8288
rect 20168 8304 20220 8356
rect 20720 8347 20772 8356
rect 20720 8313 20729 8347
rect 20729 8313 20763 8347
rect 20763 8313 20772 8347
rect 20720 8304 20772 8313
rect 20812 8304 20864 8356
rect 23756 8347 23808 8356
rect 23756 8313 23765 8347
rect 23765 8313 23799 8347
rect 23799 8313 23808 8347
rect 23756 8304 23808 8313
rect 19340 8236 19392 8288
rect 21548 8236 21600 8288
rect 23388 8236 23440 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 8944 8032 8996 8084
rect 8300 7964 8352 8016
rect 11796 8032 11848 8084
rect 15292 8032 15344 8084
rect 17224 8032 17276 8084
rect 23388 8075 23440 8084
rect 12716 7964 12768 8016
rect 14372 7964 14424 8016
rect 19340 7964 19392 8016
rect 21456 7964 21508 8016
rect 23388 8041 23397 8075
rect 23397 8041 23431 8075
rect 23431 8041 23440 8075
rect 23388 8032 23440 8041
rect 23756 8032 23808 8084
rect 26056 8032 26108 8084
rect 27804 8032 27856 8084
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 6920 7828 6972 7880
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10508 7828 10560 7880
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 13452 7896 13504 7948
rect 14280 7896 14332 7948
rect 17040 7896 17092 7948
rect 17132 7896 17184 7948
rect 17868 7896 17920 7948
rect 17960 7896 18012 7948
rect 18144 7939 18196 7948
rect 18144 7905 18153 7939
rect 18153 7905 18187 7939
rect 18187 7905 18196 7939
rect 18144 7896 18196 7905
rect 19156 7896 19208 7948
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 24860 7964 24912 8016
rect 22284 7896 22336 7948
rect 12624 7871 12676 7880
rect 12624 7837 12633 7871
rect 12633 7837 12667 7871
rect 12667 7837 12676 7871
rect 12624 7828 12676 7837
rect 6460 7735 6512 7744
rect 6460 7701 6469 7735
rect 6469 7701 6503 7735
rect 6503 7701 6512 7735
rect 6460 7692 6512 7701
rect 6552 7692 6604 7744
rect 12164 7692 12216 7744
rect 14188 7760 14240 7812
rect 16120 7760 16172 7812
rect 16396 7803 16448 7812
rect 16396 7769 16405 7803
rect 16405 7769 16439 7803
rect 16439 7769 16448 7803
rect 16396 7760 16448 7769
rect 16672 7760 16724 7812
rect 17868 7803 17920 7812
rect 17868 7769 17877 7803
rect 17877 7769 17911 7803
rect 17911 7769 17920 7803
rect 17868 7760 17920 7769
rect 19708 7803 19760 7812
rect 16580 7692 16632 7744
rect 19708 7769 19717 7803
rect 19717 7769 19751 7803
rect 19751 7769 19760 7803
rect 19708 7760 19760 7769
rect 19800 7760 19852 7812
rect 23296 7896 23348 7948
rect 23756 7828 23808 7880
rect 24124 7896 24176 7948
rect 24584 7896 24636 7948
rect 18052 7692 18104 7744
rect 25964 7760 26016 7812
rect 26792 7803 26844 7812
rect 26792 7769 26801 7803
rect 26801 7769 26835 7803
rect 26835 7769 26844 7803
rect 26792 7760 26844 7769
rect 27804 7760 27856 7812
rect 22284 7692 22336 7744
rect 26056 7692 26108 7744
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 12440 7488 12492 7540
rect 13452 7488 13504 7540
rect 17684 7488 17736 7540
rect 17868 7488 17920 7540
rect 20904 7531 20956 7540
rect 8484 7463 8536 7472
rect 8484 7429 8493 7463
rect 8493 7429 8527 7463
rect 8527 7429 8536 7463
rect 8484 7420 8536 7429
rect 8668 7420 8720 7472
rect 11244 7420 11296 7472
rect 15752 7463 15804 7472
rect 15752 7429 15761 7463
rect 15761 7429 15795 7463
rect 15795 7429 15804 7463
rect 15752 7420 15804 7429
rect 16120 7420 16172 7472
rect 18788 7420 18840 7472
rect 20904 7497 20913 7531
rect 20913 7497 20947 7531
rect 20947 7497 20956 7531
rect 20904 7488 20956 7497
rect 21640 7488 21692 7540
rect 22744 7420 22796 7472
rect 22928 7488 22980 7540
rect 28264 7488 28316 7540
rect 24860 7420 24912 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 11060 7352 11112 7404
rect 12164 7352 12216 7404
rect 18696 7352 18748 7404
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 21364 7352 21416 7404
rect 22652 7352 22704 7404
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 23480 7352 23532 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 28172 7395 28224 7404
rect 11704 7327 11756 7336
rect 6828 7216 6880 7268
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 11980 7284 12032 7336
rect 11796 7216 11848 7268
rect 11888 7216 11940 7268
rect 13268 7284 13320 7336
rect 14648 7284 14700 7336
rect 16304 7284 16356 7336
rect 16856 7284 16908 7336
rect 17408 7284 17460 7336
rect 18236 7284 18288 7336
rect 21640 7284 21692 7336
rect 23572 7284 23624 7336
rect 24400 7327 24452 7336
rect 24400 7293 24409 7327
rect 24409 7293 24443 7327
rect 24443 7293 24452 7327
rect 24400 7284 24452 7293
rect 24860 7284 24912 7336
rect 28172 7361 28181 7395
rect 28181 7361 28215 7395
rect 28215 7361 28224 7395
rect 28172 7352 28224 7361
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 10784 7148 10836 7200
rect 11244 7148 11296 7200
rect 12440 7148 12492 7200
rect 12624 7148 12676 7200
rect 12808 7148 12860 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 15660 7148 15712 7200
rect 18880 7148 18932 7200
rect 19156 7148 19208 7200
rect 24124 7216 24176 7268
rect 27620 7148 27672 7200
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 8576 6944 8628 6996
rect 7656 6876 7708 6928
rect 11244 6944 11296 6996
rect 11704 6944 11756 6996
rect 11796 6944 11848 6996
rect 14464 6944 14516 6996
rect 18236 6944 18288 6996
rect 18512 6944 18564 6996
rect 20076 6944 20128 6996
rect 10140 6876 10192 6928
rect 12440 6876 12492 6928
rect 15660 6876 15712 6928
rect 16396 6876 16448 6928
rect 8852 6808 8904 6860
rect 17408 6808 17460 6860
rect 17500 6808 17552 6860
rect 7748 6740 7800 6792
rect 8760 6740 8812 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11796 6740 11848 6792
rect 12624 6740 12676 6792
rect 13912 6740 13964 6792
rect 15200 6740 15252 6792
rect 8484 6672 8536 6724
rect 9496 6672 9548 6724
rect 12900 6672 12952 6724
rect 16488 6740 16540 6792
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 16856 6672 16908 6724
rect 16580 6604 16632 6656
rect 17224 6604 17276 6656
rect 18512 6740 18564 6792
rect 18696 6808 18748 6860
rect 19340 6808 19392 6860
rect 20628 6808 20680 6860
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 22192 6851 22244 6860
rect 22192 6817 22201 6851
rect 22201 6817 22235 6851
rect 22235 6817 22244 6851
rect 22192 6808 22244 6817
rect 22652 6808 22704 6860
rect 23296 6808 23348 6860
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 18972 6740 19024 6792
rect 20352 6740 20404 6792
rect 19984 6672 20036 6724
rect 20444 6672 20496 6724
rect 20812 6672 20864 6724
rect 18144 6604 18196 6656
rect 21364 6604 21416 6656
rect 22284 6672 22336 6724
rect 23112 6715 23164 6724
rect 23112 6681 23121 6715
rect 23121 6681 23155 6715
rect 23155 6681 23164 6715
rect 23112 6672 23164 6681
rect 23388 6672 23440 6724
rect 24492 6808 24544 6860
rect 24584 6740 24636 6792
rect 26240 6740 26292 6792
rect 25412 6672 25464 6724
rect 27620 6672 27672 6724
rect 26516 6604 26568 6656
rect 29920 6740 29972 6792
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 7748 6400 7800 6452
rect 11060 6400 11112 6452
rect 5724 6332 5776 6384
rect 8668 6332 8720 6384
rect 9772 6332 9824 6384
rect 6828 6264 6880 6316
rect 7656 6264 7708 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 14556 6400 14608 6452
rect 14740 6400 14792 6452
rect 15016 6400 15068 6452
rect 16304 6400 16356 6452
rect 17316 6400 17368 6452
rect 18972 6400 19024 6452
rect 19156 6443 19208 6452
rect 19156 6409 19165 6443
rect 19165 6409 19199 6443
rect 19199 6409 19208 6443
rect 19156 6400 19208 6409
rect 19340 6400 19392 6452
rect 20444 6400 20496 6452
rect 12532 6332 12584 6384
rect 14372 6332 14424 6384
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 13176 6239 13228 6248
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 13728 6196 13780 6248
rect 14188 6264 14240 6316
rect 17132 6264 17184 6316
rect 14740 6239 14792 6248
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 9772 6128 9824 6180
rect 13084 6128 13136 6180
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 20352 6332 20404 6384
rect 19248 6264 19300 6316
rect 18236 6196 18288 6248
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 20628 6264 20680 6316
rect 23204 6332 23256 6384
rect 23664 6332 23716 6384
rect 24860 6332 24912 6384
rect 25136 6332 25188 6384
rect 20812 6264 20864 6316
rect 21548 6264 21600 6316
rect 23480 6264 23532 6316
rect 24768 6264 24820 6316
rect 18144 6128 18196 6180
rect 18880 6128 18932 6180
rect 21364 6196 21416 6248
rect 22560 6196 22612 6248
rect 22928 6196 22980 6248
rect 24676 6196 24728 6248
rect 25688 6239 25740 6248
rect 25688 6205 25697 6239
rect 25697 6205 25731 6239
rect 25731 6205 25740 6239
rect 25688 6196 25740 6205
rect 26608 6307 26660 6316
rect 26608 6273 26617 6307
rect 26617 6273 26651 6307
rect 26651 6273 26660 6307
rect 26608 6264 26660 6273
rect 27252 6264 27304 6316
rect 27804 6196 27856 6248
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 11888 6060 11940 6112
rect 15752 6060 15804 6112
rect 16856 6060 16908 6112
rect 20076 6060 20128 6112
rect 26240 6128 26292 6180
rect 28264 6171 28316 6180
rect 28264 6137 28273 6171
rect 28273 6137 28307 6171
rect 28307 6137 28316 6171
rect 28264 6128 28316 6137
rect 23664 6060 23716 6112
rect 28080 6060 28132 6112
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 8852 5856 8904 5908
rect 10968 5856 11020 5908
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 14464 5856 14516 5908
rect 12348 5788 12400 5840
rect 13084 5831 13136 5840
rect 13084 5797 13093 5831
rect 13093 5797 13127 5831
rect 13127 5797 13136 5831
rect 13084 5788 13136 5797
rect 13176 5788 13228 5840
rect 6552 5720 6604 5772
rect 10508 5720 10560 5772
rect 12532 5720 12584 5772
rect 15016 5763 15068 5772
rect 15016 5729 15025 5763
rect 15025 5729 15059 5763
rect 15059 5729 15068 5763
rect 15016 5720 15068 5729
rect 18880 5788 18932 5840
rect 19064 5856 19116 5908
rect 19616 5856 19668 5908
rect 23112 5856 23164 5908
rect 24952 5856 25004 5908
rect 25044 5856 25096 5908
rect 26608 5899 26660 5908
rect 26608 5865 26617 5899
rect 26617 5865 26651 5899
rect 26651 5865 26660 5899
rect 26608 5856 26660 5865
rect 27252 5899 27304 5908
rect 27252 5865 27261 5899
rect 27261 5865 27295 5899
rect 27295 5865 27304 5899
rect 27252 5856 27304 5865
rect 19892 5788 19944 5840
rect 20352 5788 20404 5840
rect 20812 5788 20864 5840
rect 21180 5788 21232 5840
rect 24676 5831 24728 5840
rect 24676 5797 24685 5831
rect 24685 5797 24719 5831
rect 24719 5797 24728 5831
rect 24676 5788 24728 5797
rect 22560 5720 22612 5772
rect 9312 5695 9364 5704
rect 3884 5584 3936 5636
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9496 5652 9548 5704
rect 11152 5652 11204 5704
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 12164 5652 12216 5704
rect 12900 5695 12952 5704
rect 12900 5661 12909 5695
rect 12909 5661 12943 5695
rect 12943 5661 12952 5695
rect 12900 5652 12952 5661
rect 13820 5652 13872 5704
rect 14464 5652 14516 5704
rect 16396 5695 16448 5704
rect 16396 5661 16405 5695
rect 16405 5661 16439 5695
rect 16439 5661 16448 5695
rect 16396 5652 16448 5661
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 19524 5652 19576 5704
rect 14648 5584 14700 5636
rect 20076 5652 20128 5704
rect 20352 5652 20404 5704
rect 20444 5652 20496 5704
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 23112 5652 23164 5704
rect 23296 5652 23348 5704
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24768 5652 24820 5704
rect 26056 5695 26108 5704
rect 26056 5661 26065 5695
rect 26065 5661 26099 5695
rect 26099 5661 26108 5695
rect 26056 5652 26108 5661
rect 27160 5695 27212 5704
rect 4252 5516 4304 5568
rect 6920 5516 6972 5568
rect 14280 5516 14332 5568
rect 20904 5584 20956 5636
rect 22744 5584 22796 5636
rect 27160 5661 27169 5695
rect 27169 5661 27203 5695
rect 27203 5661 27212 5695
rect 27160 5652 27212 5661
rect 21180 5516 21232 5568
rect 23664 5559 23716 5568
rect 23664 5525 23673 5559
rect 23673 5525 23707 5559
rect 23707 5525 23716 5559
rect 23664 5516 23716 5525
rect 26056 5516 26108 5568
rect 27896 5559 27948 5568
rect 27896 5525 27905 5559
rect 27905 5525 27939 5559
rect 27939 5525 27948 5559
rect 27896 5516 27948 5525
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 9864 5312 9916 5364
rect 11428 5312 11480 5364
rect 13728 5312 13780 5364
rect 14280 5312 14332 5364
rect 14740 5312 14792 5364
rect 17500 5312 17552 5364
rect 21088 5312 21140 5364
rect 21272 5312 21324 5364
rect 6460 5244 6512 5296
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 8944 5176 8996 5228
rect 14556 5244 14608 5296
rect 16028 5244 16080 5296
rect 18052 5244 18104 5296
rect 19340 5287 19392 5296
rect 19340 5253 19349 5287
rect 19349 5253 19383 5287
rect 19383 5253 19392 5287
rect 19340 5244 19392 5253
rect 23020 5244 23072 5296
rect 12348 5176 12400 5228
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 14280 5176 14332 5228
rect 15568 5176 15620 5228
rect 16856 5176 16908 5228
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 17316 5176 17368 5228
rect 18972 5176 19024 5228
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 23664 5176 23716 5228
rect 26056 5287 26108 5296
rect 26056 5253 26065 5287
rect 26065 5253 26099 5287
rect 26099 5253 26108 5287
rect 26056 5244 26108 5253
rect 26240 5244 26292 5296
rect 28080 5219 28132 5228
rect 28080 5185 28089 5219
rect 28089 5185 28123 5219
rect 28123 5185 28132 5219
rect 28080 5176 28132 5185
rect 15384 5108 15436 5160
rect 17868 5108 17920 5160
rect 11980 5040 12032 5092
rect 12992 5040 13044 5092
rect 19156 5040 19208 5092
rect 19432 5108 19484 5160
rect 20812 5151 20864 5160
rect 20812 5117 20821 5151
rect 20821 5117 20855 5151
rect 20855 5117 20864 5151
rect 20812 5108 20864 5117
rect 22744 5151 22796 5160
rect 20076 5040 20128 5092
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 12072 4972 12124 5024
rect 13544 5015 13596 5024
rect 13544 4981 13553 5015
rect 13553 4981 13587 5015
rect 13587 4981 13596 5015
rect 13544 4972 13596 4981
rect 14004 4972 14056 5024
rect 14648 4972 14700 5024
rect 20352 4972 20404 5024
rect 20720 5040 20772 5092
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 24676 5108 24728 5160
rect 27620 5108 27672 5160
rect 22928 5083 22980 5092
rect 22928 5049 22937 5083
rect 22937 5049 22971 5083
rect 22971 5049 22980 5083
rect 22928 5040 22980 5049
rect 22376 4972 22428 5024
rect 25872 4972 25924 5024
rect 28264 5015 28316 5024
rect 28264 4981 28273 5015
rect 28273 4981 28307 5015
rect 28307 4981 28316 5015
rect 28264 4972 28316 4981
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 9588 4768 9640 4820
rect 12164 4811 12216 4820
rect 12164 4777 12173 4811
rect 12173 4777 12207 4811
rect 12207 4777 12216 4811
rect 12164 4768 12216 4777
rect 13728 4768 13780 4820
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 17684 4768 17736 4820
rect 20812 4768 20864 4820
rect 20996 4768 21048 4820
rect 22376 4811 22428 4820
rect 22376 4777 22385 4811
rect 22385 4777 22419 4811
rect 22419 4777 22428 4811
rect 22376 4768 22428 4777
rect 23020 4811 23072 4820
rect 23020 4777 23029 4811
rect 23029 4777 23063 4811
rect 23063 4777 23072 4811
rect 23020 4768 23072 4777
rect 23204 4768 23256 4820
rect 26240 4768 26292 4820
rect 27160 4768 27212 4820
rect 27620 4811 27672 4820
rect 27620 4777 27629 4811
rect 27629 4777 27663 4811
rect 27663 4777 27672 4811
rect 27620 4768 27672 4777
rect 14188 4700 14240 4752
rect 14740 4700 14792 4752
rect 9680 4632 9732 4684
rect 6920 4564 6972 4616
rect 8668 4564 8720 4616
rect 12992 4564 13044 4616
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14648 4564 14700 4616
rect 11060 4496 11112 4548
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 11704 4428 11756 4480
rect 15200 4428 15252 4480
rect 18236 4632 18288 4684
rect 19708 4700 19760 4752
rect 20352 4700 20404 4752
rect 22836 4700 22888 4752
rect 24952 4700 25004 4752
rect 20536 4632 20588 4684
rect 18144 4564 18196 4616
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 20812 4564 20864 4616
rect 22284 4607 22336 4616
rect 19248 4496 19300 4548
rect 19984 4496 20036 4548
rect 22284 4573 22293 4607
rect 22293 4573 22327 4607
rect 22327 4573 22336 4607
rect 22284 4564 22336 4573
rect 26792 4632 26844 4684
rect 22192 4496 22244 4548
rect 23848 4564 23900 4616
rect 23940 4564 23992 4616
rect 25136 4564 25188 4616
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 25872 4564 25924 4573
rect 27528 4607 27580 4616
rect 27528 4573 27537 4607
rect 27537 4573 27571 4607
rect 27571 4573 27580 4607
rect 27528 4564 27580 4573
rect 27252 4496 27304 4548
rect 28080 4428 28132 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 17868 4224 17920 4276
rect 13544 4199 13596 4208
rect 13544 4165 13553 4199
rect 13553 4165 13587 4199
rect 13587 4165 13596 4199
rect 13544 4156 13596 4165
rect 7380 4088 7432 4140
rect 8944 4088 8996 4140
rect 11060 4088 11112 4140
rect 11244 4088 11296 4140
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 14188 4088 14240 4140
rect 14832 4088 14884 4140
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 14648 4020 14700 4072
rect 15568 4020 15620 4072
rect 9680 3952 9732 4004
rect 12256 3952 12308 4004
rect 5724 3884 5776 3936
rect 11980 3884 12032 3936
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 17960 4156 18012 4208
rect 18052 4088 18104 4140
rect 22744 4224 22796 4276
rect 23940 4267 23992 4276
rect 23940 4233 23949 4267
rect 23949 4233 23983 4267
rect 23983 4233 23992 4267
rect 23940 4224 23992 4233
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 19800 4088 19852 4140
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20904 4131 20956 4140
rect 20168 4088 20220 4097
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 22652 4020 22704 4072
rect 14556 3927 14608 3936
rect 12164 3884 12216 3893
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 17040 3884 17092 3936
rect 19340 3952 19392 4004
rect 19800 3952 19852 4004
rect 21640 3952 21692 4004
rect 23388 4131 23440 4140
rect 23388 4097 23397 4131
rect 23397 4097 23431 4131
rect 23431 4097 23440 4131
rect 23388 4088 23440 4097
rect 25964 4088 26016 4140
rect 24124 4020 24176 4072
rect 27804 4131 27856 4140
rect 27804 4097 27813 4131
rect 27813 4097 27847 4131
rect 27847 4097 27856 4131
rect 27804 4088 27856 4097
rect 25596 3952 25648 4004
rect 19708 3884 19760 3936
rect 20444 3884 20496 3936
rect 24032 3884 24084 3936
rect 26424 3952 26476 4004
rect 25780 3884 25832 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 12900 3680 12952 3732
rect 13728 3680 13780 3732
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 19616 3680 19668 3732
rect 18788 3612 18840 3664
rect 19340 3612 19392 3664
rect 14832 3544 14884 3596
rect 21456 3680 21508 3732
rect 21640 3680 21692 3732
rect 22376 3723 22428 3732
rect 21180 3655 21232 3664
rect 21180 3621 21189 3655
rect 21189 3621 21223 3655
rect 21223 3621 21232 3655
rect 21180 3612 21232 3621
rect 21548 3612 21600 3664
rect 22376 3689 22385 3723
rect 22385 3689 22419 3723
rect 22419 3689 22428 3723
rect 22376 3680 22428 3689
rect 23572 3680 23624 3732
rect 25044 3680 25096 3732
rect 26240 3723 26292 3732
rect 3976 3476 4028 3528
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12072 3476 12124 3528
rect 13452 3476 13504 3528
rect 15200 3476 15252 3528
rect 17592 3476 17644 3528
rect 17868 3476 17920 3528
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19524 3476 19576 3528
rect 20444 3476 20496 3528
rect 23296 3476 23348 3528
rect 26240 3689 26249 3723
rect 26249 3689 26283 3723
rect 26283 3689 26292 3723
rect 26240 3680 26292 3689
rect 27804 3680 27856 3732
rect 25780 3587 25832 3596
rect 25780 3553 25789 3587
rect 25789 3553 25823 3587
rect 25823 3553 25832 3587
rect 25780 3544 25832 3553
rect 25688 3476 25740 3528
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 27896 3476 27948 3528
rect 12440 3408 12492 3460
rect 14188 3408 14240 3460
rect 16672 3408 16724 3460
rect 19432 3408 19484 3460
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 17500 3340 17552 3392
rect 19248 3340 19300 3392
rect 23388 3340 23440 3392
rect 29920 3340 29972 3392
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 3884 3136 3936 3188
rect 5540 3136 5592 3188
rect 11888 3136 11940 3188
rect 14096 3136 14148 3188
rect 6000 3068 6052 3120
rect 2780 3000 2832 3052
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 15936 3068 15988 3120
rect 18144 3136 18196 3188
rect 18880 3136 18932 3188
rect 20812 3136 20864 3188
rect 22192 3136 22244 3188
rect 23388 3179 23440 3188
rect 8392 2932 8444 2984
rect 12164 3000 12216 3052
rect 13084 3000 13136 3052
rect 14556 3000 14608 3052
rect 7656 2864 7708 2916
rect 664 2796 716 2848
rect 5724 2796 5776 2848
rect 10416 2796 10468 2848
rect 16672 3000 16724 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 11244 2864 11296 2916
rect 18236 3000 18288 3052
rect 19800 3068 19852 3120
rect 20628 3000 20680 3052
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 23388 3145 23397 3179
rect 23397 3145 23431 3179
rect 23431 3145 23440 3179
rect 23388 3136 23440 3145
rect 25136 3136 25188 3188
rect 27528 3136 27580 3188
rect 25872 3068 25924 3120
rect 26424 3043 26476 3052
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 21548 2932 21600 2984
rect 19340 2864 19392 2916
rect 21456 2864 21508 2916
rect 26424 3009 26433 3043
rect 26433 3009 26467 3043
rect 26467 3009 26476 3043
rect 26424 3000 26476 3009
rect 28080 3043 28132 3052
rect 28080 3009 28089 3043
rect 28089 3009 28123 3043
rect 28123 3009 28132 3043
rect 28080 3000 28132 3009
rect 29092 2932 29144 2984
rect 12348 2796 12400 2848
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 15752 2796 15804 2848
rect 18788 2839 18840 2848
rect 18788 2805 18797 2839
rect 18797 2805 18831 2839
rect 18831 2805 18840 2839
rect 18788 2796 18840 2805
rect 19708 2796 19760 2848
rect 20260 2796 20312 2848
rect 27804 2796 27856 2848
rect 28356 2796 28408 2848
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 9036 2592 9088 2644
rect 9312 2592 9364 2644
rect 11152 2592 11204 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 18696 2592 18748 2644
rect 19524 2592 19576 2644
rect 20536 2635 20588 2644
rect 20536 2601 20545 2635
rect 20545 2601 20579 2635
rect 20579 2601 20588 2635
rect 20536 2592 20588 2601
rect 22652 2635 22704 2644
rect 22652 2601 22661 2635
rect 22661 2601 22695 2635
rect 22695 2601 22704 2635
rect 22652 2592 22704 2601
rect 24584 2635 24636 2644
rect 24584 2601 24593 2635
rect 24593 2601 24627 2635
rect 24627 2601 24636 2635
rect 24584 2592 24636 2601
rect 25872 2635 25924 2644
rect 25872 2601 25881 2635
rect 25881 2601 25915 2635
rect 25915 2601 25924 2635
rect 25872 2592 25924 2601
rect 25964 2592 26016 2644
rect 4252 2524 4304 2576
rect 1952 2388 2004 2440
rect 14464 2456 14516 2508
rect 22284 2524 22336 2576
rect 27252 2524 27304 2576
rect 5540 2388 5592 2440
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 7656 2388 7708 2440
rect 7748 2388 7800 2440
rect 9036 2388 9088 2440
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11612 2388 11664 2440
rect 12256 2388 12308 2440
rect 14648 2388 14700 2440
rect 15752 2388 15804 2440
rect 16120 2388 16172 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18788 2388 18840 2440
rect 20 2252 72 2304
rect 11796 2320 11848 2372
rect 20536 2388 20588 2440
rect 21456 2388 21508 2440
rect 22284 2388 22336 2440
rect 23204 2388 23256 2440
rect 24492 2388 24544 2440
rect 25412 2431 25464 2440
rect 25412 2397 25421 2431
rect 25421 2397 25455 2431
rect 25455 2397 25464 2431
rect 25412 2388 25464 2397
rect 25780 2388 25832 2440
rect 26424 2388 26476 2440
rect 27804 2431 27856 2440
rect 27804 2397 27813 2431
rect 27813 2397 27847 2431
rect 27847 2397 27856 2431
rect 27804 2388 27856 2397
rect 3240 2252 3292 2304
rect 4528 2252 4580 2304
rect 5816 2252 5868 2304
rect 6460 2252 6512 2304
rect 10324 2252 10376 2304
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 13544 2252 13596 2304
rect 14740 2252 14792 2304
rect 17408 2252 17460 2304
rect 27712 2252 27764 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 18696 1368 18748 1420
rect 20536 1368 20588 1420
<< metal2 >>
rect 662 29322 718 29800
rect 662 29294 1072 29322
rect 662 29200 718 29294
rect 1044 27606 1072 29294
rect 1950 29200 2006 29800
rect 2778 29336 2834 29345
rect 2778 29271 2834 29280
rect 3238 29322 3294 29800
rect 3882 29322 3938 29800
rect 5170 29322 5226 29800
rect 6458 29322 6514 29800
rect 7746 29322 7802 29800
rect 3238 29294 3464 29322
rect 1032 27600 1084 27606
rect 1032 27542 1084 27548
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 1860 27396 1912 27402
rect 1860 27338 1912 27344
rect 1688 27305 1716 27338
rect 1674 27296 1730 27305
rect 1674 27231 1730 27240
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1780 25945 1808 26318
rect 1766 25936 1822 25945
rect 1766 25871 1822 25880
rect 1768 24812 1820 24818
rect 1768 24754 1820 24760
rect 1780 24585 1808 24754
rect 1766 24576 1822 24585
rect 1766 24511 1822 24520
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1780 23225 1808 23666
rect 1766 23216 1822 23225
rect 1766 23151 1822 23160
rect 1872 22710 1900 27338
rect 1964 26994 1992 29200
rect 2792 27130 2820 29271
rect 3238 29200 3294 29294
rect 3146 27976 3202 27985
rect 3146 27911 3202 27920
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 3160 26994 3188 27911
rect 3436 27470 3464 29294
rect 3882 29294 4108 29322
rect 3882 29200 3938 29294
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3424 27464 3476 27470
rect 4080 27452 4108 29294
rect 5170 29294 5488 29322
rect 5170 29200 5226 29294
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 5460 27470 5488 29294
rect 6458 29294 6776 29322
rect 6458 29200 6514 29294
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 4160 27464 4212 27470
rect 4080 27424 4160 27452
rect 3424 27406 3476 27412
rect 4160 27406 4212 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 3252 27130 3280 27406
rect 3240 27124 3292 27130
rect 3240 27066 3292 27072
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 3148 26988 3200 26994
rect 3148 26930 3200 26936
rect 4252 26988 4304 26994
rect 4252 26930 4304 26936
rect 4264 26586 4292 26930
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4908 26586 4936 26862
rect 4252 26580 4304 26586
rect 4252 26522 4304 26528
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 5092 26042 5120 26318
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 1860 22704 1912 22710
rect 1860 22646 1912 22652
rect 1768 22024 1820 22030
rect 1768 21966 1820 21972
rect 1780 21865 1808 21966
rect 1766 21856 1822 21865
rect 1766 21791 1822 21800
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1768 19848 1820 19854
rect 1766 19816 1768 19825
rect 1820 19816 1822 19825
rect 1766 19751 1822 19760
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1780 18465 1808 18566
rect 1766 18456 1822 18465
rect 1766 18391 1822 18400
rect 1766 17096 1822 17105
rect 1766 17031 1768 17040
rect 1820 17031 1822 17040
rect 1768 17002 1820 17008
rect 3712 16114 3740 19654
rect 3988 16726 4016 20742
rect 4080 19854 4108 24550
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 6104 20942 6132 27542
rect 6748 27470 6776 29294
rect 7746 29294 8064 29322
rect 7746 29200 7802 29294
rect 7288 27532 7340 27538
rect 7288 27474 7340 27480
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6460 27328 6512 27334
rect 6460 27270 6512 27276
rect 6472 25906 6500 27270
rect 6460 25900 6512 25906
rect 6460 25842 6512 25848
rect 7300 21554 7328 27474
rect 8036 27470 8064 29294
rect 9034 29200 9090 29800
rect 10322 29200 10378 29800
rect 10966 29200 11022 29800
rect 12254 29322 12310 29800
rect 12254 29294 12388 29322
rect 12254 29200 12310 29294
rect 9048 27470 9076 29200
rect 10336 27606 10364 29200
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 10416 27464 10468 27470
rect 10980 27452 11008 29200
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11060 27464 11112 27470
rect 10980 27424 11060 27452
rect 10416 27406 10468 27412
rect 12360 27452 12388 29294
rect 13542 29200 13598 29800
rect 14830 29322 14886 29800
rect 14830 29294 15148 29322
rect 14830 29200 14886 29294
rect 13556 27606 13584 29200
rect 15120 27606 15148 29294
rect 16118 29200 16174 29800
rect 16762 29200 16818 29800
rect 18050 29200 18106 29800
rect 19338 29322 19394 29800
rect 19338 29294 19748 29322
rect 19338 29200 19394 29294
rect 16132 27606 16160 29200
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 12440 27464 12492 27470
rect 12360 27424 12440 27452
rect 11060 27406 11112 27412
rect 12440 27406 12492 27412
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 8312 23118 8340 26794
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8404 24206 8432 24754
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 8404 23662 8432 24142
rect 9232 23866 9260 24142
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9324 23730 9352 26454
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 9600 22658 9628 27270
rect 10428 26858 10456 27406
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 10416 26852 10468 26858
rect 10416 26794 10468 26800
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 9784 24682 9812 25842
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 9772 24676 9824 24682
rect 9772 24618 9824 24624
rect 9876 24342 9904 24754
rect 9864 24336 9916 24342
rect 9864 24278 9916 24284
rect 9600 22642 9812 22658
rect 9600 22636 9824 22642
rect 9600 22630 9772 22636
rect 9772 22578 9824 22584
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8772 22030 8800 22374
rect 9140 22166 9168 22510
rect 9128 22160 9180 22166
rect 9128 22102 9180 22108
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7392 21690 7420 21898
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 7380 21684 7432 21690
rect 7432 21644 7512 21672
rect 7380 21626 7432 21632
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 5080 20324 5132 20330
rect 5080 20266 5132 20272
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 5092 20058 5120 20266
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 17202 5396 17478
rect 5552 17202 5580 18022
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 5184 16794 5212 17138
rect 5736 17066 5764 20198
rect 6104 20058 6132 20334
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 1780 15745 1808 16050
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 1766 15736 1822 15745
rect 4423 15739 4731 15748
rect 1766 15671 1822 15680
rect 6196 15570 6224 20742
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6748 19378 6776 19790
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6748 18902 6776 19314
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6748 18358 6776 18838
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6840 17882 6868 18702
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6932 16454 6960 17274
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7024 16590 7052 16662
rect 7116 16590 7144 18634
rect 7392 18290 7420 19110
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7484 18222 7512 21644
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 8772 20466 8800 21830
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7208 16794 7236 17138
rect 7472 17128 7524 17134
rect 7392 17088 7472 17116
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 7116 16250 7144 16526
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 1768 14408 1820 14414
rect 1766 14376 1768 14385
rect 5816 14408 5868 14414
rect 1820 14376 1822 14385
rect 5816 14350 5868 14356
rect 1766 14311 1822 14320
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1780 13705 1808 13874
rect 1766 13696 1822 13705
rect 1766 13631 1822 13640
rect 3252 13326 3280 14010
rect 4908 13938 4936 14214
rect 5828 14074 5856 14350
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 6564 13938 6592 15846
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13530 4200 13806
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4264 12986 4292 13262
rect 4356 12986 4384 13262
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1780 12345 1808 12786
rect 4816 12714 4844 13126
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1596 11354 1624 11630
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10985 1808 11086
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9625 1808 9862
rect 3620 9722 3648 9998
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 4080 9042 4108 12582
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4816 10062 4844 12650
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5736 11354 5764 12174
rect 5920 11898 5948 12786
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6012 11762 6040 13194
rect 6380 12306 6408 13874
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6472 13530 6500 13806
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6472 12850 6500 13466
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6656 12102 6684 13398
rect 7208 13394 7236 13670
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12850 6776 13126
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6840 12442 6868 13262
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9586 4936 9862
rect 6656 9586 6684 12038
rect 7208 11762 7236 12174
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 11150 7236 11494
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7300 10810 7328 11086
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 5920 8974 5948 9318
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 1780 8498 1808 8774
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1766 8256 1822 8265
rect 1596 7410 1624 8230
rect 1766 8191 1822 8200
rect 1780 7886 1808 8191
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 6905 1808 7142
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 5736 6390 5764 8774
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7886 6960 8230
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 1766 6216 1822 6225
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4865 1808 4966
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1780 3398 1808 3431
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 3896 3194 3924 5578
rect 4172 5234 4200 6054
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 3534 4016 4966
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 32 800 60 2246
rect 676 800 704 2790
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1964 800 1992 2382
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 2792 785 2820 2994
rect 3160 2145 3188 2994
rect 4264 2582 4292 5510
rect 6472 5302 6500 7686
rect 6564 5778 6592 7686
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6840 6322 6868 7210
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 6932 4622 6960 5510
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 5552 2446 5580 3130
rect 5736 3058 5764 3878
rect 6012 3126 6040 4422
rect 7392 4146 7420 17088
rect 7472 17070 7524 17076
rect 7760 15638 7788 20198
rect 9140 19854 9168 22102
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9876 20466 9904 20742
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 9232 18834 9260 19654
rect 9968 19378 9996 21490
rect 10060 20466 10088 21830
rect 10244 20942 10272 26726
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 24274 10364 25094
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10428 23186 10456 23462
rect 10612 23322 10640 24006
rect 10704 23594 10732 24754
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10416 23180 10468 23186
rect 10416 23122 10468 23128
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10336 22098 10364 22374
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10520 22030 10548 22374
rect 10888 22234 10916 24686
rect 11072 24614 11100 25162
rect 11164 24682 11192 25230
rect 11152 24676 11204 24682
rect 11152 24618 11204 24624
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11072 23186 11100 23666
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 11256 23118 11284 25638
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11716 25294 11744 27270
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 25974 11836 26862
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11900 25974 11928 26522
rect 11992 26382 12020 27338
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12728 26382 12756 27270
rect 13188 27130 13216 27406
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13832 26450 13860 26726
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 11980 26240 12032 26246
rect 11980 26182 12032 26188
rect 11796 25968 11848 25974
rect 11796 25910 11848 25916
rect 11888 25968 11940 25974
rect 11888 25910 11940 25916
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11808 24818 11836 25094
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11900 24154 11928 25638
rect 11992 24954 12020 26182
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11992 24274 12020 24890
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11900 24126 12020 24154
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11808 22642 11836 23462
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11900 22778 11928 23054
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10336 21010 10364 21286
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 8312 18426 8340 18566
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 8312 17270 8340 18362
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 17882 8432 18226
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16590 8064 17070
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 8404 16114 8432 17614
rect 8588 16726 8616 18158
rect 9324 17882 9352 18702
rect 9876 18290 9904 19110
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9416 17746 9444 17818
rect 9692 17746 9720 18022
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9048 16017 9076 16050
rect 9232 16046 9260 17614
rect 9876 16658 9904 18090
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9220 16040 9272 16046
rect 9034 16008 9090 16017
rect 9220 15982 9272 15988
rect 9034 15943 9090 15952
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 9324 15502 9352 16050
rect 9784 16046 9812 16186
rect 9772 16040 9824 16046
rect 9968 16017 9996 19314
rect 10336 18834 10364 20742
rect 10520 20602 10548 20742
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10520 19802 10548 20538
rect 10428 19774 10548 19802
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10428 18970 10456 19774
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19378 10548 19654
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 10508 16040 10560 16046
rect 9772 15982 9824 15988
rect 9954 16008 10010 16017
rect 10244 15988 10508 15994
rect 10244 15982 10560 15988
rect 10244 15978 10548 15982
rect 9954 15943 10010 15952
rect 10232 15972 10548 15978
rect 10284 15966 10548 15972
rect 10232 15914 10284 15920
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9770 15600 9826 15609
rect 9770 15535 9826 15544
rect 9784 15502 9812 15535
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 7760 15162 7788 15438
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7668 12442 7696 13330
rect 8312 13326 8340 15302
rect 8404 14618 8432 15370
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8772 13938 8800 14282
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7484 8498 7512 11562
rect 7760 10674 7788 12310
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 8496 11898 8524 13806
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 8312 10810 8340 11630
rect 8496 11354 8524 11630
rect 8772 11558 8800 11766
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7760 7886 7788 10610
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 8312 8634 8340 8842
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8300 8016 8352 8022
rect 8404 8004 8432 9522
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8352 7976 8432 8004
rect 8300 7958 8352 7964
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 8496 7562 8524 8910
rect 8680 8498 8708 9318
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8404 7534 8524 7562
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 6322 7696 6870
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6458 7788 6734
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 8404 2990 8432 7534
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8496 6730 8524 7414
rect 8588 7002 8616 7822
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8680 6390 8708 7414
rect 8772 6798 8800 8298
rect 8864 6866 8892 13262
rect 9048 12782 9076 15370
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13462 9168 13670
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9232 12442 9260 12922
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9324 12374 9352 14962
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 12918 9444 13670
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9324 11354 9352 12310
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9416 11218 9444 11494
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9586 9260 9862
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9324 9450 9352 11018
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9324 8514 9352 8910
rect 9416 8634 9444 11154
rect 9508 10810 9536 13806
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12918 9628 13126
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9692 12238 9720 14826
rect 9784 12238 9812 15438
rect 9968 14618 9996 15642
rect 10612 15502 10640 16118
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10152 14482 10180 14758
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10414 14512 10470 14521
rect 10140 14476 10192 14482
rect 10414 14447 10470 14456
rect 10140 14418 10192 14424
rect 10428 14414 10456 14447
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10244 13938 10272 14214
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 10244 12170 10272 13262
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11762 9628 12038
rect 10244 11898 10272 12106
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10520 11830 10548 14554
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11354 9628 11494
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9692 11218 9720 11562
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 10152 10146 10180 11766
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10152 10130 10272 10146
rect 10152 10124 10284 10130
rect 10152 10118 10232 10124
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9508 8514 9536 8570
rect 9324 8486 9536 8514
rect 9876 8498 9904 8842
rect 9864 8492 9916 8498
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8956 8090 8984 8366
rect 9324 8362 9352 8486
rect 9864 8434 9916 8440
rect 10152 8430 10180 10118
rect 10232 10066 10284 10072
rect 10428 9586 10456 11018
rect 10612 9602 10640 13942
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10704 11286 10732 11766
rect 10796 11286 10824 19790
rect 10888 18290 10916 22170
rect 10980 21554 11008 22578
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 11072 22094 11100 22510
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11072 22066 11192 22094
rect 11164 21962 11192 22066
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 20602 11008 21490
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10980 19514 11008 20402
rect 11072 20398 11100 21830
rect 11164 20942 11192 21898
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 11072 18222 11100 19382
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11164 17762 11192 19654
rect 10980 17734 11192 17762
rect 10980 17542 11008 17734
rect 11256 17678 11284 21966
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11716 20466 11744 22442
rect 11992 22030 12020 24126
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 20942 11928 21286
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11716 19174 11744 20198
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11992 19514 12020 19790
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10968 16448 11020 16454
rect 10874 16416 10930 16425
rect 10968 16390 11020 16396
rect 10874 16351 10930 16360
rect 10888 15162 10916 16351
rect 10980 15910 11008 16390
rect 11072 16096 11100 17546
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17202 11192 17478
rect 11808 17338 11836 18702
rect 11900 18290 11928 18702
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11900 17202 11928 18090
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17678 12020 18022
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11256 16590 11284 17002
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11244 16108 11296 16114
rect 11072 16068 11192 16096
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10980 14906 11008 15846
rect 11072 15026 11100 15914
rect 11164 15706 11192 16068
rect 11244 16050 11296 16056
rect 11256 15706 11284 16050
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 15162 11192 15438
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10980 14878 11284 14906
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12442 11100 13262
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10796 11150 10824 11222
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10888 11014 10916 11766
rect 11164 11098 11192 12582
rect 11256 11234 11284 14878
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11532 12646 11560 13262
rect 11716 12918 11744 16662
rect 11992 16153 12020 17478
rect 12084 17218 12112 22918
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12176 21146 12204 21966
rect 12268 21350 12296 26250
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 12452 25265 12480 26182
rect 13372 25974 13400 26182
rect 13924 26042 13952 26930
rect 14280 26852 14332 26858
rect 14280 26794 14332 26800
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13268 25832 13320 25838
rect 13268 25774 13320 25780
rect 13280 25430 13308 25774
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 13176 25424 13228 25430
rect 13176 25366 13228 25372
rect 13268 25424 13320 25430
rect 13268 25366 13320 25372
rect 13084 25288 13136 25294
rect 12438 25256 12494 25265
rect 13084 25230 13136 25236
rect 12438 25191 12494 25200
rect 12452 23186 12480 25191
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12636 24070 12664 25094
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12176 20058 12204 20878
rect 12360 20346 12388 22578
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21486 12480 21966
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12268 20318 12388 20346
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12176 18426 12204 19178
rect 12268 19122 12296 20318
rect 12452 20262 12480 21286
rect 12544 20942 12572 22510
rect 12820 22094 12848 24142
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23730 12940 24006
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13004 23662 13032 24550
rect 13096 24410 13124 25230
rect 13188 24818 13216 25366
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12820 22066 13032 22094
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12636 21622 12664 21830
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12268 19094 12388 19122
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12268 18290 12296 18566
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12360 17785 12388 19094
rect 12346 17776 12402 17785
rect 12346 17711 12402 17720
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17338 12388 17614
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12084 17190 12388 17218
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 12084 16250 12112 16458
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11978 16144 12034 16153
rect 11978 16079 12034 16088
rect 12256 16108 12308 16114
rect 11992 14498 12020 16079
rect 12256 16050 12308 16056
rect 12268 15881 12296 16050
rect 12254 15872 12310 15881
rect 12254 15807 12310 15816
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11992 14470 12112 14498
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11808 13394 11836 13942
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11716 12434 11744 12854
rect 11808 12442 11836 12854
rect 11624 12406 11744 12434
rect 11796 12436 11848 12442
rect 11624 11642 11652 12406
rect 11796 12378 11848 12384
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11900 12306 11928 12378
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11762 11744 12038
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11624 11614 11744 11642
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11256 11218 11376 11234
rect 11256 11212 11388 11218
rect 11256 11206 11336 11212
rect 11336 11154 11388 11160
rect 10980 11070 11192 11098
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10266 10916 10950
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10796 9722 10824 9998
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10416 9580 10468 9586
rect 10612 9574 10824 9602
rect 10416 9522 10468 9528
rect 10140 8424 10192 8430
rect 10336 8401 10364 9522
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8498 10456 8774
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10140 8366 10192 8372
rect 10322 8392 10378 8401
rect 9312 8356 9364 8362
rect 10322 8327 10378 8336
rect 9312 8298 9364 8304
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9496 7880 9548 7886
rect 9548 7840 9720 7868
rect 9496 7822 9548 7828
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8864 5914 8892 6802
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4622 8708 4966
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8956 4146 8984 5170
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5736 2446 5764 2790
rect 7668 2446 7696 2858
rect 9048 2650 9076 6258
rect 9508 5710 9536 6666
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9324 2650 9352 5646
rect 9600 4826 9628 6734
rect 9692 6202 9720 7840
rect 9784 7410 9812 8230
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9784 6390 9812 7346
rect 10152 6934 10180 7822
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9692 6186 9812 6202
rect 9692 6180 9824 6186
rect 9692 6174 9772 6180
rect 9772 6122 9824 6128
rect 9876 5370 9904 6258
rect 10520 5778 10548 7822
rect 10612 6662 10640 8978
rect 10796 8430 10824 9574
rect 10888 9178 10916 9998
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 6798 10824 7142
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10980 5914 11008 11070
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11164 9722 11192 10610
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11716 10248 11744 11614
rect 11808 10470 11836 12174
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 10810 11928 11630
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11716 10220 11836 10248
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11256 8974 11284 9522
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11716 9178 11744 10066
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 7954 11284 8774
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11808 8090 11836 10220
rect 11992 9518 12020 14350
rect 12084 14006 12112 14470
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 11218 12112 11494
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 12176 9110 12204 15302
rect 12268 15094 12296 15807
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12360 14940 12388 17190
rect 12452 16658 12480 20198
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12636 19378 12664 19654
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12728 19258 12756 21626
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12636 19230 12756 19258
rect 12636 17218 12664 19230
rect 12820 18086 12848 20742
rect 13004 20602 13032 22066
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12544 17202 12664 17218
rect 12532 17196 12664 17202
rect 12584 17190 12664 17196
rect 12532 17138 12584 17144
rect 12544 16969 12572 17138
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12530 16960 12586 16969
rect 12530 16895 12586 16904
rect 12636 16794 12664 17070
rect 12714 16960 12770 16969
rect 12714 16895 12770 16904
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16250 12480 16390
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12440 14952 12492 14958
rect 12360 14912 12440 14940
rect 12440 14894 12492 14900
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 12238 12480 14758
rect 12544 13190 12572 16730
rect 12728 16114 12756 16895
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12532 12844 12584 12850
rect 12636 12832 12664 13194
rect 12584 12804 12664 12832
rect 12532 12786 12584 12792
rect 12728 12434 12756 15438
rect 12820 13870 12848 18022
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12912 15502 12940 17614
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 17066 13032 17546
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13096 15586 13124 22578
rect 13188 19417 13216 24142
rect 13740 22642 13768 25230
rect 13924 23186 13952 25434
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24818 14136 25094
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13636 22500 13688 22506
rect 13636 22442 13688 22448
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13280 19514 13308 19722
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13372 19446 13400 21014
rect 13450 20904 13506 20913
rect 13450 20839 13506 20848
rect 13464 20398 13492 20839
rect 13556 20398 13584 21490
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13360 19440 13412 19446
rect 13174 19408 13230 19417
rect 13360 19382 13412 19388
rect 13174 19343 13230 19352
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13004 15558 13124 15586
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 13004 15026 13032 15558
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13096 14074 13124 15438
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 13188 13802 13216 16050
rect 13280 15366 13308 18770
rect 13372 17338 13400 19382
rect 13556 19378 13584 19654
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13648 19310 13676 22442
rect 13740 22234 13768 22578
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13832 22166 13860 23054
rect 14016 22574 14044 23258
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 14200 22234 14228 26318
rect 14292 25702 14320 26794
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14384 25498 14412 27406
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 14752 26994 14780 27270
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 15672 27062 15700 27270
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14556 26784 14608 26790
rect 14556 26726 14608 26732
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 14568 25906 14596 26726
rect 15292 26512 15344 26518
rect 15292 26454 15344 26460
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 15304 25906 15332 26454
rect 15764 26382 15792 26726
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 15120 25226 15148 25638
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 15752 25220 15804 25226
rect 15752 25162 15804 25168
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24410 14412 25094
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 15764 24954 15792 25162
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14384 22506 14412 23054
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13648 17882 13676 18634
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13740 17678 13768 21830
rect 13832 21554 13860 22102
rect 14292 22098 14320 22374
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14384 21690 14412 21898
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13924 18426 13952 19246
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13372 15434 13400 17070
rect 13464 16425 13492 17206
rect 13450 16416 13506 16425
rect 13450 16351 13506 16360
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13464 15162 13492 16186
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15570 13584 15846
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13464 14482 13492 14826
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12866 13032 13126
rect 13004 12838 13216 12866
rect 13004 12782 13032 12838
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12544 12406 12756 12434
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12268 10674 12296 11290
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8566 12020 8910
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11256 7478 11284 7890
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 6458 11100 7346
rect 11992 7342 12020 8502
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7410 12204 7686
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 7002 11284 7142
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11716 7002 11744 7278
rect 11796 7268 11848 7274
rect 11796 7210 11848 7216
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11808 7002 11836 7210
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 4010 9720 4626
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 4146 11100 4490
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 10428 2446 10456 2790
rect 11164 2650 11192 5646
rect 11440 5370 11468 5646
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 4146 11744 4422
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11256 2922 11284 4082
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 3146 2136 3202 2145
rect 3146 2071 3202 2080
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 5828 800 5856 2246
rect 6472 800 6500 2246
rect 7760 800 7788 2382
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 9048 800 9076 2382
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 800 10364 2246
rect 11624 800 11652 2382
rect 11808 2378 11836 6734
rect 11900 6118 11928 7210
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 12360 5930 12388 11018
rect 12452 9654 12480 12174
rect 12544 11694 12572 12406
rect 12820 12186 12848 12718
rect 13096 12646 13124 12718
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13096 12306 13124 12582
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12728 12158 12848 12186
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12452 7546 12480 9114
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6934 12480 7142
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12544 6390 12572 11630
rect 12728 11558 12756 12158
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12636 11150 12664 11222
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12820 10810 12848 12038
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10538 12940 12174
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 13004 11354 13032 11630
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 13004 10470 13032 11086
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12728 10266 12756 10406
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 13096 10130 13124 11494
rect 13188 10538 13216 12838
rect 13556 12306 13584 15302
rect 13648 14006 13676 16118
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13648 12918 13676 13738
rect 13832 13530 13860 14758
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11898 13492 12038
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13280 11558 13308 11834
rect 13726 11792 13782 11801
rect 13726 11727 13782 11736
rect 13740 11626 13768 11727
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9489 12848 9522
rect 12806 9480 12862 9489
rect 12806 9415 12862 9424
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 7886 12664 9318
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6798 12664 7142
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12728 6322 12756 7958
rect 12820 7206 12848 8842
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12912 6730 12940 9930
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12268 5902 12388 5930
rect 12164 5704 12216 5710
rect 11978 5672 12034 5681
rect 12164 5646 12216 5652
rect 11978 5607 12034 5616
rect 11992 5098 12020 5607
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11900 3194 11928 4014
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11992 3534 12020 3878
rect 12084 3534 12112 4966
rect 12176 4826 12204 5646
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12268 4162 12296 5902
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12360 5234 12388 5782
rect 12544 5778 12572 6190
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12268 4134 12388 4162
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12176 3058 12204 3878
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12268 2446 12296 3946
rect 12360 3346 12388 4134
rect 12912 3738 12940 5646
rect 13004 5098 13032 8978
rect 13096 8566 13124 9318
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 6254 13216 8434
rect 13280 7342 13308 9998
rect 13372 9178 13400 10746
rect 13452 10668 13504 10674
rect 13556 10656 13584 11086
rect 13504 10628 13584 10656
rect 13452 10610 13504 10616
rect 13450 10568 13506 10577
rect 13450 10503 13506 10512
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13464 8974 13492 10503
rect 13452 8968 13504 8974
rect 13556 8945 13584 10628
rect 13648 9450 13676 11154
rect 13832 11014 13860 13466
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13740 10742 13768 10950
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13452 8910 13504 8916
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13648 8786 13676 9114
rect 13556 8758 13676 8786
rect 13556 8362 13584 8758
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13648 8537 13676 8570
rect 13634 8528 13690 8537
rect 13634 8463 13690 8472
rect 13740 8362 13768 9522
rect 13924 8838 13952 18226
rect 14108 14396 14136 19790
rect 14384 19514 14412 20198
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14384 18834 14412 19450
rect 14476 19394 14504 21490
rect 14568 19514 14596 24754
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 23662 14688 24550
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 14936 23322 14964 23462
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14752 22642 14780 22918
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 20942 14688 21830
rect 14752 21010 14780 22374
rect 15212 22166 15240 24006
rect 15304 23186 15332 24142
rect 15948 23798 15976 27270
rect 16776 27062 16804 29200
rect 18064 27606 18092 29200
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16120 26852 16172 26858
rect 16120 26794 16172 26800
rect 16132 24206 16160 26794
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16684 26450 16712 26726
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16868 25498 16896 27406
rect 17776 27396 17828 27402
rect 17776 27338 17828 27344
rect 17788 26994 17816 27338
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 16948 26920 17000 26926
rect 16948 26862 17000 26868
rect 16960 26586 16988 26862
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 17144 25786 17172 26930
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 16960 25758 17172 25786
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16488 25288 16540 25294
rect 16486 25256 16488 25265
rect 16540 25256 16542 25265
rect 16486 25191 16542 25200
rect 16500 24750 16528 25191
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15028 21962 15056 22034
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15028 21457 15056 21490
rect 15108 21480 15160 21486
rect 15014 21448 15070 21457
rect 15108 21422 15160 21428
rect 15014 21383 15070 21392
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14648 20936 14700 20942
rect 15120 20924 15148 21422
rect 15212 21078 15240 22102
rect 15396 21962 15424 23598
rect 15488 22710 15516 23666
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 15764 22710 15792 22918
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15948 22098 15976 23734
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15200 21072 15252 21078
rect 15200 21014 15252 21020
rect 15120 20896 15240 20924
rect 14648 20878 14700 20884
rect 15212 20806 15240 20896
rect 15580 20874 15608 21898
rect 15752 21616 15804 21622
rect 15752 21558 15804 21564
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 20058 14780 20334
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14476 19366 14688 19394
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14476 18358 14504 18566
rect 14568 18358 14596 18702
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14200 16250 14228 17206
rect 14292 16658 14320 17614
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14188 14408 14240 14414
rect 14108 14368 14188 14396
rect 14188 14350 14240 14356
rect 14200 13938 14228 14350
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 13938 14320 14214
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14292 13462 14320 13670
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14108 11830 14136 12310
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8498 13952 8774
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7546 13492 7890
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13096 5846 13124 6122
rect 13188 5846 13216 6190
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12990 4720 13046 4729
rect 12990 4655 13046 4664
rect 13004 4622 13032 4655
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12452 3346 12480 3402
rect 12360 3318 12480 3346
rect 12360 2854 12388 3318
rect 13096 3058 13124 5782
rect 13464 3534 13492 7482
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 6322 13676 7142
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13740 5370 13768 6190
rect 13832 5710 13860 8434
rect 13924 6798 13952 8434
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4214 13584 4966
rect 13740 4826 13768 5170
rect 14016 5030 14044 11630
rect 14384 11354 14412 18158
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16726 14596 17002
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14464 14952 14516 14958
rect 14660 14929 14688 19366
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 15212 17814 15240 20266
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16250 14780 17002
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14464 14894 14516 14900
rect 14646 14920 14702 14929
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10169 14320 10542
rect 14278 10160 14334 10169
rect 14278 10095 14334 10104
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13740 3738 13768 4558
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 14108 3194 14136 9318
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14200 8430 14228 9046
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14200 7818 14228 8366
rect 14292 7954 14320 8910
rect 14476 8294 14504 14894
rect 14556 14884 14608 14890
rect 14646 14855 14702 14864
rect 14556 14826 14608 14832
rect 14568 14074 14596 14826
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14568 12434 14596 13806
rect 14752 12714 14780 15370
rect 15212 15366 15240 17750
rect 15396 16658 15424 20742
rect 15672 20466 15700 21286
rect 15764 21146 15792 21558
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 16040 19938 16068 21966
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 15764 19910 16068 19938
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 18290 15516 18702
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15580 18426 15608 18634
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15672 18290 15700 19654
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15396 15434 15424 16594
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14844 14414 14872 14894
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 15304 14074 15332 14350
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15212 13530 15240 13942
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 15396 12986 15424 13262
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14568 12406 14688 12434
rect 14660 11694 14688 12406
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 9926 14596 11290
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14752 10674 14780 11086
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 15304 10130 15332 12582
rect 15488 11354 15516 16050
rect 15672 15978 15700 16050
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9722 14780 9862
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 9178 15148 9522
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14752 8838 14780 9046
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 8294 14780 8366
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14384 8022 14412 8230
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14476 7002 14504 8230
rect 14844 7970 14872 8502
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 14568 7942 14872 7970
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14568 6882 14596 7942
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14476 6854 14596 6882
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14476 6338 14504 6854
rect 14554 6760 14610 6769
rect 14554 6695 14610 6704
rect 14568 6458 14596 6695
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14200 4758 14228 6258
rect 14384 5914 14412 6326
rect 14476 6310 14596 6338
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14476 5710 14504 5850
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 5370 14320 5510
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14568 5302 14596 6310
rect 14660 5642 14688 7278
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6458 14780 7142
rect 15212 6798 15240 8434
rect 15304 8090 15332 9930
rect 15580 9586 15608 11290
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15566 9480 15622 9489
rect 15566 9415 15622 9424
rect 15382 8800 15438 8809
rect 15382 8735 15438 8744
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14752 5370 14780 6190
rect 15028 5778 15056 6394
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14292 4826 14320 5170
rect 15396 5166 15424 8735
rect 15580 5234 15608 9415
rect 15672 8498 15700 14486
rect 15764 13394 15792 19910
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19514 16068 19790
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15934 18864 15990 18873
rect 15934 18799 15936 18808
rect 15988 18799 15990 18808
rect 15936 18770 15988 18776
rect 16132 18290 16160 19994
rect 16224 18766 16252 23598
rect 16316 23050 16344 24278
rect 16960 23730 16988 25758
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 17144 25362 17172 25638
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16500 21894 16528 22918
rect 16868 22710 16896 22986
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21146 16620 21830
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16776 20874 16804 22374
rect 16856 22160 16908 22166
rect 16856 22102 16908 22108
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15856 16658 15884 17682
rect 15948 16658 15976 18226
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 14414 15884 15438
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14278 15884 14350
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15764 11898 15792 12854
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15752 11144 15804 11150
rect 15750 11112 15752 11121
rect 15804 11112 15806 11121
rect 15856 11082 15884 13330
rect 15948 12442 15976 14962
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15750 11047 15806 11056
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15948 9994 15976 12106
rect 16040 10538 16068 17274
rect 16132 16454 16160 17614
rect 16224 16454 16252 18566
rect 16316 18290 16344 19110
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16592 17202 16620 17614
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 6934 15700 7142
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15764 6118 15792 7414
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14660 4622 14688 4966
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14200 3466 14228 4082
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 14476 2514 14504 4558
rect 14648 4072 14700 4078
rect 14752 4026 14780 4694
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14700 4020 14780 4026
rect 14648 4014 14780 4020
rect 14660 3998 14780 4014
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3058 14596 3878
rect 14752 3738 14780 3998
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14844 3602 14872 4082
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 15212 3534 15240 4422
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15580 3738 15608 4014
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 15948 3126 15976 9930
rect 16132 9874 16160 11018
rect 16040 9846 16160 9874
rect 16040 5302 16068 9846
rect 16224 9042 16252 16390
rect 16316 15434 16344 16594
rect 16394 15872 16450 15881
rect 16394 15807 16450 15816
rect 16408 15434 16436 15807
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16316 11354 16344 15370
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16500 14822 16528 15030
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16500 13841 16528 14282
rect 16592 14074 16620 15302
rect 16684 14822 16712 20810
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19786 16804 20198
rect 16868 19922 16896 22102
rect 17052 21146 17080 22578
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16960 18358 16988 19246
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 17052 17814 17080 18294
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17144 17270 17172 20402
rect 17236 18222 17264 25842
rect 17696 24410 17724 26862
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 17960 25696 18012 25702
rect 17960 25638 18012 25644
rect 17684 24404 17736 24410
rect 17604 24364 17684 24392
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17512 23118 17540 23462
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17512 20466 17540 22578
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17420 19281 17448 19314
rect 17406 19272 17462 19281
rect 17406 19207 17462 19216
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17420 18358 17448 18566
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17144 16590 17172 17206
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 16250 17172 16390
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 14618 16712 14758
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16868 14482 16896 14894
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16486 13832 16542 13841
rect 16486 13767 16542 13776
rect 16592 13716 16620 14010
rect 16960 13870 16988 15574
rect 17052 15162 17080 15982
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17236 14482 17264 18158
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17420 15065 17448 17138
rect 17512 16182 17540 19654
rect 17604 19378 17632 24364
rect 17684 24346 17736 24352
rect 17972 23730 18000 25638
rect 18156 25294 18184 26182
rect 18708 25838 18736 26726
rect 18800 26450 18828 26998
rect 18880 26512 18932 26518
rect 18880 26454 18932 26460
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18248 25498 18276 25774
rect 18892 25702 18920 26454
rect 18972 26376 19024 26382
rect 18972 26318 19024 26324
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18800 24206 18828 24686
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17696 23118 17724 23666
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17788 22080 17816 23462
rect 18156 23322 18184 24142
rect 18604 24064 18656 24070
rect 18656 24024 18736 24052
rect 18604 24006 18656 24012
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17880 22642 17908 22918
rect 18708 22778 18736 24024
rect 18800 23594 18828 24142
rect 18892 23798 18920 25638
rect 18984 25294 19012 26318
rect 19064 26308 19116 26314
rect 19064 26250 19116 26256
rect 18972 25288 19024 25294
rect 18972 25230 19024 25236
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 18788 23588 18840 23594
rect 18788 23530 18840 23536
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 17696 22052 17816 22080
rect 18052 22092 18104 22098
rect 17696 21486 17724 22052
rect 18052 22034 18104 22040
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17788 21622 17816 21898
rect 17776 21616 17828 21622
rect 17776 21558 17828 21564
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17788 20058 17816 21422
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17788 19854 17816 19994
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17604 17678 17632 19314
rect 17880 18698 17908 21286
rect 17972 20466 18000 21422
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17972 20058 18000 20402
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17972 19378 18000 19994
rect 18064 19718 18092 22034
rect 18708 22030 18736 22714
rect 18788 22568 18840 22574
rect 18786 22536 18788 22545
rect 18840 22536 18842 22545
rect 18786 22471 18842 22480
rect 18892 22438 18920 22918
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18510 21720 18566 21729
rect 18510 21655 18566 21664
rect 18524 21622 18552 21655
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18142 20632 18198 20641
rect 18248 20602 18276 21422
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18708 20942 18736 21966
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18142 20567 18144 20576
rect 18196 20567 18198 20576
rect 18236 20596 18288 20602
rect 18144 20538 18196 20544
rect 18236 20538 18288 20544
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18144 19848 18196 19854
rect 18142 19816 18144 19825
rect 18196 19816 18198 19825
rect 18142 19751 18198 19760
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17972 17814 18000 18838
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 18064 17746 18092 18158
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 17338 17632 17478
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17406 15056 17462 15065
rect 17406 14991 17462 15000
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17328 14362 17356 14418
rect 17420 14414 17448 14991
rect 17236 14334 17356 14362
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16408 13688 16620 13716
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16408 9674 16436 13688
rect 16960 13530 16988 13806
rect 17040 13796 17092 13802
rect 17040 13738 17092 13744
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16488 13320 16540 13326
rect 16670 13288 16726 13297
rect 16540 13268 16670 13274
rect 16488 13262 16670 13268
rect 16500 13246 16670 13262
rect 16670 13223 16726 13232
rect 16856 13252 16908 13258
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16592 12345 16620 12718
rect 16578 12336 16634 12345
rect 16578 12271 16580 12280
rect 16632 12271 16634 12280
rect 16580 12242 16632 12248
rect 16592 12211 16620 12242
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16316 9646 16436 9674
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16132 8634 16160 8842
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16132 7478 16160 7754
rect 16120 7472 16172 7478
rect 16120 7414 16172 7420
rect 16316 7342 16344 9646
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 7818 16436 8774
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16500 7018 16528 10474
rect 16592 8242 16620 12106
rect 16684 9586 16712 13223
rect 16856 13194 16908 13200
rect 16764 11892 16816 11898
rect 16868 11880 16896 13194
rect 16948 12640 17000 12646
rect 16946 12608 16948 12617
rect 17000 12608 17002 12617
rect 16946 12543 17002 12552
rect 17052 12434 17080 13738
rect 17236 12434 17264 14334
rect 17420 14278 17448 14350
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17512 13462 17540 16118
rect 17604 15502 17632 16526
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17880 16402 17908 17070
rect 17972 16590 18000 17546
rect 18064 17202 18092 17682
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18156 16590 18184 18702
rect 18248 17678 18276 19926
rect 18432 19904 18460 19994
rect 18604 19916 18656 19922
rect 18432 19876 18604 19904
rect 18604 19858 18656 19864
rect 18696 19848 18748 19854
rect 18694 19816 18696 19825
rect 18748 19816 18750 19825
rect 18694 19751 18750 19760
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19446 18736 19654
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18328 18624 18380 18630
rect 18432 18612 18460 18702
rect 18380 18584 18460 18612
rect 18328 18566 18380 18572
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18616 17105 18644 17206
rect 18602 17096 18658 17105
rect 18602 17031 18658 17040
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17052 12406 17172 12434
rect 17236 12406 17356 12434
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16816 11852 16896 11880
rect 16764 11834 16816 11840
rect 16960 11778 16988 12242
rect 16868 11750 16988 11778
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16764 9104 16816 9110
rect 16762 9072 16764 9081
rect 16816 9072 16818 9081
rect 16762 9007 16818 9016
rect 16592 8214 16804 8242
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16316 6990 16528 7018
rect 16316 6458 16344 6990
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16408 5710 16436 6870
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16500 5710 16528 6734
rect 16592 6662 16620 7686
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16396 5704 16448 5710
rect 16394 5672 16396 5681
rect 16488 5704 16540 5710
rect 16448 5672 16450 5681
rect 16488 5646 16540 5652
rect 16394 5607 16450 5616
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 16684 3466 16712 7754
rect 16776 6712 16804 8214
rect 16868 7342 16896 11750
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16960 10674 16988 11562
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16960 8634 16988 9862
rect 17052 9625 17080 10134
rect 17144 10044 17172 12406
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 12102 17264 12174
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17328 11762 17356 12406
rect 17420 12306 17448 13194
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 11620 17276 11626
rect 17224 11562 17276 11568
rect 17236 11286 17264 11562
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17222 11112 17278 11121
rect 17222 11047 17224 11056
rect 17276 11047 17278 11056
rect 17224 11018 17276 11024
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17236 10606 17264 10746
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17224 10056 17276 10062
rect 17144 10016 17224 10044
rect 17038 9616 17094 9625
rect 17038 9551 17094 9560
rect 17144 9466 17172 10016
rect 17224 9998 17276 10004
rect 17224 9648 17276 9654
rect 17222 9616 17224 9625
rect 17276 9616 17278 9625
rect 17222 9551 17278 9560
rect 17052 9438 17172 9466
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17052 7954 17080 9438
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 8498 17172 9318
rect 17222 8528 17278 8537
rect 17132 8492 17184 8498
rect 17222 8463 17278 8472
rect 17132 8434 17184 8440
rect 17236 8430 17264 8463
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 17144 6798 17172 7890
rect 17236 6798 17264 8026
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16856 6724 16908 6730
rect 16776 6684 16856 6712
rect 16856 6666 16908 6672
rect 16868 6118 16896 6666
rect 17144 6322 17172 6734
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 17144 5234 17172 6258
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17132 5228 17184 5234
rect 17236 5216 17264 6598
rect 17328 6458 17356 11698
rect 17420 11558 17448 12038
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17406 11248 17462 11257
rect 17406 11183 17408 11192
rect 17460 11183 17462 11192
rect 17408 11154 17460 11160
rect 17512 10810 17540 12106
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9654 17448 9998
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17420 8566 17448 8842
rect 17408 8560 17460 8566
rect 17406 8528 17408 8537
rect 17460 8528 17462 8537
rect 17406 8463 17462 8472
rect 17408 7336 17460 7342
rect 17406 7304 17408 7313
rect 17460 7304 17462 7313
rect 17406 7239 17462 7248
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17420 6254 17448 6802
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17512 5370 17540 6802
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17316 5228 17368 5234
rect 17236 5188 17316 5216
rect 17132 5170 17184 5176
rect 17316 5170 17368 5176
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 16684 3058 16712 3402
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14660 2446 14688 2790
rect 15764 2446 15792 2790
rect 16868 2650 16896 5170
rect 17604 4808 17632 14486
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 11880 17724 14350
rect 17788 13802 17816 16390
rect 17880 16374 18000 16402
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17880 15609 17908 16050
rect 17866 15600 17922 15609
rect 17866 15535 17922 15544
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17880 14482 17908 15438
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 14278 17908 14418
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17972 14074 18000 16374
rect 18156 15502 18184 16526
rect 18708 16114 18736 17682
rect 18800 17542 18828 22170
rect 18892 18306 18920 22170
rect 18984 21486 19012 25230
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19076 21332 19104 26250
rect 19248 25220 19300 25226
rect 19248 25162 19300 25168
rect 19260 24750 19288 25162
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19352 24698 19380 27066
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19444 26586 19472 26930
rect 19628 26586 19656 27406
rect 19720 26994 19748 29294
rect 20626 29200 20682 29800
rect 21914 29200 21970 29800
rect 23202 29322 23258 29800
rect 23846 29322 23902 29800
rect 23202 29294 23428 29322
rect 23202 29200 23258 29294
rect 20640 27554 20668 29200
rect 20720 27600 20772 27606
rect 20640 27548 20720 27554
rect 20640 27542 20772 27548
rect 20640 27526 20760 27542
rect 21364 27464 21416 27470
rect 21928 27452 21956 29200
rect 23400 27554 23428 29294
rect 23846 29294 24256 29322
rect 23846 29200 23902 29294
rect 23480 27600 23532 27606
rect 23400 27548 23480 27554
rect 23400 27542 23532 27548
rect 23400 27526 23520 27542
rect 22100 27464 22152 27470
rect 21928 27424 22100 27452
rect 21364 27406 21416 27412
rect 22100 27406 22152 27412
rect 19708 26988 19760 26994
rect 19708 26930 19760 26936
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 19708 26852 19760 26858
rect 19708 26794 19760 26800
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19444 25974 19472 26318
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19352 24670 19472 24698
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 19168 24154 19196 24278
rect 19168 24126 19288 24154
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 19168 23798 19196 24006
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 19168 22234 19196 23054
rect 19260 22794 19288 24126
rect 19352 22982 19380 24550
rect 19444 23746 19472 24670
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19536 24313 19564 24550
rect 19616 24336 19668 24342
rect 19522 24304 19578 24313
rect 19616 24278 19668 24284
rect 19522 24239 19578 24248
rect 19628 24206 19656 24278
rect 19720 24274 19748 26794
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19812 24342 19840 24686
rect 19800 24336 19852 24342
rect 19800 24278 19852 24284
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19616 24200 19668 24206
rect 19614 24168 19616 24177
rect 19668 24168 19670 24177
rect 19614 24103 19670 24112
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19444 23718 19564 23746
rect 19536 23662 19564 23718
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19260 22766 19380 22794
rect 19444 22778 19472 23598
rect 19628 23066 19656 24006
rect 19720 23866 19748 24210
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19720 23474 19748 23598
rect 19904 23497 19932 26726
rect 20732 26586 20760 26862
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19996 24206 20024 25230
rect 20180 25158 20208 26318
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 20272 24970 20300 25230
rect 20180 24942 20300 24970
rect 20904 24948 20956 24954
rect 20180 24818 20208 24942
rect 20904 24890 20956 24896
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 24274 20116 24550
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19890 23488 19946 23497
rect 19720 23446 19840 23474
rect 19706 23352 19762 23361
rect 19706 23287 19762 23296
rect 19536 23050 19656 23066
rect 19524 23044 19656 23050
rect 19576 23038 19656 23044
rect 19524 22986 19576 22992
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 19352 22094 19380 22766
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19444 22234 19472 22510
rect 19628 22438 19656 23038
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19352 22066 19472 22094
rect 19248 21480 19300 21486
rect 19246 21448 19248 21457
rect 19300 21448 19302 21457
rect 19246 21383 19302 21392
rect 18984 21304 19104 21332
rect 18984 18834 19012 21304
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19076 18902 19104 20198
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 19062 18320 19118 18329
rect 18892 18278 19062 18306
rect 19062 18255 19118 18264
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18708 15570 18736 16050
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18248 15026 18276 15506
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 15094 18644 15302
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18156 13818 18184 14894
rect 18248 13988 18276 14962
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18800 14414 18828 15438
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18328 14000 18380 14006
rect 18248 13960 18328 13988
rect 18328 13942 18380 13948
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 18064 13790 18184 13818
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12170 17816 12786
rect 18064 12238 18092 13790
rect 18524 13734 18552 13806
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18156 13433 18184 13670
rect 18142 13424 18198 13433
rect 18142 13359 18198 13368
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18156 12986 18184 13262
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18156 12442 18184 12786
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17696 11852 17908 11880
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 11150 17816 11494
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10130 17816 10950
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 8634 17816 9454
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17880 7954 17908 11852
rect 18248 11801 18276 13670
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18708 12918 18736 14010
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18708 12238 18736 12854
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18696 12096 18748 12102
rect 18800 12050 18828 13806
rect 18892 13433 18920 18158
rect 18970 16824 19026 16833
rect 18970 16759 19026 16768
rect 18984 16726 19012 16759
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18970 16144 19026 16153
rect 18970 16079 19026 16088
rect 18984 16046 19012 16079
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 19076 14958 19104 18255
rect 19168 17921 19196 20742
rect 19260 19922 19288 20946
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20346 19380 20878
rect 19444 20466 19472 22066
rect 19536 22030 19564 22374
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19616 21412 19668 21418
rect 19616 21354 19668 21360
rect 19628 21146 19656 21354
rect 19720 21350 19748 23287
rect 19812 23050 19840 23446
rect 19890 23423 19946 23432
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19904 22778 19932 23258
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19536 20369 19564 20878
rect 19720 20534 19748 21286
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19522 20360 19578 20369
rect 19352 20330 19472 20346
rect 19352 20324 19484 20330
rect 19352 20318 19432 20324
rect 19522 20295 19578 20304
rect 19432 20266 19484 20272
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19260 18834 19288 19858
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19154 17912 19210 17921
rect 19154 17847 19210 17856
rect 19154 16688 19210 16697
rect 19260 16658 19288 18770
rect 19352 16726 19380 20198
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19444 18068 19472 19790
rect 19628 19718 19656 20402
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19536 18193 19564 18362
rect 19522 18184 19578 18193
rect 19522 18119 19578 18128
rect 19616 18080 19668 18086
rect 19444 18040 19616 18068
rect 19616 18022 19668 18028
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19154 16623 19210 16632
rect 19248 16652 19300 16658
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 18878 13424 18934 13433
rect 19168 13394 19196 16623
rect 19248 16594 19300 16600
rect 19248 16176 19300 16182
rect 19246 16144 19248 16153
rect 19300 16144 19302 16153
rect 19246 16079 19302 16088
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19260 14482 19288 15506
rect 19352 15434 19380 16662
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19522 16416 19578 16425
rect 19522 16351 19578 16360
rect 19536 16046 19564 16351
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19628 15434 19656 16458
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19628 14890 19656 15370
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19260 13818 19288 14418
rect 19628 14414 19656 14826
rect 19720 14793 19748 16934
rect 19706 14784 19762 14793
rect 19706 14719 19762 14728
rect 19340 14408 19392 14414
rect 19616 14408 19668 14414
rect 19392 14368 19564 14396
rect 19340 14350 19392 14356
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19260 13790 19380 13818
rect 19352 13394 19380 13790
rect 19444 13705 19472 13942
rect 19430 13696 19486 13705
rect 19430 13631 19486 13640
rect 19430 13560 19486 13569
rect 19430 13495 19486 13504
rect 18878 13359 18934 13368
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18748 12044 18828 12050
rect 18696 12038 18828 12044
rect 18708 12022 18828 12038
rect 18234 11792 18290 11801
rect 18052 11756 18104 11762
rect 18234 11727 18290 11736
rect 18052 11698 18104 11704
rect 18064 11354 18092 11698
rect 18708 11694 18736 12022
rect 18786 11792 18842 11801
rect 18786 11727 18842 11736
rect 18800 11694 18828 11727
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18156 11286 18184 11630
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10538 18000 10950
rect 18248 10606 18276 11630
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 18064 10130 18092 10542
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 18694 10160 18750 10169
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18064 9674 18092 10066
rect 17972 9646 18092 9674
rect 17972 9586 18000 9646
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17972 9042 18000 9522
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17972 8566 18000 8978
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 18064 8430 18092 9114
rect 18156 8922 18184 10134
rect 18694 10095 18750 10104
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18340 9722 18368 9862
rect 18432 9722 18460 9930
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18248 9489 18276 9590
rect 18234 9480 18290 9489
rect 18234 9415 18290 9424
rect 18248 9024 18276 9415
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18420 9036 18472 9042
rect 18248 8996 18420 9024
rect 18420 8978 18472 8984
rect 18156 8894 18276 8922
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18156 7954 18184 8774
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17880 7546 17908 7754
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17696 7449 17724 7482
rect 17682 7440 17738 7449
rect 17682 7375 17738 7384
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17684 4820 17736 4826
rect 17604 4780 17684 4808
rect 17684 4762 17736 4768
rect 17880 4282 17908 5102
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 3058 17080 3878
rect 17880 3534 17908 4218
rect 17972 4214 18000 7890
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 5302 18092 7686
rect 18248 7426 18276 8894
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18156 7398 18276 7426
rect 18708 7410 18736 10095
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18800 8945 18828 9454
rect 18786 8936 18842 8945
rect 18786 8871 18842 8880
rect 18788 8832 18840 8838
rect 18786 8800 18788 8809
rect 18840 8800 18842 8809
rect 18786 8735 18842 8744
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18696 7404 18748 7410
rect 18156 6662 18184 7398
rect 18696 7346 18748 7352
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18248 7002 18276 7278
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18524 6798 18552 6938
rect 18708 6866 18736 7346
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6186 18184 6598
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 18248 4690 18276 6190
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 18050 4176 18106 4185
rect 18050 4111 18052 4120
rect 18104 4111 18106 4120
rect 18052 4082 18104 4088
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17512 2446 17540 3334
rect 17604 3058 17632 3470
rect 18156 3194 18184 4558
rect 18234 4176 18290 4185
rect 18234 4111 18290 4120
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18248 3058 18276 4111
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18708 2650 18736 6190
rect 18800 3670 18828 7414
rect 18892 7206 18920 13126
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18984 9926 19012 11766
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18984 6458 19012 6734
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18892 5846 18920 6122
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18984 5234 19012 6394
rect 19076 5914 19104 10542
rect 19168 9110 19196 13330
rect 19352 12850 19380 13330
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19260 10606 19288 12582
rect 19352 12306 19380 12786
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19444 11506 19472 13495
rect 19352 11478 19472 11506
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19352 9994 19380 11478
rect 19536 11370 19564 14368
rect 19616 14350 19668 14356
rect 19614 13832 19670 13841
rect 19614 13767 19670 13776
rect 19628 13258 19656 13767
rect 19706 13560 19762 13569
rect 19706 13495 19762 13504
rect 19720 13258 19748 13495
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19720 12617 19748 12854
rect 19812 12782 19840 22714
rect 19892 22500 19944 22506
rect 19892 22442 19944 22448
rect 19904 22234 19932 22442
rect 19892 22228 19944 22234
rect 19892 22170 19944 22176
rect 19890 20496 19946 20505
rect 19890 20431 19946 20440
rect 19904 19786 19932 20431
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19904 19174 19932 19343
rect 19996 19310 20024 24142
rect 20180 23730 20208 24754
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 20088 22166 20116 22442
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 20180 21729 20208 23666
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20272 22166 20300 22510
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20166 21720 20222 21729
rect 20166 21655 20222 21664
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20088 20330 20116 21490
rect 20272 21457 20300 21626
rect 20258 21448 20314 21457
rect 20258 21383 20314 21392
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19904 18358 19932 18634
rect 19996 18426 20024 19246
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19904 16998 19932 17478
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19904 16674 19932 16934
rect 20088 16776 20116 20266
rect 20180 19281 20208 21082
rect 20166 19272 20222 19281
rect 20166 19207 20222 19216
rect 20180 17338 20208 19207
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20272 17241 20300 21286
rect 20456 20398 20484 24006
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18426 20484 19110
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20258 17232 20314 17241
rect 20258 17167 20314 17176
rect 20088 16748 20208 16776
rect 19904 16658 20116 16674
rect 19904 16652 20128 16658
rect 19904 16646 20076 16652
rect 20076 16594 20128 16600
rect 20076 15020 20128 15026
rect 20180 15008 20208 16748
rect 20350 16552 20406 16561
rect 20350 16487 20406 16496
rect 20364 16454 20392 16487
rect 20352 16448 20404 16454
rect 20444 16448 20496 16454
rect 20352 16390 20404 16396
rect 20442 16416 20444 16425
rect 20496 16416 20498 16425
rect 20442 16351 20498 16360
rect 20260 16040 20312 16046
rect 20258 16008 20260 16017
rect 20312 16008 20314 16017
rect 20258 15943 20314 15952
rect 20128 14980 20208 15008
rect 20076 14962 20128 14968
rect 20088 14657 20116 14962
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20074 14648 20130 14657
rect 20074 14583 20130 14592
rect 20088 13852 20116 14583
rect 20180 13977 20208 14758
rect 20166 13968 20222 13977
rect 20166 13903 20222 13912
rect 20088 13824 20208 13852
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19706 12608 19762 12617
rect 19706 12543 19762 12552
rect 19720 11898 19748 12543
rect 19812 12294 20024 12322
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19812 11778 19840 12294
rect 19996 12170 20024 12294
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19444 11342 19564 11370
rect 19720 11750 19840 11778
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19444 8498 19472 11342
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19628 10674 19656 11154
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19720 8430 19748 11750
rect 19904 11150 19932 12106
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19800 11144 19852 11150
rect 19798 11112 19800 11121
rect 19892 11144 19944 11150
rect 19852 11112 19854 11121
rect 19892 11086 19944 11092
rect 19798 11047 19854 11056
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19168 7410 19196 7890
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19168 6458 19196 7142
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19168 5098 19196 6394
rect 19260 6322 19288 8366
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 8022 19380 8230
rect 19720 8106 19748 8366
rect 19628 8078 19748 8106
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6458 19380 6802
rect 19628 6769 19656 8078
rect 19996 7993 20024 11834
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 20088 9722 20116 9930
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20088 8945 20116 9318
rect 20074 8936 20130 8945
rect 20074 8871 20130 8880
rect 20180 8514 20208 13824
rect 20272 10742 20300 15943
rect 20444 15904 20496 15910
rect 20364 15852 20444 15858
rect 20364 15846 20496 15852
rect 20364 15830 20484 15846
rect 20364 15094 20392 15830
rect 20444 15156 20496 15162
rect 20548 15144 20576 23598
rect 20824 23497 20852 24550
rect 20810 23488 20866 23497
rect 20810 23423 20866 23432
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20732 21690 20760 22102
rect 20824 21962 20852 22918
rect 20916 22522 20944 24890
rect 21008 24410 21036 25842
rect 21100 24818 21128 25842
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 20994 24168 21050 24177
rect 20994 24103 21050 24112
rect 21008 22642 21036 24103
rect 21100 23730 21128 24754
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21100 23186 21128 23666
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21192 23118 21220 26726
rect 21376 26586 21404 27406
rect 24228 27402 24256 29294
rect 25134 29200 25190 29800
rect 26422 29200 26478 29800
rect 27710 29200 27766 29800
rect 28998 29322 29054 29800
rect 29642 29322 29698 29800
rect 28644 29294 29054 29322
rect 25148 27538 25176 29200
rect 26238 28656 26294 28665
rect 26238 28591 26294 28600
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 25136 27532 25188 27538
rect 25136 27474 25188 27480
rect 24216 27396 24268 27402
rect 24216 27338 24268 27344
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21560 26382 21588 27270
rect 21652 26994 21680 27270
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 22664 27062 22692 27270
rect 22652 27056 22704 27062
rect 22652 26998 22704 27004
rect 21640 26988 21692 26994
rect 21640 26930 21692 26936
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21456 26308 21508 26314
rect 21456 26250 21508 26256
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21376 25362 21404 25638
rect 21468 25378 21496 26250
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 21560 25498 21588 25706
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21364 25356 21416 25362
rect 21468 25350 21588 25378
rect 21364 25298 21416 25304
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21284 23526 21312 24686
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21364 23520 21416 23526
rect 21468 23497 21496 24142
rect 21364 23462 21416 23468
rect 21454 23488 21510 23497
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21284 23118 21312 23258
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21088 23044 21140 23050
rect 21088 22986 21140 22992
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20916 22494 21036 22522
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20812 21956 20864 21962
rect 20812 21898 20864 21904
rect 20810 21720 20866 21729
rect 20720 21684 20772 21690
rect 20810 21655 20866 21664
rect 20720 21626 20772 21632
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20640 17542 20668 21082
rect 20824 20618 20852 21655
rect 20916 20754 20944 22374
rect 21008 22098 21036 22494
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 21100 21978 21128 22986
rect 21272 22568 21324 22574
rect 21376 22545 21404 23462
rect 21454 23423 21510 23432
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21272 22510 21324 22516
rect 21362 22536 21418 22545
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 21192 22166 21220 22442
rect 21180 22160 21232 22166
rect 21180 22102 21232 22108
rect 21100 21950 21220 21978
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21100 20874 21128 21830
rect 21192 20913 21220 21950
rect 21284 21729 21312 22510
rect 21362 22471 21418 22480
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21270 21720 21326 21729
rect 21270 21655 21326 21664
rect 21270 21584 21326 21593
rect 21270 21519 21326 21528
rect 21178 20904 21234 20913
rect 21088 20868 21140 20874
rect 21178 20839 21234 20848
rect 21088 20810 21140 20816
rect 20916 20726 21036 20754
rect 20824 20590 20944 20618
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19174 20760 20198
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20640 16810 20668 17274
rect 20732 16946 20760 17274
rect 20824 17202 20852 19314
rect 20916 18766 20944 20590
rect 21008 19446 21036 20726
rect 21284 19854 21312 21519
rect 21376 20777 21404 21898
rect 21362 20768 21418 20777
rect 21362 20703 21418 20712
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21376 20262 21404 20538
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20732 16918 20852 16946
rect 20824 16833 20852 16918
rect 20810 16824 20866 16833
rect 20640 16782 20760 16810
rect 20732 16726 20760 16782
rect 20810 16759 20866 16768
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20496 15116 20576 15144
rect 20444 15098 20496 15104
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20364 14346 20392 15030
rect 20548 14822 20576 15116
rect 20626 15056 20682 15065
rect 20626 14991 20628 15000
rect 20680 14991 20682 15000
rect 20628 14962 20680 14968
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20732 14385 20760 15370
rect 20718 14376 20774 14385
rect 20352 14340 20404 14346
rect 20718 14311 20774 14320
rect 20352 14282 20404 14288
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20456 12481 20484 13466
rect 20548 12753 20576 14214
rect 20640 14074 20668 14214
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20534 12744 20590 12753
rect 20534 12679 20590 12688
rect 20442 12472 20498 12481
rect 20442 12407 20498 12416
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20640 11218 20668 12242
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20442 10432 20498 10441
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20088 8486 20208 8514
rect 19982 7984 20038 7993
rect 19720 7942 19982 7970
rect 19720 7818 19748 7942
rect 19982 7919 20038 7928
rect 19996 7859 20024 7919
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19800 7812 19852 7818
rect 19800 7754 19852 7760
rect 19614 6760 19670 6769
rect 19614 6695 19670 6704
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19628 5914 19656 6190
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18892 3194 18920 3470
rect 19260 3398 19288 4490
rect 19352 4010 19380 5238
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19338 3768 19394 3777
rect 19338 3703 19394 3712
rect 19352 3670 19380 3703
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19444 3466 19472 5102
rect 19536 3534 19564 5646
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19628 3738 19656 4558
rect 19720 3942 19748 4694
rect 19812 4146 19840 7754
rect 20088 7002 20116 8486
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19982 6760 20038 6769
rect 19982 6695 19984 6704
rect 20036 6695 20038 6704
rect 19984 6666 20036 6672
rect 19890 6216 19946 6225
rect 20088 6202 20116 6938
rect 19890 6151 19946 6160
rect 19996 6174 20116 6202
rect 19904 5846 19932 6151
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19996 4554 20024 6174
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20088 5953 20116 6054
rect 20074 5944 20130 5953
rect 20074 5879 20130 5888
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20088 5098 20116 5646
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 20180 4146 20208 8298
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 19800 4004 19852 4010
rect 19800 3946 19852 3952
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18800 2446 18828 2790
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 12912 800 12940 2246
rect 13556 800 13584 2246
rect 14752 1306 14780 2246
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 14752 1278 14872 1306
rect 14844 800 14872 1278
rect 16132 800 16160 2382
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17420 800 17448 2246
rect 18696 1420 18748 1426
rect 18696 1362 18748 1368
rect 18708 800 18736 1362
rect 19352 800 19380 2858
rect 19536 2650 19564 2926
rect 19720 2854 19748 3878
rect 19812 3126 19840 3946
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 20272 2854 20300 9522
rect 20364 8634 20392 10406
rect 20442 10367 20498 10376
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20364 8129 20392 8434
rect 20350 8120 20406 8129
rect 20350 8055 20406 8064
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20364 6390 20392 6734
rect 20456 6730 20484 10367
rect 20548 10169 20576 10542
rect 20534 10160 20590 10169
rect 20640 10130 20668 11154
rect 20732 10606 20760 13806
rect 20824 13569 20852 16759
rect 20916 14006 20944 18702
rect 21272 18692 21324 18698
rect 21192 18652 21272 18680
rect 21192 17542 21220 18652
rect 21272 18634 21324 18640
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21100 16114 21128 17138
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20810 13560 20866 13569
rect 20810 13495 20866 13504
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20824 13297 20852 13398
rect 20810 13288 20866 13297
rect 20810 13223 20866 13232
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12434 20852 12650
rect 20824 12406 20944 12434
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20534 10095 20590 10104
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20640 9704 20668 10066
rect 20640 9676 20760 9704
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20548 8838 20576 9522
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 8838 20668 9318
rect 20732 9042 20760 9676
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8650 20668 8774
rect 20548 8622 20668 8650
rect 20732 8634 20760 8978
rect 20824 8974 20852 11494
rect 20916 9897 20944 12406
rect 21008 12306 21036 16050
rect 21100 13938 21128 16050
rect 21192 14618 21220 17478
rect 21376 17338 21404 19654
rect 21468 19378 21496 23122
rect 21560 19990 21588 25350
rect 22112 25265 22140 25638
rect 22098 25256 22154 25265
rect 22098 25191 22154 25200
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22204 24410 22232 24686
rect 22572 24614 22600 26726
rect 22664 26586 22692 26862
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22756 26382 22784 26726
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22664 25401 22692 25774
rect 22650 25392 22706 25401
rect 22650 25327 22706 25336
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24886 22784 25230
rect 22744 24880 22796 24886
rect 22744 24822 22796 24828
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22374 24032 22430 24041
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 22204 23662 22232 24006
rect 22374 23967 22430 23976
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 21185 21680 23054
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 22204 21622 22232 22374
rect 22388 21962 22416 23967
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22468 23792 22520 23798
rect 22468 23734 22520 23740
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 21638 21176 21694 21185
rect 21638 21111 21694 21120
rect 21824 21004 21876 21010
rect 21652 20964 21824 20992
rect 21652 20602 21680 20964
rect 21824 20946 21876 20952
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21560 19446 21588 19926
rect 21652 19922 21680 20402
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 21914 19952 21970 19961
rect 21640 19916 21692 19922
rect 22020 19922 22048 20334
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 21914 19887 21970 19896
rect 22008 19916 22060 19922
rect 21640 19858 21692 19864
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21652 19378 21680 19858
rect 21928 19786 21956 19887
rect 22008 19858 22060 19864
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21652 17746 21680 19314
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 22204 18408 22232 19994
rect 22020 18380 22232 18408
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21468 16794 21496 17274
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21192 13734 21220 14282
rect 21284 14074 21312 16458
rect 21560 16454 21588 17546
rect 21652 17202 21680 17682
rect 22020 17610 22048 18380
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21652 16658 21680 17138
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21836 16522 21864 17274
rect 22296 17134 22324 21286
rect 22388 19961 22416 21898
rect 22480 20602 22508 23734
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22572 22030 22600 22578
rect 22560 22024 22612 22030
rect 22664 22012 22692 23802
rect 22744 22704 22796 22710
rect 22742 22672 22744 22681
rect 22796 22672 22798 22681
rect 22742 22607 22798 22616
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22756 22166 22784 22374
rect 22744 22160 22796 22166
rect 22744 22102 22796 22108
rect 22664 21984 22784 22012
rect 22560 21966 22612 21972
rect 22572 21554 22600 21966
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22374 19952 22430 19961
rect 22374 19887 22430 19896
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 22480 19514 22508 19722
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22756 19334 22784 21984
rect 22848 21010 22876 26182
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 22940 24342 22968 24618
rect 22928 24336 22980 24342
rect 22928 24278 22980 24284
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 22642 22968 23462
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 22926 22128 22982 22137
rect 22926 22063 22928 22072
rect 22980 22063 22982 22072
rect 22928 22034 22980 22040
rect 23032 21729 23060 26930
rect 23400 26858 23428 27270
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 23124 24206 23152 24278
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23018 21720 23074 21729
rect 23018 21655 23074 21664
rect 23032 21622 23060 21655
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 23032 21457 23060 21558
rect 23018 21448 23074 21457
rect 23018 21383 23074 21392
rect 23124 21146 23152 24142
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22848 19825 22876 20742
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22834 19816 22890 19825
rect 22834 19751 22890 19760
rect 23032 19514 23060 20198
rect 23124 20058 23152 20266
rect 23112 20052 23164 20058
rect 23112 19994 23164 20000
rect 23216 19768 23244 25094
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23308 23798 23336 24686
rect 23400 24274 23428 25638
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23584 24206 23612 26318
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23296 23792 23348 23798
rect 23294 23760 23296 23769
rect 23348 23760 23350 23769
rect 23294 23695 23350 23704
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 20618 23336 22918
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23400 21486 23428 21898
rect 23492 21622 23520 23530
rect 23768 23118 23796 25298
rect 23860 24818 23888 26726
rect 24124 25832 24176 25838
rect 24124 25774 24176 25780
rect 23940 24880 23992 24886
rect 23940 24822 23992 24828
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23572 22568 23624 22574
rect 23676 22545 23704 22986
rect 23860 22794 23888 24142
rect 23768 22766 23888 22794
rect 23572 22510 23624 22516
rect 23662 22536 23718 22545
rect 23584 22234 23612 22510
rect 23662 22471 23718 22480
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23768 22094 23796 22766
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23584 22066 23796 22094
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23584 21486 23612 22066
rect 23754 21992 23810 22001
rect 23754 21927 23810 21936
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23570 21176 23626 21185
rect 23570 21111 23626 21120
rect 23308 20590 23520 20618
rect 23492 20534 23520 20590
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23584 20398 23612 21111
rect 23572 20392 23624 20398
rect 23492 20352 23572 20380
rect 23296 19780 23348 19786
rect 23216 19740 23296 19768
rect 23296 19722 23348 19728
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22756 19306 22968 19334
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22848 18970 22876 19110
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22374 17912 22430 17921
rect 22374 17847 22430 17856
rect 22388 17610 22416 17847
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22374 17232 22430 17241
rect 22374 17167 22430 17176
rect 22284 17128 22336 17134
rect 22006 17096 22062 17105
rect 21916 17060 21968 17066
rect 22284 17070 22336 17076
rect 22006 17031 22008 17040
rect 21916 17002 21968 17008
rect 22060 17031 22062 17040
rect 22008 17002 22060 17008
rect 21928 16658 21956 17002
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22388 16522 22416 17167
rect 22468 17128 22520 17134
rect 22520 17088 22784 17116
rect 22468 17070 22520 17076
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22466 16688 22522 16697
rect 22572 16658 22600 16934
rect 22466 16623 22468 16632
rect 22520 16623 22522 16632
rect 22560 16652 22612 16658
rect 22468 16594 22520 16600
rect 22560 16594 22612 16600
rect 22466 16552 22522 16561
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 22376 16516 22428 16522
rect 22466 16487 22522 16496
rect 22376 16458 22428 16464
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21652 16130 21680 16458
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 21928 16153 21956 16186
rect 22480 16182 22508 16487
rect 22468 16176 22520 16182
rect 21914 16144 21970 16153
rect 21652 16102 21864 16130
rect 21732 15972 21784 15978
rect 21732 15914 21784 15920
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21546 15736 21602 15745
rect 21546 15671 21548 15680
rect 21600 15671 21602 15680
rect 21548 15642 21600 15648
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21376 14929 21404 14962
rect 21362 14920 21418 14929
rect 21362 14855 21418 14864
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 20902 9888 20958 9897
rect 20902 9823 20958 9832
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20720 8628 20772 8634
rect 20548 7449 20576 8622
rect 20720 8570 20772 8576
rect 20718 8528 20774 8537
rect 20824 8498 20852 8910
rect 20718 8463 20720 8472
rect 20772 8463 20774 8472
rect 20812 8492 20864 8498
rect 20720 8434 20772 8440
rect 20812 8434 20864 8440
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20626 7848 20682 7857
rect 20626 7783 20682 7792
rect 20534 7440 20590 7449
rect 20534 7375 20590 7384
rect 20640 6866 20668 7783
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20444 6724 20496 6730
rect 20496 6684 20576 6712
rect 20444 6666 20496 6672
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20352 6384 20404 6390
rect 20352 6326 20404 6332
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20364 5710 20392 5782
rect 20456 5710 20484 6394
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20548 5556 20576 6684
rect 20628 6316 20680 6322
rect 20732 6304 20760 8298
rect 20824 6730 20852 8298
rect 20916 7546 20944 9658
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20680 6276 20760 6304
rect 20812 6316 20864 6322
rect 20628 6258 20680 6264
rect 20812 6258 20864 6264
rect 20824 5846 20852 6258
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20916 5642 20944 7482
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20548 5528 20760 5556
rect 20732 5098 20760 5528
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4758 20392 4966
rect 20824 4826 20852 5102
rect 21008 4826 21036 12106
rect 21100 11694 21128 13670
rect 21178 13560 21234 13569
rect 21178 13495 21234 13504
rect 21192 13462 21220 13495
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21192 13190 21220 13398
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21284 12209 21312 13874
rect 21362 13696 21418 13705
rect 21362 13631 21418 13640
rect 21270 12200 21326 12209
rect 21270 12135 21326 12144
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 21178 11248 21234 11257
rect 21178 11183 21234 11192
rect 21088 11144 21140 11150
rect 21086 11112 21088 11121
rect 21140 11112 21142 11121
rect 21192 11082 21220 11183
rect 21086 11047 21142 11056
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21192 10033 21220 10746
rect 21284 10674 21312 12135
rect 21376 10810 21404 13631
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21468 10554 21496 14282
rect 21560 13258 21588 15302
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21560 12374 21588 13194
rect 21652 12986 21680 15846
rect 21744 15366 21772 15914
rect 21836 15586 21864 16102
rect 22468 16118 22520 16124
rect 22558 16144 22614 16153
rect 21914 16079 21970 16088
rect 22558 16079 22614 16088
rect 22572 16046 22600 16079
rect 22100 16040 22152 16046
rect 22468 16040 22520 16046
rect 22100 15982 22152 15988
rect 22466 16008 22468 16017
rect 22560 16040 22612 16046
rect 22520 16008 22522 16017
rect 22112 15706 22140 15982
rect 22560 15982 22612 15988
rect 22466 15943 22522 15952
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 15745 22232 15846
rect 22190 15736 22246 15745
rect 22100 15700 22152 15706
rect 22190 15671 22246 15680
rect 22284 15700 22336 15706
rect 22100 15642 22152 15648
rect 22284 15642 22336 15648
rect 21836 15558 21956 15586
rect 21822 15464 21878 15473
rect 21928 15434 21956 15558
rect 21822 15399 21824 15408
rect 21876 15399 21878 15408
rect 21916 15428 21968 15434
rect 21824 15370 21876 15376
rect 21916 15370 21968 15376
rect 21732 15360 21784 15366
rect 22112 15348 22140 15642
rect 22296 15473 22324 15642
rect 22282 15464 22338 15473
rect 22282 15399 22338 15408
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22112 15320 22232 15348
rect 21732 15302 21784 15308
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 22204 15026 22232 15320
rect 22388 15162 22416 15370
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22020 13394 22048 13806
rect 22098 13424 22154 13433
rect 22008 13388 22060 13394
rect 22098 13359 22100 13368
rect 22008 13330 22060 13336
rect 22152 13359 22154 13368
rect 22100 13330 22152 13336
rect 22190 13288 22246 13297
rect 22190 13223 22246 13232
rect 22204 13190 22232 13223
rect 22296 13190 22324 14826
rect 22652 14544 22704 14550
rect 22652 14486 22704 14492
rect 22558 14376 22614 14385
rect 22558 14311 22614 14320
rect 22374 13832 22430 13841
rect 22374 13767 22430 13776
rect 22388 13734 22416 13767
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 22284 12912 22336 12918
rect 22282 12880 22284 12889
rect 22336 12880 22338 12889
rect 22282 12815 22338 12824
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22204 12434 22232 12718
rect 22572 12442 22600 14311
rect 22560 12436 22612 12442
rect 22204 12406 22324 12434
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 22296 12238 22324 12406
rect 22560 12378 22612 12384
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11558 21588 12106
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 22192 11824 22244 11830
rect 22190 11792 22192 11801
rect 22244 11792 22246 11801
rect 22008 11756 22060 11762
rect 22190 11727 22246 11736
rect 22008 11698 22060 11704
rect 22020 11642 22048 11698
rect 22296 11642 22324 12174
rect 22664 12170 22692 14486
rect 22756 13569 22784 17088
rect 22848 15162 22876 18634
rect 22940 15570 22968 19306
rect 23204 19304 23256 19310
rect 23202 19272 23204 19281
rect 23296 19304 23348 19310
rect 23256 19272 23258 19281
rect 23296 19246 23348 19252
rect 23202 19207 23258 19216
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23124 16504 23152 18566
rect 23216 18426 23244 19110
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23308 18154 23336 19246
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23400 18329 23428 18838
rect 23386 18320 23442 18329
rect 23386 18255 23442 18264
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 16794 23428 17478
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23204 16516 23256 16522
rect 23124 16476 23204 16504
rect 23204 16458 23256 16464
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22742 13560 22798 13569
rect 22742 13495 22798 13504
rect 22848 12918 22876 14214
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 22926 12880 22982 12889
rect 22652 12164 22704 12170
rect 22652 12106 22704 12112
rect 22376 11824 22428 11830
rect 22558 11792 22614 11801
rect 22428 11772 22508 11778
rect 22376 11766 22508 11772
rect 22388 11750 22508 11766
rect 22020 11614 22324 11642
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 22296 11218 22324 11614
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 21640 11076 21692 11082
rect 21560 11036 21640 11064
rect 21560 10690 21588 11036
rect 21640 11018 21692 11024
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 22190 10840 22246 10849
rect 22190 10775 22246 10784
rect 21560 10662 21680 10690
rect 21376 10526 21496 10554
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21178 10024 21234 10033
rect 21088 9988 21140 9994
rect 21178 9959 21234 9968
rect 21088 9930 21140 9936
rect 21100 5370 21128 9930
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 5846 21220 8842
rect 21284 6866 21312 9658
rect 21376 9518 21404 10526
rect 21560 9926 21588 10542
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21468 9382 21496 9862
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21652 9194 21680 10662
rect 22204 10554 22232 10775
rect 22296 10742 22324 11154
rect 22284 10736 22336 10742
rect 22376 10736 22428 10742
rect 22284 10678 22336 10684
rect 22374 10704 22376 10713
rect 22428 10704 22430 10713
rect 22296 10588 22324 10678
rect 22374 10639 22430 10648
rect 22296 10560 22416 10588
rect 22112 10538 22232 10554
rect 22100 10532 22232 10538
rect 22152 10526 22232 10532
rect 22100 10474 22152 10480
rect 22098 10296 22154 10305
rect 22388 10282 22416 10560
rect 22098 10231 22100 10240
rect 22152 10231 22154 10240
rect 22296 10254 22416 10282
rect 22100 10202 22152 10208
rect 22190 10160 22246 10169
rect 22190 10095 22246 10104
rect 22204 9994 22232 10095
rect 22296 10062 22324 10254
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 22296 9586 22324 9998
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22480 9518 22508 11750
rect 22558 11727 22614 11736
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 21560 9166 21680 9194
rect 21364 9036 21416 9042
rect 21416 8996 21496 9024
rect 21364 8978 21416 8984
rect 21468 8566 21496 8996
rect 21456 8560 21508 8566
rect 21362 8528 21418 8537
rect 21456 8502 21508 8508
rect 21362 8463 21364 8472
rect 21416 8463 21418 8472
rect 21364 8434 21416 8440
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21468 8106 21496 8366
rect 21560 8294 21588 9166
rect 21638 9072 21694 9081
rect 22480 9042 22508 9454
rect 21638 9007 21640 9016
rect 21692 9007 21694 9016
rect 22468 9036 22520 9042
rect 21640 8978 21692 8984
rect 22468 8978 22520 8984
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21468 8078 21588 8106
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21362 7440 21418 7449
rect 21362 7375 21364 7384
rect 21416 7375 21418 7384
rect 21364 7346 21416 7352
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20456 3534 20484 3878
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20548 2650 20576 4626
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 3194 20852 4558
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20916 3777 20944 4082
rect 20902 3768 20958 3777
rect 20902 3703 20958 3712
rect 21192 3670 21220 5510
rect 21284 5370 21312 6802
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6254 21404 6598
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21468 3738 21496 7958
rect 21560 6322 21588 8078
rect 21652 7954 21680 8570
rect 22020 8498 22048 8570
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21652 7342 21680 7482
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 22204 6866 22232 8502
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22296 7857 22324 7890
rect 22282 7848 22338 7857
rect 22282 7783 22338 7792
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22296 6730 22324 7686
rect 22388 6769 22416 8910
rect 22572 8906 22600 11727
rect 22664 11354 22692 12106
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22664 9897 22692 10066
rect 22650 9888 22706 9897
rect 22650 9823 22706 9832
rect 22650 9072 22706 9081
rect 22650 9007 22706 9016
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22664 8430 22692 9007
rect 22848 8974 22876 12854
rect 22926 12815 22982 12824
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22652 8424 22704 8430
rect 22572 8384 22652 8412
rect 22466 8120 22522 8129
rect 22466 8055 22522 8064
rect 22374 6760 22430 6769
rect 22284 6724 22336 6730
rect 22374 6695 22430 6704
rect 22284 6666 22336 6672
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 22284 5704 22336 5710
rect 22480 5692 22508 8055
rect 22572 6338 22600 8384
rect 22652 8366 22704 8372
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 6866 22692 7346
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22572 6310 22692 6338
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22572 5778 22600 6190
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22336 5664 22508 5692
rect 22284 5646 22336 5652
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 22558 5264 22614 5273
rect 22558 5199 22560 5208
rect 22612 5199 22614 5208
rect 22560 5170 22612 5176
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22388 4826 22416 4966
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21640 4004 21692 4010
rect 21640 3946 21692 3952
rect 21652 3738 21680 3946
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20810 3088 20866 3097
rect 20628 3052 20680 3058
rect 20810 3023 20812 3032
rect 20628 2994 20680 3000
rect 20864 3023 20866 3032
rect 20812 2994 20864 3000
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20548 1426 20576 2382
rect 20536 1420 20588 1426
rect 20536 1362 20588 1368
rect 20640 800 20668 2994
rect 21560 2990 21588 3606
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 22204 3194 22232 4490
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 21548 2984 21600 2990
rect 21548 2926 21600 2932
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21468 2446 21496 2858
rect 22296 2582 22324 4558
rect 22664 4185 22692 6310
rect 22756 5642 22784 7414
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22756 4282 22784 5102
rect 22848 4758 22876 8502
rect 22940 7546 22968 12815
rect 23032 11898 23060 15574
rect 23492 15162 23520 20352
rect 23572 20334 23624 20340
rect 23768 19378 23796 21927
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23584 18086 23612 18362
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23112 15088 23164 15094
rect 23110 15056 23112 15065
rect 23164 15056 23166 15065
rect 23110 14991 23166 15000
rect 23294 14784 23350 14793
rect 23294 14719 23350 14728
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23112 13320 23164 13326
rect 23216 13297 23244 13398
rect 23112 13262 23164 13268
rect 23202 13288 23258 13297
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 23018 11248 23074 11257
rect 23018 11183 23020 11192
rect 23072 11183 23074 11192
rect 23020 11154 23072 11160
rect 23124 9110 23152 13262
rect 23202 13223 23258 13232
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 23216 10130 23244 12582
rect 23308 11830 23336 14719
rect 23478 14648 23534 14657
rect 23584 14618 23612 17546
rect 23860 17218 23888 22646
rect 23952 21026 23980 24822
rect 24136 23866 24164 25774
rect 24504 25294 24532 26726
rect 24952 26240 25004 26246
rect 24952 26182 25004 26188
rect 24964 25906 24992 26182
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24584 24608 24636 24614
rect 24584 24550 24636 24556
rect 24596 24274 24624 24550
rect 24780 24410 24808 25706
rect 25056 25378 25084 27270
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 24964 25350 25084 25378
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24584 24268 24636 24274
rect 24584 24210 24636 24216
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24676 23792 24728 23798
rect 24676 23734 24728 23740
rect 24032 23588 24084 23594
rect 24032 23530 24084 23536
rect 24044 21350 24072 23530
rect 24688 23322 24716 23734
rect 24964 23662 24992 25350
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 25504 25288 25556 25294
rect 25504 25230 25556 25236
rect 25056 23730 25084 25230
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25148 23730 25176 25094
rect 25424 24886 25452 25230
rect 25412 24880 25464 24886
rect 25412 24822 25464 24828
rect 25516 24682 25544 25230
rect 25504 24676 25556 24682
rect 25504 24618 25556 24624
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25228 24064 25280 24070
rect 25320 24064 25372 24070
rect 25228 24006 25280 24012
rect 25318 24032 25320 24041
rect 25372 24032 25374 24041
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 24952 23656 25004 23662
rect 24952 23598 25004 23604
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24136 21146 24164 21966
rect 24216 21956 24268 21962
rect 24216 21898 24268 21904
rect 24228 21418 24256 21898
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 23952 20998 24164 21026
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 23676 17190 23888 17218
rect 23478 14583 23534 14592
rect 23572 14612 23624 14618
rect 23492 14414 23520 14583
rect 23572 14554 23624 14560
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23570 13968 23626 13977
rect 23570 13903 23626 13912
rect 23584 13394 23612 13903
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23676 12374 23704 17190
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23768 12434 23796 16594
rect 23952 15910 23980 18158
rect 24044 16998 24072 20878
rect 24136 17134 24164 20998
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 24228 18193 24256 18634
rect 24214 18184 24270 18193
rect 24214 18119 24270 18128
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24136 16697 24164 17070
rect 24122 16688 24178 16697
rect 24122 16623 24178 16632
rect 24228 16538 24256 18119
rect 24412 17882 24440 22170
rect 24504 21622 24532 23054
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 21622 24624 21830
rect 24688 21690 24716 22374
rect 24964 22094 24992 23122
rect 24872 22066 24992 22094
rect 24872 21690 24900 22066
rect 25056 21894 25084 23666
rect 25240 23610 25268 24006
rect 25318 23967 25374 23976
rect 25148 23582 25268 23610
rect 25516 23610 25544 24074
rect 25608 23798 25636 27270
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 25872 26512 25924 26518
rect 25872 26454 25924 26460
rect 25688 25696 25740 25702
rect 25688 25638 25740 25644
rect 25700 25430 25728 25638
rect 25688 25424 25740 25430
rect 25688 25366 25740 25372
rect 25884 24818 25912 26454
rect 25976 26450 26004 26726
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 26068 24750 26096 26726
rect 26252 26382 26280 28591
rect 26436 27470 26464 29200
rect 27528 27668 27580 27674
rect 27528 27610 27580 27616
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27160 27328 27212 27334
rect 27160 27270 27212 27276
rect 27172 27062 27200 27270
rect 27160 27056 27212 27062
rect 27160 26998 27212 27004
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26528 26314 26556 26930
rect 27356 26586 27384 26930
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 26884 26376 26936 26382
rect 26884 26318 26936 26324
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 26516 26308 26568 26314
rect 26516 26250 26568 26256
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25700 23866 25728 24142
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25516 23582 25636 23610
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24492 21616 24544 21622
rect 24492 21558 24544 21564
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 24688 21554 24716 21626
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24504 19786 24532 21422
rect 24688 20262 24716 21490
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24780 21010 24808 21422
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24688 19922 24716 20198
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24492 19780 24544 19786
rect 24492 19722 24544 19728
rect 24688 19378 24716 19858
rect 24676 19372 24728 19378
rect 24596 19332 24676 19360
rect 24596 18834 24624 19332
rect 24676 19314 24728 19320
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 24596 18086 24624 18770
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24320 17542 24348 17818
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24136 16510 24256 16538
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 24044 14074 24072 15982
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 24136 13954 24164 16510
rect 24412 16232 24440 17818
rect 24596 17746 24624 18022
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24504 17134 24532 17682
rect 24596 17202 24624 17682
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24596 16658 24624 17138
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24492 16244 24544 16250
rect 24412 16204 24492 16232
rect 24492 16186 24544 16192
rect 24596 16182 24624 16594
rect 24584 16176 24636 16182
rect 24584 16118 24636 16124
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 23952 13926 24164 13954
rect 23768 12406 23888 12434
rect 23664 12368 23716 12374
rect 23716 12316 23796 12322
rect 23664 12310 23796 12316
rect 23676 12294 23796 12310
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23492 10674 23520 12038
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23584 10441 23612 12038
rect 23676 11354 23704 12174
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23570 10432 23626 10441
rect 23570 10367 23626 10376
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23768 9194 23796 12294
rect 23860 11830 23888 12406
rect 23952 11898 23980 13926
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 23952 11082 23980 11630
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 24044 10266 24072 11630
rect 24136 10742 24164 12922
rect 24228 12918 24256 15642
rect 24596 15638 24624 16118
rect 24780 15910 24808 20946
rect 25056 20482 25084 21830
rect 24872 20454 25084 20482
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24872 14958 24900 20454
rect 25044 20392 25096 20398
rect 25044 20334 25096 20340
rect 25056 19310 25084 20334
rect 25148 19446 25176 23582
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25608 22710 25636 23582
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25872 22976 25924 22982
rect 25872 22918 25924 22924
rect 25700 22778 25728 22918
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 25596 22704 25648 22710
rect 25596 22646 25648 22652
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25332 21593 25360 21898
rect 25318 21584 25374 21593
rect 25318 21519 25374 21528
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25136 19440 25188 19446
rect 25136 19382 25188 19388
rect 25044 19304 25096 19310
rect 24950 19272 25006 19281
rect 25044 19246 25096 19252
rect 24950 19207 25006 19216
rect 24964 19122 24992 19207
rect 24964 19094 25084 19122
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 24964 17649 24992 17750
rect 24950 17640 25006 17649
rect 24950 17575 25006 17584
rect 25056 15162 25084 19094
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25148 17270 25176 18362
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 25148 16182 25176 16458
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 25134 15872 25190 15881
rect 25134 15807 25190 15816
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 24952 15088 25004 15094
rect 25004 15036 25084 15042
rect 24952 15030 25084 15036
rect 24964 15014 25084 15030
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24596 14414 24624 14894
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24320 12986 24348 13126
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12186 24348 12786
rect 24400 12232 24452 12238
rect 24228 12158 24348 12186
rect 24398 12200 24400 12209
rect 24452 12200 24454 12209
rect 24228 11014 24256 12158
rect 24398 12135 24454 12144
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24214 10840 24270 10849
rect 24214 10775 24270 10784
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 24228 10674 24256 10775
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24136 10169 24164 10542
rect 24320 10538 24348 12038
rect 24504 11354 24532 13942
rect 24596 13870 24624 14350
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24596 12850 24624 13806
rect 24780 13530 24808 14282
rect 24872 14006 24900 14758
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24964 13258 24992 14418
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 25056 13138 25084 15014
rect 25148 14464 25176 15807
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25148 14436 25268 14464
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 24964 13110 25084 13138
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24780 12850 24808 12922
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24596 11762 24624 12786
rect 24858 12472 24914 12481
rect 24858 12407 24914 12416
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24400 11280 24452 11286
rect 24400 11222 24452 11228
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24228 10305 24256 10406
rect 24214 10296 24270 10305
rect 24214 10231 24270 10240
rect 24216 10192 24268 10198
rect 24122 10160 24178 10169
rect 24216 10134 24268 10140
rect 24122 10095 24178 10104
rect 23768 9166 23980 9194
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23202 8120 23258 8129
rect 23202 8055 23258 8064
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23216 7410 23244 8055
rect 23308 7954 23336 8910
rect 23754 8392 23810 8401
rect 23754 8327 23756 8336
rect 23808 8327 23810 8336
rect 23756 8298 23808 8304
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 8090 23428 8230
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23768 7886 23796 8026
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 22940 5098 22968 6190
rect 23124 5914 23152 6666
rect 23204 6384 23256 6390
rect 23204 6326 23256 6332
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23110 5808 23166 5817
rect 23110 5743 23166 5752
rect 23124 5710 23152 5743
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23020 5296 23072 5302
rect 23020 5238 23072 5244
rect 22928 5092 22980 5098
rect 22928 5034 22980 5040
rect 23032 4826 23060 5238
rect 23216 4826 23244 6326
rect 23308 5710 23336 6802
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22650 4176 22706 4185
rect 22376 4140 22428 4146
rect 22650 4111 22706 4120
rect 22376 4082 22428 4088
rect 22388 3738 22416 4082
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22664 2650 22692 4014
rect 23308 3534 23336 5646
rect 23400 4146 23428 6666
rect 23492 6322 23520 7346
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23584 3738 23612 7278
rect 23754 6896 23810 6905
rect 23754 6831 23756 6840
rect 23808 6831 23810 6840
rect 23756 6802 23808 6808
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 23676 6118 23704 6326
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23676 5234 23704 5510
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23860 4622 23888 8978
rect 23952 4706 23980 9166
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24136 7954 24164 8570
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24136 7410 24164 7890
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 23952 4678 24072 4706
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23952 4282 23980 4558
rect 23940 4276 23992 4282
rect 23940 4218 23992 4224
rect 24044 3942 24072 4678
rect 24136 4078 24164 7210
rect 24228 5817 24256 10134
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24320 9178 24348 9318
rect 24308 9172 24360 9178
rect 24308 9114 24360 9120
rect 24412 7342 24440 11222
rect 24596 10674 24624 11698
rect 24780 11150 24808 12174
rect 24872 11694 24900 12407
rect 24964 11694 24992 13110
rect 25042 12608 25098 12617
rect 25042 12543 25098 12552
rect 25056 12306 25084 12543
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 10130 24624 10610
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24504 6866 24532 10066
rect 24596 9586 24624 10066
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24596 9024 24624 9522
rect 24676 9036 24728 9042
rect 24596 8996 24676 9024
rect 24596 8430 24624 8996
rect 24676 8978 24728 8984
rect 24780 8974 24808 11086
rect 25148 9738 25176 14282
rect 25240 14074 25268 14436
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25608 13394 25636 21966
rect 25700 20505 25728 22374
rect 25884 21729 25912 22918
rect 25870 21720 25926 21729
rect 25870 21655 25926 21664
rect 25780 21412 25832 21418
rect 25780 21354 25832 21360
rect 25686 20496 25742 20505
rect 25686 20431 25742 20440
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25240 12646 25268 13330
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25596 12640 25648 12646
rect 25596 12582 25648 12588
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 24964 9710 25176 9738
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24872 9081 24900 9114
rect 24858 9072 24914 9081
rect 24858 9007 24914 9016
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24766 8392 24822 8401
rect 24596 7954 24624 8366
rect 24964 8378 24992 9710
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24822 8350 24992 8378
rect 24766 8327 24822 8336
rect 24860 8016 24912 8022
rect 24860 7958 24912 7964
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24596 6798 24624 7890
rect 24872 7478 24900 7958
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24872 6390 24900 7278
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24688 5953 24716 6190
rect 24674 5944 24730 5953
rect 24674 5879 24730 5888
rect 24688 5846 24716 5879
rect 24676 5840 24728 5846
rect 24214 5808 24270 5817
rect 24676 5782 24728 5788
rect 24214 5743 24270 5752
rect 24780 5710 24808 6258
rect 25056 5914 25084 9590
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25318 8936 25374 8945
rect 25136 8900 25188 8906
rect 25318 8871 25374 8880
rect 25136 8842 25188 8848
rect 25148 6390 25176 8842
rect 25332 8566 25360 8871
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25410 6896 25466 6905
rect 25410 6831 25466 6840
rect 25424 6730 25452 6831
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23400 3194 23428 3334
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 24596 2650 24624 5646
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24688 4282 24716 5102
rect 24964 4758 24992 5850
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 25042 4040 25098 4049
rect 25042 3975 25098 3984
rect 25056 3738 25084 3975
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 25148 3194 25176 4558
rect 25608 4010 25636 12582
rect 25686 11656 25742 11665
rect 25686 11591 25742 11600
rect 25700 6254 25728 11591
rect 25792 10266 25820 21354
rect 25884 18358 25912 21655
rect 25976 20058 26004 24550
rect 26068 24274 26096 24550
rect 26056 24268 26108 24274
rect 26056 24210 26108 24216
rect 26424 24200 26476 24206
rect 26424 24142 26476 24148
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 26068 19990 26096 23666
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26252 23118 26280 23462
rect 26436 23322 26464 24142
rect 26424 23316 26476 23322
rect 26424 23258 26476 23264
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26252 21554 26280 21966
rect 26528 21962 26556 26250
rect 26700 26240 26752 26246
rect 26700 26182 26752 26188
rect 26712 25906 26740 26182
rect 26896 25945 26924 26318
rect 26882 25936 26938 25945
rect 26700 25900 26752 25906
rect 26882 25871 26938 25880
rect 26700 25842 26752 25848
rect 26792 25288 26844 25294
rect 26792 25230 26844 25236
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 26252 21010 26280 21490
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26056 19984 26108 19990
rect 26056 19926 26108 19932
rect 26436 19514 26464 20538
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 26252 17610 26280 18906
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26436 16130 26464 19450
rect 26528 18902 26556 21898
rect 26516 18896 26568 18902
rect 26516 18838 26568 18844
rect 26620 16658 26648 23462
rect 26700 19780 26752 19786
rect 26700 19722 26752 19728
rect 26712 17134 26740 19722
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26344 16102 26464 16130
rect 26344 15706 26372 16102
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 26332 15700 26384 15706
rect 26332 15642 26384 15648
rect 25872 15428 25924 15434
rect 25872 15370 25924 15376
rect 25884 12170 25912 15370
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 25964 13796 26016 13802
rect 25964 13738 26016 13744
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25884 9897 25912 9930
rect 25870 9888 25926 9897
rect 25870 9823 25926 9832
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25792 4026 25820 9454
rect 25976 7818 26004 13738
rect 26068 11121 26096 14418
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26160 13870 26188 14282
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 26160 13394 26188 13466
rect 26252 13462 26280 14758
rect 26330 13696 26386 13705
rect 26330 13631 26386 13640
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26344 13394 26372 13631
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26160 11218 26188 13330
rect 26344 12986 26372 13330
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26344 12434 26372 12922
rect 26436 12646 26464 15982
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26620 14521 26648 14894
rect 26606 14512 26662 14521
rect 26606 14447 26662 14456
rect 26712 14090 26740 15846
rect 26804 14618 26832 25230
rect 27264 24410 27292 26318
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27356 24818 27384 25638
rect 27448 25498 27476 27406
rect 27540 27130 27568 27610
rect 27724 27606 27752 29200
rect 27712 27600 27764 27606
rect 27712 27542 27764 27548
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27540 26042 27568 26930
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27436 25492 27488 25498
rect 27436 25434 27488 25440
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27540 24585 27568 25774
rect 27526 24576 27582 24585
rect 27526 24511 27582 24520
rect 27724 24410 27752 25842
rect 27908 25498 27936 26862
rect 28644 26586 28672 29294
rect 28998 29200 29054 29294
rect 29288 29294 29698 29322
rect 29288 27674 29316 29294
rect 29642 29200 29698 29294
rect 29276 27668 29328 27674
rect 29276 27610 29328 27616
rect 29918 27296 29974 27305
rect 28734 27228 29042 27237
rect 29918 27231 29974 27240
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 29932 27130 29960 27231
rect 29920 27124 29972 27130
rect 29920 27066 29972 27072
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 27712 24404 27764 24410
rect 27712 24346 27764 24352
rect 27710 24304 27766 24313
rect 27710 24239 27766 24248
rect 27158 22672 27214 22681
rect 27158 22607 27214 22616
rect 27172 21554 27200 22607
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27632 20874 27660 22170
rect 27724 22098 27752 24239
rect 27816 23594 27844 25230
rect 28172 25220 28224 25226
rect 28172 25162 28224 25168
rect 28184 24818 28212 25162
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 27804 23588 27856 23594
rect 27804 23530 27856 23536
rect 28368 23225 28396 23666
rect 28354 23216 28410 23225
rect 28354 23151 28410 23160
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27620 20868 27672 20874
rect 27620 20810 27672 20816
rect 27710 19408 27766 19417
rect 27710 19343 27766 19352
rect 27620 19236 27672 19242
rect 27620 19178 27672 19184
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26882 14512 26938 14521
rect 26882 14447 26938 14456
rect 26620 14062 26740 14090
rect 26620 12986 26648 14062
rect 26700 14000 26752 14006
rect 26700 13942 26752 13948
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26252 12406 26372 12434
rect 26252 12238 26280 12406
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26252 11218 26280 12174
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 26528 11558 26556 12106
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26528 11370 26556 11494
rect 26436 11354 26556 11370
rect 26424 11348 26556 11354
rect 26476 11342 26556 11348
rect 26424 11290 26476 11296
rect 26620 11218 26648 12922
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26054 11112 26110 11121
rect 26054 11047 26110 11056
rect 26068 9926 26096 11047
rect 26608 10804 26660 10810
rect 26608 10746 26660 10752
rect 26238 10568 26294 10577
rect 26238 10503 26294 10512
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 26068 8090 26096 9862
rect 26252 9586 26280 10503
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26330 10024 26386 10033
rect 26330 9959 26386 9968
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26344 8566 26372 9959
rect 26436 9042 26464 10202
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26332 8560 26384 8566
rect 26332 8502 26384 8508
rect 26528 8430 26556 10406
rect 26620 9518 26648 10746
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26712 8242 26740 13942
rect 26790 12744 26846 12753
rect 26790 12679 26846 12688
rect 26804 8906 26832 12679
rect 26792 8900 26844 8906
rect 26792 8842 26844 8848
rect 26712 8214 26832 8242
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26238 7984 26294 7993
rect 26238 7919 26294 7928
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 26068 5710 26096 7686
rect 26252 6798 26280 7919
rect 26804 7818 26832 8214
rect 26792 7812 26844 7818
rect 26792 7754 26844 7760
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26528 6225 26556 6598
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26514 6216 26570 6225
rect 26240 6180 26292 6186
rect 26514 6151 26570 6160
rect 26240 6122 26292 6128
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26068 5302 26096 5510
rect 26252 5302 26280 6122
rect 26620 5914 26648 6258
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 26240 5296 26292 5302
rect 26240 5238 26292 5244
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 25884 4622 25912 4966
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 25596 4004 25648 4010
rect 25596 3946 25648 3952
rect 25700 3998 25820 4026
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25700 3534 25728 3998
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 25792 3602 25820 3878
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 25884 2650 25912 3062
rect 25976 2650 26004 4082
rect 26252 3738 26280 4762
rect 26804 4690 26832 7754
rect 26896 6905 26924 14447
rect 27080 10033 27108 18838
rect 27632 16522 27660 19178
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27724 15570 27752 19343
rect 27816 18873 27844 22918
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 27908 20602 27936 22578
rect 28262 22536 28318 22545
rect 28262 22471 28264 22480
rect 28316 22471 28318 22480
rect 28264 22442 28316 22448
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 28092 20466 28120 21286
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 27986 20360 28042 20369
rect 27986 20295 28042 20304
rect 28000 18970 28028 20295
rect 28184 20058 28212 21422
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 28276 21185 28304 21286
rect 28262 21176 28318 21185
rect 28262 21111 28318 21120
rect 28264 20868 28316 20874
rect 28264 20810 28316 20816
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28276 19904 28304 20810
rect 28184 19876 28304 19904
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 27802 18864 27858 18873
rect 27802 18799 27858 18808
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27172 13530 27200 14962
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27632 13734 27660 14758
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 27632 12434 27660 13330
rect 27632 12406 27752 12434
rect 27066 10024 27122 10033
rect 27066 9959 27122 9968
rect 27724 9674 27752 12406
rect 27816 10606 27844 15370
rect 27908 13394 27936 17682
rect 28184 17542 28212 19876
rect 28356 19848 28408 19854
rect 28354 19816 28356 19825
rect 28408 19816 28410 19825
rect 28354 19751 28410 19760
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 28000 15026 28028 16934
rect 28080 16516 28132 16522
rect 28080 16458 28132 16464
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27724 9646 27844 9674
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27632 9042 27660 9318
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27816 8537 27844 9646
rect 27908 9450 27936 13126
rect 28092 10826 28120 16458
rect 28184 15586 28212 17478
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28368 17105 28396 17138
rect 28354 17096 28410 17105
rect 28354 17031 28410 17040
rect 28264 15904 28316 15910
rect 28264 15846 28316 15852
rect 28276 15745 28304 15846
rect 28262 15736 28318 15745
rect 28262 15671 28318 15680
rect 28184 15558 28304 15586
rect 28172 12640 28224 12646
rect 28172 12582 28224 12588
rect 28000 10798 28120 10826
rect 28000 9586 28028 10798
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27896 9444 27948 9450
rect 27896 9386 27948 9392
rect 28092 8634 28120 10610
rect 28080 8628 28132 8634
rect 28080 8570 28132 8576
rect 27802 8528 27858 8537
rect 27802 8463 27858 8472
rect 27816 8090 27844 8463
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 26882 6896 26938 6905
rect 26882 6831 26938 6840
rect 27632 6730 27660 7142
rect 27620 6724 27672 6730
rect 27620 6666 27672 6672
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 27264 5914 27292 6258
rect 27816 6254 27844 7754
rect 28184 7410 28212 12582
rect 28276 10962 28304 15558
rect 28354 15056 28410 15065
rect 28354 14991 28410 15000
rect 28368 14414 28396 14991
rect 28460 14618 28488 23054
rect 28552 16114 28580 24550
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 29932 18465 29960 18702
rect 29918 18456 29974 18465
rect 29918 18391 29974 18400
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28368 12345 28396 12786
rect 28354 12336 28410 12345
rect 28354 12271 28410 12280
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 29918 10976 29974 10985
rect 28276 10934 28396 10962
rect 28368 10146 28396 10934
rect 28734 10908 29042 10917
rect 29918 10911 29974 10920
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 29932 10810 29960 10911
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 28276 10118 28396 10146
rect 28276 9178 28304 10118
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 28368 9625 28396 9998
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28354 9616 28410 9625
rect 28354 9551 28410 9560
rect 28448 9580 28500 9586
rect 28448 9522 28500 9528
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28460 8945 28488 9522
rect 28446 8936 28502 8945
rect 28446 8871 28502 8880
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28276 7546 28304 8434
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 29918 7576 29974 7585
rect 28264 7540 28316 7546
rect 29918 7511 29974 7520
rect 28264 7482 28316 7488
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 29932 6798 29960 7511
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 28262 6216 28318 6225
rect 28262 6151 28264 6160
rect 28316 6151 28318 6160
rect 28264 6122 28316 6128
rect 28080 6112 28132 6118
rect 28080 6054 28132 6060
rect 27252 5908 27304 5914
rect 27252 5850 27304 5856
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27172 4826 27200 5646
rect 27896 5568 27948 5574
rect 27896 5510 27948 5516
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27632 4826 27660 5102
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27252 4548 27304 4554
rect 27252 4490 27304 4496
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26436 3058 26464 3946
rect 26976 3528 27028 3534
rect 26974 3496 26976 3505
rect 27028 3496 27030 3505
rect 26974 3431 27030 3440
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 25964 2644 26016 2650
rect 25964 2586 26016 2592
rect 27264 2582 27292 4490
rect 27540 3194 27568 4558
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 27816 3738 27844 4082
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 27908 3534 27936 5510
rect 28092 5234 28120 6054
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28264 5024 28316 5030
rect 28264 4966 28316 4972
rect 28276 4865 28304 4966
rect 28262 4856 28318 4865
rect 28262 4791 28318 4800
rect 28080 4480 28132 4486
rect 28080 4422 28132 4428
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 28092 3058 28120 4422
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 27252 2576 27304 2582
rect 27252 2518 27304 2524
rect 27816 2446 27844 2790
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 22296 1442 22324 2382
rect 21928 1414 22324 1442
rect 21928 800 21956 1414
rect 23216 800 23244 2382
rect 24504 800 24532 2382
rect 25424 1465 25452 2382
rect 25410 1456 25466 1465
rect 25410 1391 25466 1400
rect 25792 800 25820 2382
rect 26436 800 26464 2382
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27724 800 27752 2246
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 6458 200 6514 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 18694 200 18750 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21914 200 21970 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28368 105 28396 2790
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 29104 1306 29132 2926
rect 29932 2145 29960 3334
rect 29918 2136 29974 2145
rect 29918 2071 29974 2080
rect 29012 1278 29132 1306
rect 29012 800 29040 1278
rect 28998 200 29054 800
rect 28354 96 28410 105
rect 28354 31 28410 40
<< via2 >>
rect 2778 29280 2834 29336
rect 1674 27240 1730 27296
rect 1766 25880 1822 25936
rect 1766 24520 1822 24576
rect 1766 23160 1822 23216
rect 3146 27920 3202 27976
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 1766 21800 1822 21856
rect 1766 20440 1822 20496
rect 1766 19796 1768 19816
rect 1768 19796 1820 19816
rect 1820 19796 1822 19816
rect 1766 19760 1822 19796
rect 1766 18400 1822 18456
rect 1766 17060 1822 17096
rect 1766 17040 1768 17060
rect 1768 17040 1820 17060
rect 1820 17040 1822 17060
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 1766 15680 1822 15736
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 1766 14356 1768 14376
rect 1768 14356 1820 14376
rect 1820 14356 1822 14376
rect 1766 14320 1822 14356
rect 1766 13640 1822 13696
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 1766 12280 1822 12336
rect 1766 10920 1822 10976
rect 1766 9560 1822 9616
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 1766 8200 1822 8256
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 1766 6840 1822 6896
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 1766 4800 1822 4856
rect 1766 3440 1822 3496
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 9034 15952 9090 16008
rect 9954 15952 10010 16008
rect 9770 15544 9826 15600
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 10414 14456 10470 14512
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 10874 16360 10930 16416
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 12438 25200 12494 25256
rect 12346 17720 12402 17776
rect 11978 16088 12034 16144
rect 12254 15816 12310 15872
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 10322 8336 10378 8392
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 12530 16904 12586 16960
rect 12714 16904 12770 16960
rect 13450 20848 13506 20904
rect 13174 19352 13230 19408
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 13450 16360 13506 16416
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 3146 2080 3202 2136
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 13726 11736 13782 11792
rect 12806 9424 12862 9480
rect 11978 5616 12034 5672
rect 13450 10512 13506 10568
rect 13542 8880 13598 8936
rect 13634 8472 13690 8528
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 16486 25236 16488 25256
rect 16488 25236 16540 25256
rect 16540 25236 16542 25256
rect 16486 25200 16542 25236
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 15014 21392 15070 21448
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 12990 4664 13046 4720
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14278 10104 14334 10160
rect 14646 14864 14702 14920
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 14554 6704 14610 6760
rect 15566 9424 15622 9480
rect 15382 8744 15438 8800
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 15934 18828 15990 18864
rect 15934 18808 15936 18828
rect 15936 18808 15988 18828
rect 15988 18808 15990 18828
rect 15750 11092 15752 11112
rect 15752 11092 15804 11112
rect 15804 11092 15806 11112
rect 15750 11056 15806 11092
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 16394 15816 16450 15872
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 17406 19216 17462 19272
rect 16486 13776 16542 13832
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18786 22516 18788 22536
rect 18788 22516 18840 22536
rect 18840 22516 18842 22536
rect 18786 22480 18842 22516
rect 18510 21664 18566 21720
rect 18142 20596 18198 20632
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18142 20576 18144 20596
rect 18144 20576 18196 20596
rect 18196 20576 18198 20596
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18142 19796 18144 19816
rect 18144 19796 18196 19816
rect 18196 19796 18198 19816
rect 18142 19760 18198 19796
rect 17406 15000 17462 15056
rect 16670 13232 16726 13288
rect 16578 12300 16634 12336
rect 16578 12280 16580 12300
rect 16580 12280 16632 12300
rect 16632 12280 16634 12300
rect 16946 12588 16948 12608
rect 16948 12588 17000 12608
rect 17000 12588 17002 12608
rect 16946 12552 17002 12588
rect 18694 19796 18696 19816
rect 18696 19796 18748 19816
rect 18748 19796 18750 19816
rect 18694 19760 18750 19796
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18602 17040 18658 17096
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 16762 9052 16764 9072
rect 16764 9052 16816 9072
rect 16816 9052 16818 9072
rect 16762 9016 16818 9052
rect 16394 5652 16396 5672
rect 16396 5652 16448 5672
rect 16448 5652 16450 5672
rect 16394 5616 16450 5652
rect 17222 11076 17278 11112
rect 17222 11056 17224 11076
rect 17224 11056 17276 11076
rect 17276 11056 17278 11076
rect 17038 9560 17094 9616
rect 17222 9596 17224 9616
rect 17224 9596 17276 9616
rect 17276 9596 17278 9616
rect 17222 9560 17278 9596
rect 17222 8472 17278 8528
rect 17406 11212 17462 11248
rect 17406 11192 17408 11212
rect 17408 11192 17460 11212
rect 17460 11192 17462 11212
rect 17406 8508 17408 8528
rect 17408 8508 17460 8528
rect 17460 8508 17462 8528
rect 17406 8472 17462 8508
rect 17406 7284 17408 7304
rect 17408 7284 17460 7304
rect 17460 7284 17462 7304
rect 17406 7248 17462 7284
rect 17866 15544 17922 15600
rect 19522 24248 19578 24304
rect 19614 24148 19616 24168
rect 19616 24148 19668 24168
rect 19668 24148 19670 24168
rect 19614 24112 19670 24148
rect 19706 23296 19762 23352
rect 19246 21428 19248 21448
rect 19248 21428 19300 21448
rect 19300 21428 19302 21448
rect 19246 21392 19302 21428
rect 19062 18264 19118 18320
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18142 13368 18198 13424
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18970 16768 19026 16824
rect 18970 16088 19026 16144
rect 19890 23432 19946 23488
rect 19522 20304 19578 20360
rect 19154 17856 19210 17912
rect 19154 16632 19210 16688
rect 19522 18128 19578 18184
rect 18878 13368 18934 13424
rect 19246 16124 19248 16144
rect 19248 16124 19300 16144
rect 19300 16124 19302 16144
rect 19246 16088 19302 16124
rect 19522 16360 19578 16416
rect 19706 14728 19762 14784
rect 19430 13640 19486 13696
rect 19430 13504 19486 13560
rect 18234 11736 18290 11792
rect 18786 11736 18842 11792
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18694 10104 18750 10160
rect 18234 9424 18290 9480
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 17682 7384 17738 7440
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18786 8880 18842 8936
rect 18786 8780 18788 8800
rect 18788 8780 18840 8800
rect 18840 8780 18842 8800
rect 18786 8744 18842 8780
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18050 4140 18106 4176
rect 18050 4120 18052 4140
rect 18052 4120 18104 4140
rect 18104 4120 18106 4140
rect 18234 4120 18290 4176
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 19614 13776 19670 13832
rect 19706 13504 19762 13560
rect 19890 20440 19946 20496
rect 19890 19352 19946 19408
rect 20166 21664 20222 21720
rect 20258 21392 20314 21448
rect 20166 19216 20222 19272
rect 20258 17176 20314 17232
rect 20350 16496 20406 16552
rect 20442 16396 20444 16416
rect 20444 16396 20496 16416
rect 20496 16396 20498 16416
rect 20442 16360 20498 16396
rect 20258 15988 20260 16008
rect 20260 15988 20312 16008
rect 20312 15988 20314 16008
rect 20258 15952 20314 15988
rect 20074 14592 20130 14648
rect 20166 13912 20222 13968
rect 19706 12552 19762 12608
rect 19798 11092 19800 11112
rect 19800 11092 19852 11112
rect 19852 11092 19854 11112
rect 19798 11056 19854 11092
rect 20074 8880 20130 8936
rect 20810 23432 20866 23488
rect 20994 24112 21050 24168
rect 26238 28600 26294 28656
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 20810 21664 20866 21720
rect 21454 23432 21510 23488
rect 21362 22480 21418 22536
rect 21270 21664 21326 21720
rect 21270 21528 21326 21584
rect 21178 20848 21234 20904
rect 21362 20712 21418 20768
rect 20810 16768 20866 16824
rect 20626 15020 20682 15056
rect 20626 15000 20628 15020
rect 20628 15000 20680 15020
rect 20680 15000 20682 15020
rect 20718 14320 20774 14376
rect 20534 12688 20590 12744
rect 20442 12416 20498 12472
rect 19982 7928 20038 7984
rect 19614 6704 19670 6760
rect 19338 3712 19394 3768
rect 19982 6724 20038 6760
rect 19982 6704 19984 6724
rect 19984 6704 20036 6724
rect 20036 6704 20038 6724
rect 19890 6160 19946 6216
rect 20074 5888 20130 5944
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 20442 10376 20498 10432
rect 20350 8064 20406 8120
rect 20534 10104 20590 10160
rect 20810 13504 20866 13560
rect 20810 13232 20866 13288
rect 22098 25200 22154 25256
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 22650 25336 22706 25392
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 22374 23976 22430 24032
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 21638 21120 21694 21176
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21914 19896 21970 19952
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 22742 22652 22744 22672
rect 22744 22652 22796 22672
rect 22796 22652 22798 22672
rect 22742 22616 22798 22652
rect 22374 19896 22430 19952
rect 22926 22092 22982 22128
rect 22926 22072 22928 22092
rect 22928 22072 22980 22092
rect 22980 22072 22982 22092
rect 23018 21664 23074 21720
rect 23018 21392 23074 21448
rect 22834 19760 22890 19816
rect 23294 23740 23296 23760
rect 23296 23740 23348 23760
rect 23348 23740 23350 23760
rect 23294 23704 23350 23740
rect 23662 22480 23718 22536
rect 23754 21936 23810 21992
rect 23570 21120 23626 21176
rect 22374 17856 22430 17912
rect 22374 17176 22430 17232
rect 22006 17060 22062 17096
rect 22006 17040 22008 17060
rect 22008 17040 22060 17060
rect 22060 17040 22062 17060
rect 22466 16652 22522 16688
rect 22466 16632 22468 16652
rect 22468 16632 22520 16652
rect 22520 16632 22522 16652
rect 22466 16496 22522 16552
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21546 15700 21602 15736
rect 21546 15680 21548 15700
rect 21548 15680 21600 15700
rect 21600 15680 21602 15700
rect 21362 14864 21418 14920
rect 20902 9832 20958 9888
rect 20718 8492 20774 8528
rect 20718 8472 20720 8492
rect 20720 8472 20772 8492
rect 20772 8472 20774 8492
rect 20626 7792 20682 7848
rect 20534 7384 20590 7440
rect 21178 13504 21234 13560
rect 21362 13640 21418 13696
rect 21270 12144 21326 12200
rect 21178 11192 21234 11248
rect 21086 11092 21088 11112
rect 21088 11092 21140 11112
rect 21140 11092 21142 11112
rect 21086 11056 21142 11092
rect 21914 16088 21970 16144
rect 22558 16088 22614 16144
rect 22466 15988 22468 16008
rect 22468 15988 22520 16008
rect 22520 15988 22522 16008
rect 22466 15952 22522 15988
rect 22190 15680 22246 15736
rect 21822 15428 21878 15464
rect 21822 15408 21824 15428
rect 21824 15408 21876 15428
rect 21876 15408 21878 15428
rect 22282 15408 22338 15464
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 22098 13388 22154 13424
rect 22098 13368 22100 13388
rect 22100 13368 22152 13388
rect 22152 13368 22154 13388
rect 22190 13232 22246 13288
rect 22558 14320 22614 14376
rect 22374 13776 22430 13832
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 22282 12860 22284 12880
rect 22284 12860 22336 12880
rect 22336 12860 22338 12880
rect 22282 12824 22338 12860
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 22190 11772 22192 11792
rect 22192 11772 22244 11792
rect 22244 11772 22246 11792
rect 22190 11736 22246 11772
rect 23202 19252 23204 19272
rect 23204 19252 23256 19272
rect 23256 19252 23258 19272
rect 23202 19216 23258 19252
rect 23386 18264 23442 18320
rect 22742 13504 22798 13560
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 22190 10784 22246 10840
rect 21178 9968 21234 10024
rect 22374 10684 22376 10704
rect 22376 10684 22428 10704
rect 22428 10684 22430 10704
rect 22374 10648 22430 10684
rect 22098 10260 22154 10296
rect 22098 10240 22100 10260
rect 22100 10240 22152 10260
rect 22152 10240 22154 10260
rect 22190 10104 22246 10160
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 22558 11736 22614 11792
rect 21362 8492 21418 8528
rect 21362 8472 21364 8492
rect 21364 8472 21416 8492
rect 21416 8472 21418 8492
rect 21638 9036 21694 9072
rect 21638 9016 21640 9036
rect 21640 9016 21692 9036
rect 21692 9016 21694 9036
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 21362 7404 21418 7440
rect 21362 7384 21364 7404
rect 21364 7384 21416 7404
rect 21416 7384 21418 7404
rect 20902 3712 20958 3768
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 22282 7792 22338 7848
rect 22650 9832 22706 9888
rect 22650 9016 22706 9072
rect 22926 12824 22982 12880
rect 22466 8064 22522 8120
rect 22374 6704 22430 6760
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 22558 5228 22614 5264
rect 22558 5208 22560 5228
rect 22560 5208 22612 5228
rect 22612 5208 22614 5228
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 20810 3052 20866 3088
rect 20810 3032 20812 3052
rect 20812 3032 20864 3052
rect 20864 3032 20866 3052
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 23110 15036 23112 15056
rect 23112 15036 23164 15056
rect 23164 15036 23166 15056
rect 23110 15000 23166 15036
rect 23294 14728 23350 14784
rect 23018 11212 23074 11248
rect 23018 11192 23020 11212
rect 23020 11192 23072 11212
rect 23072 11192 23074 11212
rect 23202 13232 23258 13288
rect 23478 14592 23534 14648
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25318 24012 25320 24032
rect 25320 24012 25372 24032
rect 25372 24012 25374 24032
rect 23570 13912 23626 13968
rect 24214 18128 24270 18184
rect 24122 16632 24178 16688
rect 25318 23976 25374 24012
rect 23570 10376 23626 10432
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25318 21528 25374 21584
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 24950 19216 25006 19272
rect 24950 17584 25006 17640
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25134 15816 25190 15872
rect 24398 12180 24400 12200
rect 24400 12180 24452 12200
rect 24452 12180 24454 12200
rect 24398 12144 24454 12180
rect 24214 10784 24270 10840
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 24858 12416 24914 12472
rect 24214 10240 24270 10296
rect 24122 10104 24178 10160
rect 23202 8064 23258 8120
rect 23754 8356 23810 8392
rect 23754 8336 23756 8356
rect 23756 8336 23808 8356
rect 23808 8336 23810 8356
rect 23110 5752 23166 5808
rect 22650 4120 22706 4176
rect 23754 6860 23810 6896
rect 23754 6840 23756 6860
rect 23756 6840 23808 6860
rect 23808 6840 23810 6860
rect 25042 12552 25098 12608
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25870 21664 25926 21720
rect 25686 20440 25742 20496
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 24858 9016 24914 9072
rect 24766 8336 24822 8392
rect 24674 5888 24730 5944
rect 24214 5752 24270 5808
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25318 8880 25374 8936
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 25410 6840 25466 6896
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 25042 3984 25098 4040
rect 25686 11600 25742 11656
rect 26882 25880 26938 25936
rect 25870 9832 25926 9888
rect 26330 13640 26386 13696
rect 26606 14456 26662 14512
rect 27526 24520 27582 24576
rect 29918 27240 29974 27296
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 27710 24248 27766 24304
rect 27158 22616 27214 22672
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28354 23160 28410 23216
rect 27710 19352 27766 19408
rect 26882 14456 26938 14512
rect 26054 11056 26110 11112
rect 26238 10512 26294 10568
rect 26330 9968 26386 10024
rect 26790 12688 26846 12744
rect 26238 7928 26294 7984
rect 26514 6160 26570 6216
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28262 22500 28318 22536
rect 28262 22480 28264 22500
rect 28264 22480 28316 22500
rect 28316 22480 28318 22500
rect 27986 20304 28042 20360
rect 28262 21120 28318 21176
rect 27802 18808 27858 18864
rect 27066 9968 27122 10024
rect 28354 19796 28356 19816
rect 28356 19796 28408 19816
rect 28408 19796 28410 19816
rect 28354 19760 28410 19796
rect 28354 17040 28410 17096
rect 28262 15680 28318 15736
rect 27802 8472 27858 8528
rect 26882 6840 26938 6896
rect 28354 15000 28410 15056
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 29918 18400 29974 18456
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28354 12280 28410 12336
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 29918 10920 29974 10976
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28354 9560 28410 9616
rect 28446 8880 28502 8936
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 29918 7520 29974 7576
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28262 6180 28318 6216
rect 28262 6160 28264 6180
rect 28264 6160 28316 6180
rect 28316 6160 28318 6180
rect 26974 3476 26976 3496
rect 26976 3476 27028 3496
rect 27028 3476 27030 3496
rect 26974 3440 27030 3476
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28262 4800 28318 4856
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 25410 1400 25466 1456
rect 2778 720 2834 776
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
rect 29918 2080 29974 2136
rect 28354 40 28410 96
<< metal3 >>
rect 200 29338 800 29368
rect 2773 29338 2839 29341
rect 200 29336 2839 29338
rect 200 29280 2778 29336
rect 2834 29280 2839 29336
rect 200 29278 2839 29280
rect 200 29248 800 29278
rect 2773 29275 2839 29278
rect 26233 28658 26299 28661
rect 29200 28658 29800 28688
rect 26233 28656 29800 28658
rect 26233 28600 26238 28656
rect 26294 28600 29800 28656
rect 26233 28598 29800 28600
rect 26233 28595 26299 28598
rect 29200 28568 29800 28598
rect 200 27978 800 28008
rect 3141 27978 3207 27981
rect 200 27976 3207 27978
rect 200 27920 3146 27976
rect 3202 27920 3207 27976
rect 200 27918 3207 27920
rect 200 27888 800 27918
rect 3141 27915 3207 27918
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 200 27298 800 27328
rect 1669 27298 1735 27301
rect 200 27296 1735 27298
rect 200 27240 1674 27296
rect 1730 27240 1735 27296
rect 200 27238 1735 27240
rect 200 27208 800 27238
rect 1669 27235 1735 27238
rect 29200 27298 29800 27328
rect 29913 27298 29979 27301
rect 29200 27296 29979 27298
rect 29200 27240 29918 27296
rect 29974 27240 29979 27296
rect 29200 27238 29979 27240
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 29200 27208 29800 27238
rect 29913 27235 29979 27238
rect 28730 27167 29046 27168
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 200 25938 800 25968
rect 1761 25938 1827 25941
rect 200 25936 1827 25938
rect 200 25880 1766 25936
rect 1822 25880 1827 25936
rect 200 25878 1827 25880
rect 200 25848 800 25878
rect 1761 25875 1827 25878
rect 26877 25938 26943 25941
rect 29200 25938 29800 25968
rect 26877 25936 29800 25938
rect 26877 25880 26882 25936
rect 26938 25880 29800 25936
rect 26877 25878 29800 25880
rect 26877 25875 26943 25878
rect 29200 25848 29800 25878
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 17350 25332 17356 25396
rect 17420 25394 17426 25396
rect 22645 25394 22711 25397
rect 17420 25392 22711 25394
rect 17420 25336 22650 25392
rect 22706 25336 22711 25392
rect 17420 25334 22711 25336
rect 17420 25332 17426 25334
rect 22645 25331 22711 25334
rect 12433 25258 12499 25261
rect 16481 25258 16547 25261
rect 12433 25256 16547 25258
rect 12433 25200 12438 25256
rect 12494 25200 16486 25256
rect 16542 25200 16547 25256
rect 12433 25198 16547 25200
rect 12433 25195 12499 25198
rect 16481 25195 16547 25198
rect 22093 25258 22159 25261
rect 23422 25258 23428 25260
rect 22093 25256 23428 25258
rect 22093 25200 22098 25256
rect 22154 25200 23428 25256
rect 22093 25198 23428 25200
rect 22093 25195 22159 25198
rect 23422 25196 23428 25198
rect 23492 25196 23498 25260
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 27521 24578 27587 24581
rect 29200 24578 29800 24608
rect 27521 24576 29800 24578
rect 27521 24520 27526 24576
rect 27582 24520 29800 24576
rect 27521 24518 29800 24520
rect 27521 24515 27587 24518
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 29200 24488 29800 24518
rect 25257 24447 25573 24448
rect 19517 24306 19583 24309
rect 27705 24306 27771 24309
rect 19517 24304 27771 24306
rect 19517 24248 19522 24304
rect 19578 24248 27710 24304
rect 27766 24248 27771 24304
rect 19517 24246 27771 24248
rect 19517 24243 19583 24246
rect 27705 24243 27771 24246
rect 19609 24170 19675 24173
rect 20989 24170 21055 24173
rect 19609 24168 21055 24170
rect 19609 24112 19614 24168
rect 19670 24112 20994 24168
rect 21050 24112 21055 24168
rect 19609 24110 21055 24112
rect 19609 24107 19675 24110
rect 20989 24107 21055 24110
rect 22369 24034 22435 24037
rect 25313 24034 25379 24037
rect 22369 24032 25379 24034
rect 22369 23976 22374 24032
rect 22430 23976 25318 24032
rect 25374 23976 25379 24032
rect 22369 23974 25379 23976
rect 22369 23971 22435 23974
rect 25313 23971 25379 23974
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 23289 23762 23355 23765
rect 23790 23762 23796 23764
rect 23289 23760 23796 23762
rect 23289 23704 23294 23760
rect 23350 23704 23796 23760
rect 23289 23702 23796 23704
rect 23289 23699 23355 23702
rect 23790 23700 23796 23702
rect 23860 23700 23866 23764
rect 19885 23490 19951 23493
rect 19704 23488 19951 23490
rect 19704 23432 19890 23488
rect 19946 23432 19951 23488
rect 19704 23430 19951 23432
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 19704 23357 19764 23430
rect 19885 23427 19951 23430
rect 20805 23492 20871 23493
rect 20805 23488 20852 23492
rect 20916 23490 20922 23492
rect 21449 23490 21515 23493
rect 22502 23490 22508 23492
rect 20805 23432 20810 23488
rect 20805 23428 20852 23432
rect 20916 23430 20962 23490
rect 21449 23488 22508 23490
rect 21449 23432 21454 23488
rect 21510 23432 22508 23488
rect 21449 23430 22508 23432
rect 20916 23428 20922 23430
rect 20805 23427 20871 23428
rect 21449 23427 21515 23430
rect 22502 23428 22508 23430
rect 22572 23428 22578 23492
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 19701 23352 19767 23357
rect 19701 23296 19706 23352
rect 19762 23296 19767 23352
rect 19701 23291 19767 23296
rect 200 23218 800 23248
rect 1761 23218 1827 23221
rect 200 23216 1827 23218
rect 200 23160 1766 23216
rect 1822 23160 1827 23216
rect 200 23158 1827 23160
rect 200 23128 800 23158
rect 1761 23155 1827 23158
rect 28349 23218 28415 23221
rect 29200 23218 29800 23248
rect 28349 23216 29800 23218
rect 28349 23160 28354 23216
rect 28410 23160 29800 23216
rect 28349 23158 29800 23160
rect 28349 23155 28415 23158
rect 29200 23128 29800 23158
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 22737 22674 22803 22677
rect 27153 22674 27219 22677
rect 22737 22672 27219 22674
rect 22737 22616 22742 22672
rect 22798 22616 27158 22672
rect 27214 22616 27219 22672
rect 22737 22614 27219 22616
rect 22737 22611 22803 22614
rect 27153 22611 27219 22614
rect 18781 22538 18847 22541
rect 21357 22538 21423 22541
rect 23657 22540 23723 22541
rect 23606 22538 23612 22540
rect 18781 22536 21423 22538
rect 18781 22480 18786 22536
rect 18842 22480 21362 22536
rect 21418 22480 21423 22536
rect 18781 22478 21423 22480
rect 23566 22478 23612 22538
rect 23676 22536 23723 22540
rect 23718 22480 23723 22536
rect 18781 22475 18847 22478
rect 21357 22475 21423 22478
rect 23606 22476 23612 22478
rect 23676 22476 23723 22480
rect 23657 22475 23723 22476
rect 28257 22538 28323 22541
rect 29200 22538 29800 22568
rect 28257 22536 29800 22538
rect 28257 22480 28262 22536
rect 28318 22480 29800 22536
rect 28257 22478 29800 22480
rect 28257 22475 28323 22478
rect 29200 22448 29800 22478
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 22921 22130 22987 22133
rect 22921 22128 23536 22130
rect 22921 22072 22926 22128
rect 22982 22072 23536 22128
rect 22921 22070 23536 22072
rect 22921 22067 22987 22070
rect 23476 21994 23536 22070
rect 23749 21994 23815 21997
rect 23476 21992 23815 21994
rect 23476 21936 23754 21992
rect 23810 21936 23815 21992
rect 23476 21934 23815 21936
rect 23749 21931 23815 21934
rect 200 21858 800 21888
rect 1761 21858 1827 21861
rect 200 21856 1827 21858
rect 200 21800 1766 21856
rect 1822 21800 1827 21856
rect 200 21798 1827 21800
rect 200 21768 800 21798
rect 1761 21795 1827 21798
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 18505 21722 18571 21725
rect 20161 21722 20227 21725
rect 18505 21720 20227 21722
rect 18505 21664 18510 21720
rect 18566 21664 20166 21720
rect 20222 21664 20227 21720
rect 18505 21662 20227 21664
rect 18505 21659 18571 21662
rect 20161 21659 20227 21662
rect 20805 21722 20871 21725
rect 21265 21722 21331 21725
rect 20805 21720 21331 21722
rect 20805 21664 20810 21720
rect 20866 21664 21270 21720
rect 21326 21664 21331 21720
rect 20805 21662 21331 21664
rect 20805 21659 20871 21662
rect 21265 21659 21331 21662
rect 23013 21722 23079 21725
rect 25865 21722 25931 21725
rect 23013 21720 25931 21722
rect 23013 21664 23018 21720
rect 23074 21664 25870 21720
rect 25926 21664 25931 21720
rect 23013 21662 25931 21664
rect 23013 21659 23079 21662
rect 25865 21659 25931 21662
rect 21265 21586 21331 21589
rect 25313 21586 25379 21589
rect 21265 21584 25379 21586
rect 21265 21528 21270 21584
rect 21326 21528 25318 21584
rect 25374 21528 25379 21584
rect 21265 21526 25379 21528
rect 21265 21523 21331 21526
rect 25313 21523 25379 21526
rect 15009 21450 15075 21453
rect 19241 21450 19307 21453
rect 15009 21448 19307 21450
rect 15009 21392 15014 21448
rect 15070 21392 19246 21448
rect 19302 21392 19307 21448
rect 15009 21390 19307 21392
rect 15009 21387 15075 21390
rect 19241 21387 19307 21390
rect 20253 21450 20319 21453
rect 23013 21450 23079 21453
rect 20253 21448 23079 21450
rect 20253 21392 20258 21448
rect 20314 21392 23018 21448
rect 23074 21392 23079 21448
rect 20253 21390 23079 21392
rect 20253 21387 20319 21390
rect 23013 21387 23079 21390
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 21633 21178 21699 21181
rect 23565 21178 23631 21181
rect 21633 21176 23631 21178
rect 21633 21120 21638 21176
rect 21694 21120 23570 21176
rect 23626 21120 23631 21176
rect 21633 21118 23631 21120
rect 21633 21115 21699 21118
rect 23565 21115 23631 21118
rect 28257 21178 28323 21181
rect 29200 21178 29800 21208
rect 28257 21176 29800 21178
rect 28257 21120 28262 21176
rect 28318 21120 29800 21176
rect 28257 21118 29800 21120
rect 28257 21115 28323 21118
rect 29200 21088 29800 21118
rect 13445 20906 13511 20909
rect 21173 20906 21239 20909
rect 13445 20904 21239 20906
rect 13445 20848 13450 20904
rect 13506 20848 21178 20904
rect 21234 20848 21239 20904
rect 13445 20846 21239 20848
rect 13445 20843 13511 20846
rect 21173 20843 21239 20846
rect 20662 20708 20668 20772
rect 20732 20770 20738 20772
rect 21357 20770 21423 20773
rect 20732 20768 21423 20770
rect 20732 20712 21362 20768
rect 21418 20712 21423 20768
rect 20732 20710 21423 20712
rect 20732 20708 20738 20710
rect 21357 20707 21423 20710
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 18137 20634 18203 20637
rect 18137 20632 19350 20634
rect 18137 20576 18142 20632
rect 18198 20576 19350 20632
rect 18137 20574 19350 20576
rect 18137 20571 18203 20574
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 19290 20498 19350 20574
rect 19885 20498 19951 20501
rect 25681 20498 25747 20501
rect 19290 20496 25747 20498
rect 19290 20440 19890 20496
rect 19946 20440 25686 20496
rect 25742 20440 25747 20496
rect 19290 20438 25747 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 19885 20435 19951 20438
rect 25681 20435 25747 20438
rect 19517 20362 19583 20365
rect 27981 20362 28047 20365
rect 19517 20360 28047 20362
rect 19517 20304 19522 20360
rect 19578 20304 27986 20360
rect 28042 20304 28047 20360
rect 19517 20302 28047 20304
rect 19517 20299 19583 20302
rect 27981 20299 28047 20302
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 21909 19954 21975 19957
rect 22369 19954 22435 19957
rect 21909 19952 22435 19954
rect 21909 19896 21914 19952
rect 21970 19896 22374 19952
rect 22430 19896 22435 19952
rect 21909 19894 22435 19896
rect 21909 19891 21975 19894
rect 22369 19891 22435 19894
rect 200 19818 800 19848
rect 1761 19818 1827 19821
rect 200 19816 1827 19818
rect 200 19760 1766 19816
rect 1822 19760 1827 19816
rect 200 19758 1827 19760
rect 200 19728 800 19758
rect 1761 19755 1827 19758
rect 18137 19818 18203 19821
rect 18689 19818 18755 19821
rect 22829 19818 22895 19821
rect 18137 19816 18755 19818
rect 18137 19760 18142 19816
rect 18198 19760 18694 19816
rect 18750 19760 18755 19816
rect 18137 19758 18755 19760
rect 18137 19755 18203 19758
rect 18689 19755 18755 19758
rect 19934 19816 22895 19818
rect 19934 19760 22834 19816
rect 22890 19760 22895 19816
rect 19934 19758 22895 19760
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 19934 19413 19994 19758
rect 22829 19755 22895 19758
rect 28349 19818 28415 19821
rect 29200 19818 29800 19848
rect 28349 19816 29800 19818
rect 28349 19760 28354 19816
rect 28410 19760 29800 19816
rect 28349 19758 29800 19760
rect 28349 19755 28415 19758
rect 29200 19728 29800 19758
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 13169 19410 13235 19413
rect 19885 19410 19994 19413
rect 13169 19408 19994 19410
rect 13169 19352 13174 19408
rect 13230 19352 19890 19408
rect 19946 19352 19994 19408
rect 13169 19350 19994 19352
rect 13169 19347 13235 19350
rect 19885 19347 19951 19350
rect 23422 19348 23428 19412
rect 23492 19410 23498 19412
rect 27705 19410 27771 19413
rect 23492 19408 27771 19410
rect 23492 19352 27710 19408
rect 27766 19352 27771 19408
rect 23492 19350 27771 19352
rect 23492 19348 23498 19350
rect 27705 19347 27771 19350
rect 17401 19274 17467 19277
rect 20161 19274 20227 19277
rect 17401 19272 20227 19274
rect 17401 19216 17406 19272
rect 17462 19216 20166 19272
rect 20222 19216 20227 19272
rect 17401 19214 20227 19216
rect 17401 19211 17467 19214
rect 20161 19211 20227 19214
rect 23197 19274 23263 19277
rect 24945 19274 25011 19277
rect 23197 19272 25011 19274
rect 23197 19216 23202 19272
rect 23258 19216 24950 19272
rect 25006 19216 25011 19272
rect 23197 19214 25011 19216
rect 23197 19211 23263 19214
rect 24945 19211 25011 19214
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 15929 18866 15995 18869
rect 27797 18866 27863 18869
rect 15929 18864 27863 18866
rect 15929 18808 15934 18864
rect 15990 18808 27802 18864
rect 27858 18808 27863 18864
rect 15929 18806 27863 18808
rect 15929 18803 15995 18806
rect 27797 18803 27863 18806
rect 7892 18528 8208 18529
rect 200 18458 800 18488
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 1761 18458 1827 18461
rect 200 18456 1827 18458
rect 200 18400 1766 18456
rect 1822 18400 1827 18456
rect 200 18398 1827 18400
rect 200 18368 800 18398
rect 1761 18395 1827 18398
rect 29200 18458 29800 18488
rect 29913 18458 29979 18461
rect 29200 18456 29979 18458
rect 29200 18400 29918 18456
rect 29974 18400 29979 18456
rect 29200 18398 29979 18400
rect 29200 18368 29800 18398
rect 29913 18395 29979 18398
rect 19057 18322 19123 18325
rect 23381 18322 23447 18325
rect 19057 18320 23447 18322
rect 19057 18264 19062 18320
rect 19118 18264 23386 18320
rect 23442 18264 23447 18320
rect 19057 18262 23447 18264
rect 19057 18259 19123 18262
rect 23381 18259 23447 18262
rect 19517 18186 19583 18189
rect 24209 18186 24275 18189
rect 19517 18184 24275 18186
rect 19517 18128 19522 18184
rect 19578 18128 24214 18184
rect 24270 18128 24275 18184
rect 19517 18126 24275 18128
rect 19517 18123 19583 18126
rect 24209 18123 24275 18126
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 19149 17914 19215 17917
rect 22369 17914 22435 17917
rect 19149 17912 22435 17914
rect 19149 17856 19154 17912
rect 19210 17856 22374 17912
rect 22430 17856 22435 17912
rect 19149 17854 22435 17856
rect 19149 17851 19215 17854
rect 22369 17851 22435 17854
rect 12341 17778 12407 17781
rect 12341 17776 12450 17778
rect 12341 17720 12346 17776
rect 12402 17720 12450 17776
rect 12341 17715 12450 17720
rect 12390 17642 12450 17715
rect 24945 17642 25011 17645
rect 12390 17640 25011 17642
rect 12390 17584 24950 17640
rect 25006 17584 25011 17640
rect 12390 17582 25011 17584
rect 24945 17579 25011 17582
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 20253 17234 20319 17237
rect 22369 17234 22435 17237
rect 20253 17232 22435 17234
rect 20253 17176 20258 17232
rect 20314 17176 22374 17232
rect 22430 17176 22435 17232
rect 20253 17174 22435 17176
rect 20253 17171 20319 17174
rect 22369 17171 22435 17174
rect 200 17098 800 17128
rect 1761 17098 1827 17101
rect 200 17096 1827 17098
rect 200 17040 1766 17096
rect 1822 17040 1827 17096
rect 200 17038 1827 17040
rect 200 17008 800 17038
rect 1761 17035 1827 17038
rect 18597 17098 18663 17101
rect 22001 17098 22067 17101
rect 18597 17096 22067 17098
rect 18597 17040 18602 17096
rect 18658 17040 22006 17096
rect 22062 17040 22067 17096
rect 18597 17038 22067 17040
rect 18597 17035 18663 17038
rect 22001 17035 22067 17038
rect 28349 17098 28415 17101
rect 29200 17098 29800 17128
rect 28349 17096 29800 17098
rect 28349 17040 28354 17096
rect 28410 17040 29800 17096
rect 28349 17038 29800 17040
rect 28349 17035 28415 17038
rect 29200 17008 29800 17038
rect 12525 16962 12591 16965
rect 12709 16962 12775 16965
rect 12525 16960 12775 16962
rect 12525 16904 12530 16960
rect 12586 16904 12714 16960
rect 12770 16904 12775 16960
rect 12525 16902 12775 16904
rect 12525 16899 12591 16902
rect 12709 16899 12775 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 18965 16826 19031 16829
rect 20805 16826 20871 16829
rect 18965 16824 20871 16826
rect 18965 16768 18970 16824
rect 19026 16768 20810 16824
rect 20866 16768 20871 16824
rect 18965 16766 20871 16768
rect 18965 16763 19031 16766
rect 20805 16763 20871 16766
rect 19149 16690 19215 16693
rect 20662 16690 20668 16692
rect 19149 16688 20668 16690
rect 19149 16632 19154 16688
rect 19210 16632 20668 16688
rect 19149 16630 20668 16632
rect 19149 16627 19215 16630
rect 20662 16628 20668 16630
rect 20732 16628 20738 16692
rect 22461 16690 22527 16693
rect 24117 16690 24183 16693
rect 22461 16688 24183 16690
rect 22461 16632 22466 16688
rect 22522 16632 24122 16688
rect 24178 16632 24183 16688
rect 22461 16630 24183 16632
rect 22461 16627 22527 16630
rect 24117 16627 24183 16630
rect 20345 16554 20411 16557
rect 22461 16554 22527 16557
rect 20345 16552 22527 16554
rect 20345 16496 20350 16552
rect 20406 16496 22466 16552
rect 22522 16496 22527 16552
rect 20345 16494 22527 16496
rect 20345 16491 20411 16494
rect 22461 16491 22527 16494
rect 10869 16418 10935 16421
rect 13445 16418 13511 16421
rect 10869 16416 13511 16418
rect 10869 16360 10874 16416
rect 10930 16360 13450 16416
rect 13506 16360 13511 16416
rect 10869 16358 13511 16360
rect 10869 16355 10935 16358
rect 13445 16355 13511 16358
rect 19517 16418 19583 16421
rect 20437 16418 20503 16421
rect 19517 16416 20503 16418
rect 19517 16360 19522 16416
rect 19578 16360 20442 16416
rect 20498 16360 20503 16416
rect 19517 16358 20503 16360
rect 19517 16355 19583 16358
rect 20437 16355 20503 16358
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 11973 16146 12039 16149
rect 18965 16146 19031 16149
rect 11973 16144 19031 16146
rect 11973 16088 11978 16144
rect 12034 16088 18970 16144
rect 19026 16088 19031 16144
rect 11973 16086 19031 16088
rect 11973 16083 12039 16086
rect 18965 16083 19031 16086
rect 19241 16146 19307 16149
rect 21909 16146 21975 16149
rect 22553 16146 22619 16149
rect 19241 16144 21834 16146
rect 19241 16088 19246 16144
rect 19302 16088 21834 16144
rect 19241 16086 21834 16088
rect 19241 16083 19307 16086
rect 9029 16010 9095 16013
rect 9949 16010 10015 16013
rect 20253 16010 20319 16013
rect 9029 16008 20319 16010
rect 9029 15952 9034 16008
rect 9090 15952 9954 16008
rect 10010 15952 20258 16008
rect 20314 15952 20319 16008
rect 9029 15950 20319 15952
rect 9029 15947 9095 15950
rect 9949 15947 10015 15950
rect 20253 15947 20319 15950
rect 12249 15874 12315 15877
rect 16389 15874 16455 15877
rect 12249 15872 16455 15874
rect 12249 15816 12254 15872
rect 12310 15816 16394 15872
rect 16450 15816 16455 15872
rect 12249 15814 16455 15816
rect 21774 15874 21834 16086
rect 21909 16144 22619 16146
rect 21909 16088 21914 16144
rect 21970 16088 22558 16144
rect 22614 16088 22619 16144
rect 21909 16086 22619 16088
rect 21909 16083 21975 16086
rect 22553 16083 22619 16086
rect 22461 16012 22527 16013
rect 22461 16008 22508 16012
rect 22572 16010 22578 16012
rect 22461 15952 22466 16008
rect 22461 15948 22508 15952
rect 22572 15950 22618 16010
rect 22572 15948 22578 15950
rect 22461 15947 22527 15948
rect 25129 15874 25195 15877
rect 21774 15872 25195 15874
rect 21774 15816 25134 15872
rect 25190 15816 25195 15872
rect 21774 15814 25195 15816
rect 12249 15811 12315 15814
rect 16389 15811 16455 15814
rect 25129 15811 25195 15814
rect 4419 15808 4735 15809
rect 200 15738 800 15768
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 21541 15738 21607 15741
rect 22185 15738 22251 15741
rect 21541 15736 22251 15738
rect 21541 15680 21546 15736
rect 21602 15680 22190 15736
rect 22246 15680 22251 15736
rect 21541 15678 22251 15680
rect 21541 15675 21607 15678
rect 22185 15675 22251 15678
rect 28257 15738 28323 15741
rect 29200 15738 29800 15768
rect 28257 15736 29800 15738
rect 28257 15680 28262 15736
rect 28318 15680 29800 15736
rect 28257 15678 29800 15680
rect 28257 15675 28323 15678
rect 29200 15648 29800 15678
rect 9765 15602 9831 15605
rect 17861 15602 17927 15605
rect 9765 15600 17927 15602
rect 9765 15544 9770 15600
rect 9826 15544 17866 15600
rect 17922 15544 17927 15600
rect 9765 15542 17927 15544
rect 9765 15539 9831 15542
rect 17861 15539 17927 15542
rect 21817 15466 21883 15469
rect 22277 15466 22343 15469
rect 21817 15464 22343 15466
rect 21817 15408 21822 15464
rect 21878 15408 22282 15464
rect 22338 15408 22343 15464
rect 21817 15406 22343 15408
rect 21817 15403 21883 15406
rect 22277 15403 22343 15406
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 17401 15058 17467 15061
rect 20621 15058 20687 15061
rect 17401 15056 20687 15058
rect 17401 15000 17406 15056
rect 17462 15000 20626 15056
rect 20682 15000 20687 15056
rect 17401 14998 20687 15000
rect 17401 14995 17467 14998
rect 20621 14995 20687 14998
rect 20846 14996 20852 15060
rect 20916 15058 20922 15060
rect 23105 15058 23171 15061
rect 20916 15056 23171 15058
rect 20916 15000 23110 15056
rect 23166 15000 23171 15056
rect 20916 14998 23171 15000
rect 20916 14996 20922 14998
rect 23105 14995 23171 14998
rect 28349 15058 28415 15061
rect 29200 15058 29800 15088
rect 28349 15056 29800 15058
rect 28349 15000 28354 15056
rect 28410 15000 29800 15056
rect 28349 14998 29800 15000
rect 28349 14995 28415 14998
rect 29200 14968 29800 14998
rect 14641 14922 14707 14925
rect 21357 14922 21423 14925
rect 14641 14920 21423 14922
rect 14641 14864 14646 14920
rect 14702 14864 21362 14920
rect 21418 14864 21423 14920
rect 14641 14862 21423 14864
rect 14641 14859 14707 14862
rect 21357 14859 21423 14862
rect 19701 14786 19767 14789
rect 23289 14786 23355 14789
rect 19701 14784 23355 14786
rect 19701 14728 19706 14784
rect 19762 14728 23294 14784
rect 23350 14728 23355 14784
rect 19701 14726 23355 14728
rect 19701 14723 19767 14726
rect 23289 14723 23355 14726
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 20069 14650 20135 14653
rect 23473 14650 23539 14653
rect 20069 14648 23539 14650
rect 20069 14592 20074 14648
rect 20130 14592 23478 14648
rect 23534 14592 23539 14648
rect 20069 14590 23539 14592
rect 20069 14587 20135 14590
rect 23473 14587 23539 14590
rect 10409 14514 10475 14517
rect 26601 14514 26667 14517
rect 26877 14514 26943 14517
rect 10409 14512 26943 14514
rect 10409 14456 10414 14512
rect 10470 14456 26606 14512
rect 26662 14456 26882 14512
rect 26938 14456 26943 14512
rect 10409 14454 26943 14456
rect 10409 14451 10475 14454
rect 26601 14451 26667 14454
rect 26877 14451 26943 14454
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 20713 14378 20779 14381
rect 22553 14378 22619 14381
rect 20713 14376 22619 14378
rect 20713 14320 20718 14376
rect 20774 14320 22558 14376
rect 22614 14320 22619 14376
rect 20713 14318 22619 14320
rect 20713 14315 20779 14318
rect 22553 14315 22619 14318
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 20161 13970 20227 13973
rect 23565 13970 23631 13973
rect 20161 13968 23631 13970
rect 20161 13912 20166 13968
rect 20222 13912 23570 13968
rect 23626 13912 23631 13968
rect 20161 13910 23631 13912
rect 20161 13907 20227 13910
rect 23565 13907 23631 13910
rect 16481 13836 16547 13837
rect 16430 13834 16436 13836
rect 16390 13774 16436 13834
rect 16500 13832 16547 13836
rect 16542 13776 16547 13832
rect 16430 13772 16436 13774
rect 16500 13772 16547 13776
rect 16481 13771 16547 13772
rect 19609 13834 19675 13837
rect 22369 13834 22435 13837
rect 19609 13832 22435 13834
rect 19609 13776 19614 13832
rect 19670 13776 22374 13832
rect 22430 13776 22435 13832
rect 19609 13774 22435 13776
rect 19609 13771 19675 13774
rect 22369 13771 22435 13774
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 19425 13698 19491 13701
rect 21357 13698 21423 13701
rect 19425 13696 21423 13698
rect 19425 13640 19430 13696
rect 19486 13640 21362 13696
rect 21418 13640 21423 13696
rect 19425 13638 21423 13640
rect 19425 13635 19491 13638
rect 21357 13635 21423 13638
rect 26325 13698 26391 13701
rect 29200 13698 29800 13728
rect 26325 13696 29800 13698
rect 26325 13640 26330 13696
rect 26386 13640 29800 13696
rect 26325 13638 29800 13640
rect 26325 13635 26391 13638
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 29200 13608 29800 13638
rect 25257 13567 25573 13568
rect 19425 13562 19491 13565
rect 19701 13562 19767 13565
rect 20805 13562 20871 13565
rect 19425 13560 20871 13562
rect 19425 13504 19430 13560
rect 19486 13504 19706 13560
rect 19762 13504 20810 13560
rect 20866 13504 20871 13560
rect 19425 13502 20871 13504
rect 19425 13499 19491 13502
rect 19701 13499 19767 13502
rect 20805 13499 20871 13502
rect 21173 13562 21239 13565
rect 22737 13562 22803 13565
rect 21173 13560 22803 13562
rect 21173 13504 21178 13560
rect 21234 13504 22742 13560
rect 22798 13504 22803 13560
rect 21173 13502 22803 13504
rect 21173 13499 21239 13502
rect 22737 13499 22803 13502
rect 18137 13426 18203 13429
rect 18873 13426 18939 13429
rect 22093 13426 22159 13429
rect 18137 13424 22159 13426
rect 18137 13368 18142 13424
rect 18198 13368 18878 13424
rect 18934 13368 22098 13424
rect 22154 13368 22159 13424
rect 18137 13366 22159 13368
rect 18137 13363 18203 13366
rect 18873 13363 18939 13366
rect 22093 13363 22159 13366
rect 16665 13290 16731 13293
rect 20805 13290 20871 13293
rect 16665 13288 20871 13290
rect 16665 13232 16670 13288
rect 16726 13232 20810 13288
rect 20866 13232 20871 13288
rect 16665 13230 20871 13232
rect 16665 13227 16731 13230
rect 20805 13227 20871 13230
rect 22185 13290 22251 13293
rect 23197 13290 23263 13293
rect 22185 13288 23263 13290
rect 22185 13232 22190 13288
rect 22246 13232 23202 13288
rect 23258 13232 23263 13288
rect 22185 13230 23263 13232
rect 22185 13227 22251 13230
rect 23197 13227 23263 13230
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 22277 12882 22343 12885
rect 22921 12882 22987 12885
rect 22277 12880 22987 12882
rect 22277 12824 22282 12880
rect 22338 12824 22926 12880
rect 22982 12824 22987 12880
rect 22277 12822 22987 12824
rect 22277 12819 22343 12822
rect 22921 12819 22987 12822
rect 20529 12746 20595 12749
rect 26785 12746 26851 12749
rect 20529 12744 26851 12746
rect 20529 12688 20534 12744
rect 20590 12688 26790 12744
rect 26846 12688 26851 12744
rect 20529 12686 26851 12688
rect 20529 12683 20595 12686
rect 26785 12683 26851 12686
rect 16941 12610 17007 12613
rect 17902 12610 17908 12612
rect 16941 12608 17908 12610
rect 16941 12552 16946 12608
rect 17002 12552 17908 12608
rect 16941 12550 17908 12552
rect 16941 12547 17007 12550
rect 17902 12548 17908 12550
rect 17972 12548 17978 12612
rect 19701 12610 19767 12613
rect 25037 12610 25103 12613
rect 19701 12608 25103 12610
rect 19701 12552 19706 12608
rect 19762 12552 25042 12608
rect 25098 12552 25103 12608
rect 19701 12550 25103 12552
rect 19701 12547 19767 12550
rect 25037 12547 25103 12550
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 20437 12474 20503 12477
rect 24853 12474 24919 12477
rect 20437 12472 24919 12474
rect 20437 12416 20442 12472
rect 20498 12416 24858 12472
rect 24914 12416 24919 12472
rect 20437 12414 24919 12416
rect 20437 12411 20503 12414
rect 24853 12411 24919 12414
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 16573 12338 16639 12341
rect 17350 12338 17356 12340
rect 16573 12336 17356 12338
rect 16573 12280 16578 12336
rect 16634 12280 17356 12336
rect 16573 12278 17356 12280
rect 16573 12275 16639 12278
rect 17350 12276 17356 12278
rect 17420 12276 17426 12340
rect 17718 12276 17724 12340
rect 17788 12338 17794 12340
rect 23606 12338 23612 12340
rect 17788 12278 23612 12338
rect 17788 12276 17794 12278
rect 23606 12276 23612 12278
rect 23676 12276 23682 12340
rect 28349 12338 28415 12341
rect 29200 12338 29800 12368
rect 28349 12336 29800 12338
rect 28349 12280 28354 12336
rect 28410 12280 29800 12336
rect 28349 12278 29800 12280
rect 28349 12275 28415 12278
rect 29200 12248 29800 12278
rect 21265 12202 21331 12205
rect 24393 12202 24459 12205
rect 21265 12200 24459 12202
rect 21265 12144 21270 12200
rect 21326 12144 24398 12200
rect 24454 12144 24459 12200
rect 21265 12142 24459 12144
rect 21265 12139 21331 12142
rect 24393 12139 24459 12142
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 13721 11794 13787 11797
rect 18229 11794 18295 11797
rect 18781 11794 18847 11797
rect 13721 11792 18847 11794
rect 13721 11736 13726 11792
rect 13782 11736 18234 11792
rect 18290 11736 18786 11792
rect 18842 11736 18847 11792
rect 13721 11734 18847 11736
rect 13721 11731 13787 11734
rect 18229 11731 18295 11734
rect 18781 11731 18847 11734
rect 22185 11794 22251 11797
rect 22553 11794 22619 11797
rect 22185 11792 22619 11794
rect 22185 11736 22190 11792
rect 22246 11736 22558 11792
rect 22614 11736 22619 11792
rect 22185 11734 22619 11736
rect 22185 11731 22251 11734
rect 22553 11731 22619 11734
rect 16430 11596 16436 11660
rect 16500 11658 16506 11660
rect 25681 11658 25747 11661
rect 16500 11656 25747 11658
rect 16500 11600 25686 11656
rect 25742 11600 25747 11656
rect 16500 11598 25747 11600
rect 16500 11596 16506 11598
rect 25681 11595 25747 11598
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 17401 11250 17467 11253
rect 17718 11250 17724 11252
rect 17401 11248 17724 11250
rect 17401 11192 17406 11248
rect 17462 11192 17724 11248
rect 17401 11190 17724 11192
rect 17401 11187 17467 11190
rect 17718 11188 17724 11190
rect 17788 11188 17794 11252
rect 21173 11250 21239 11253
rect 23013 11250 23079 11253
rect 21173 11248 23079 11250
rect 21173 11192 21178 11248
rect 21234 11192 23018 11248
rect 23074 11192 23079 11248
rect 21173 11190 23079 11192
rect 21173 11187 21239 11190
rect 23013 11187 23079 11190
rect 15745 11114 15811 11117
rect 17217 11114 17283 11117
rect 15745 11112 17283 11114
rect 15745 11056 15750 11112
rect 15806 11056 17222 11112
rect 17278 11056 17283 11112
rect 15745 11054 17283 11056
rect 15745 11051 15811 11054
rect 17217 11051 17283 11054
rect 19793 11114 19859 11117
rect 20846 11114 20852 11116
rect 19793 11112 20852 11114
rect 19793 11056 19798 11112
rect 19854 11056 20852 11112
rect 19793 11054 20852 11056
rect 19793 11051 19859 11054
rect 20846 11052 20852 11054
rect 20916 11052 20922 11116
rect 21081 11114 21147 11117
rect 26049 11114 26115 11117
rect 21081 11112 26115 11114
rect 21081 11056 21086 11112
rect 21142 11056 26054 11112
rect 26110 11056 26115 11112
rect 21081 11054 26115 11056
rect 21081 11051 21147 11054
rect 26049 11051 26115 11054
rect 200 10978 800 11008
rect 1761 10978 1827 10981
rect 200 10976 1827 10978
rect 200 10920 1766 10976
rect 1822 10920 1827 10976
rect 200 10918 1827 10920
rect 200 10888 800 10918
rect 1761 10915 1827 10918
rect 29200 10978 29800 11008
rect 29913 10978 29979 10981
rect 29200 10976 29979 10978
rect 29200 10920 29918 10976
rect 29974 10920 29979 10976
rect 29200 10918 29979 10920
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 29200 10888 29800 10918
rect 29913 10915 29979 10918
rect 28730 10847 29046 10848
rect 22185 10842 22251 10845
rect 24209 10842 24275 10845
rect 22185 10840 24275 10842
rect 22185 10784 22190 10840
rect 22246 10784 24214 10840
rect 24270 10784 24275 10840
rect 22185 10782 24275 10784
rect 22185 10779 22251 10782
rect 24209 10779 24275 10782
rect 18086 10706 18092 10708
rect 13494 10646 18092 10706
rect 13494 10573 13554 10646
rect 18086 10644 18092 10646
rect 18156 10706 18162 10708
rect 22369 10706 22435 10709
rect 18156 10704 22435 10706
rect 18156 10648 22374 10704
rect 22430 10648 22435 10704
rect 18156 10646 22435 10648
rect 18156 10644 18162 10646
rect 22369 10643 22435 10646
rect 13445 10568 13554 10573
rect 13445 10512 13450 10568
rect 13506 10512 13554 10568
rect 13445 10510 13554 10512
rect 13445 10507 13511 10510
rect 17902 10508 17908 10572
rect 17972 10570 17978 10572
rect 26233 10570 26299 10573
rect 17972 10568 26299 10570
rect 17972 10512 26238 10568
rect 26294 10512 26299 10568
rect 17972 10510 26299 10512
rect 17972 10508 17978 10510
rect 26233 10507 26299 10510
rect 20437 10434 20503 10437
rect 23565 10434 23631 10437
rect 20437 10432 23631 10434
rect 20437 10376 20442 10432
rect 20498 10376 23570 10432
rect 23626 10376 23631 10432
rect 20437 10374 23631 10376
rect 20437 10371 20503 10374
rect 23565 10371 23631 10374
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 22093 10298 22159 10301
rect 24209 10298 24275 10301
rect 22093 10296 24275 10298
rect 22093 10240 22098 10296
rect 22154 10240 24214 10296
rect 24270 10240 24275 10296
rect 22093 10238 24275 10240
rect 22093 10235 22159 10238
rect 24209 10235 24275 10238
rect 14273 10162 14339 10165
rect 18689 10162 18755 10165
rect 14273 10160 18755 10162
rect 14273 10104 14278 10160
rect 14334 10104 18694 10160
rect 18750 10104 18755 10160
rect 14273 10102 18755 10104
rect 14273 10099 14339 10102
rect 18689 10099 18755 10102
rect 20529 10162 20595 10165
rect 22185 10162 22251 10165
rect 24117 10162 24183 10165
rect 20529 10160 24183 10162
rect 20529 10104 20534 10160
rect 20590 10104 22190 10160
rect 22246 10104 24122 10160
rect 24178 10104 24183 10160
rect 20529 10102 24183 10104
rect 20529 10099 20595 10102
rect 22185 10099 22251 10102
rect 24117 10099 24183 10102
rect 21173 10026 21239 10029
rect 26325 10026 26391 10029
rect 27061 10026 27127 10029
rect 21173 10024 27127 10026
rect 21173 9968 21178 10024
rect 21234 9968 26330 10024
rect 26386 9968 27066 10024
rect 27122 9968 27127 10024
rect 21173 9966 27127 9968
rect 21173 9963 21239 9966
rect 26325 9963 26391 9966
rect 27061 9963 27127 9966
rect 20662 9828 20668 9892
rect 20732 9890 20738 9892
rect 20897 9890 20963 9893
rect 20732 9888 20963 9890
rect 20732 9832 20902 9888
rect 20958 9832 20963 9888
rect 20732 9830 20963 9832
rect 20732 9828 20738 9830
rect 20897 9827 20963 9830
rect 22645 9890 22711 9893
rect 25865 9890 25931 9893
rect 22645 9888 25931 9890
rect 22645 9832 22650 9888
rect 22706 9832 25870 9888
rect 25926 9832 25931 9888
rect 22645 9830 25931 9832
rect 22645 9827 22711 9830
rect 25865 9827 25931 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 200 9618 800 9648
rect 1761 9618 1827 9621
rect 200 9616 1827 9618
rect 200 9560 1766 9616
rect 1822 9560 1827 9616
rect 200 9558 1827 9560
rect 200 9528 800 9558
rect 1761 9555 1827 9558
rect 17033 9618 17099 9621
rect 17217 9618 17283 9621
rect 17033 9616 17283 9618
rect 17033 9560 17038 9616
rect 17094 9560 17222 9616
rect 17278 9560 17283 9616
rect 17033 9558 17283 9560
rect 17033 9555 17099 9558
rect 17217 9555 17283 9558
rect 28349 9618 28415 9621
rect 29200 9618 29800 9648
rect 28349 9616 29800 9618
rect 28349 9560 28354 9616
rect 28410 9560 29800 9616
rect 28349 9558 29800 9560
rect 28349 9555 28415 9558
rect 29200 9528 29800 9558
rect 12801 9482 12867 9485
rect 15561 9482 15627 9485
rect 18229 9482 18295 9485
rect 12801 9480 18295 9482
rect 12801 9424 12806 9480
rect 12862 9424 15566 9480
rect 15622 9424 18234 9480
rect 18290 9424 18295 9480
rect 12801 9422 18295 9424
rect 12801 9419 12867 9422
rect 15561 9419 15627 9422
rect 18229 9419 18295 9422
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 16757 9074 16823 9077
rect 21633 9074 21699 9077
rect 16757 9072 21699 9074
rect 16757 9016 16762 9072
rect 16818 9016 21638 9072
rect 21694 9016 21699 9072
rect 16757 9014 21699 9016
rect 16757 9011 16823 9014
rect 21633 9011 21699 9014
rect 22645 9074 22711 9077
rect 24853 9074 24919 9077
rect 22645 9072 24919 9074
rect 22645 9016 22650 9072
rect 22706 9016 24858 9072
rect 24914 9016 24919 9072
rect 22645 9014 24919 9016
rect 22645 9011 22711 9014
rect 24853 9011 24919 9014
rect 13537 8938 13603 8941
rect 18781 8938 18847 8941
rect 13537 8936 18847 8938
rect 13537 8880 13542 8936
rect 13598 8880 18786 8936
rect 18842 8880 18847 8936
rect 13537 8878 18847 8880
rect 13537 8875 13603 8878
rect 18781 8875 18847 8878
rect 20069 8938 20135 8941
rect 25313 8938 25379 8941
rect 20069 8936 25379 8938
rect 20069 8880 20074 8936
rect 20130 8880 25318 8936
rect 25374 8880 25379 8936
rect 20069 8878 25379 8880
rect 20069 8875 20135 8878
rect 25313 8875 25379 8878
rect 28441 8938 28507 8941
rect 29200 8938 29800 8968
rect 28441 8936 29800 8938
rect 28441 8880 28446 8936
rect 28502 8880 29800 8936
rect 28441 8878 29800 8880
rect 28441 8875 28507 8878
rect 29200 8848 29800 8878
rect 15377 8802 15443 8805
rect 18781 8802 18847 8805
rect 15377 8800 18847 8802
rect 15377 8744 15382 8800
rect 15438 8744 18786 8800
rect 18842 8744 18847 8800
rect 15377 8742 18847 8744
rect 15377 8739 15443 8742
rect 18781 8739 18847 8742
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 13629 8530 13695 8533
rect 17217 8530 17283 8533
rect 13629 8528 17283 8530
rect 13629 8472 13634 8528
rect 13690 8472 17222 8528
rect 17278 8472 17283 8528
rect 13629 8470 17283 8472
rect 13629 8467 13695 8470
rect 17217 8467 17283 8470
rect 17401 8530 17467 8533
rect 20713 8532 20779 8533
rect 20662 8530 20668 8532
rect 17401 8528 20668 8530
rect 20732 8528 20779 8532
rect 17401 8472 17406 8528
rect 17462 8472 20668 8528
rect 20774 8472 20779 8528
rect 17401 8470 20668 8472
rect 17401 8467 17467 8470
rect 20662 8468 20668 8470
rect 20732 8468 20779 8472
rect 20713 8467 20779 8468
rect 21357 8530 21423 8533
rect 27797 8530 27863 8533
rect 21357 8528 27863 8530
rect 21357 8472 21362 8528
rect 21418 8472 27802 8528
rect 27858 8472 27863 8528
rect 21357 8470 27863 8472
rect 21357 8467 21423 8470
rect 27797 8467 27863 8470
rect 10317 8394 10383 8397
rect 12934 8394 12940 8396
rect 10317 8392 12940 8394
rect 10317 8336 10322 8392
rect 10378 8336 12940 8392
rect 10317 8334 12940 8336
rect 10317 8331 10383 8334
rect 12934 8332 12940 8334
rect 13004 8394 13010 8396
rect 23749 8394 23815 8397
rect 24761 8394 24827 8397
rect 13004 8392 24827 8394
rect 13004 8336 23754 8392
rect 23810 8336 24766 8392
rect 24822 8336 24827 8392
rect 13004 8334 24827 8336
rect 13004 8332 13010 8334
rect 23749 8331 23815 8334
rect 24761 8331 24827 8334
rect 200 8258 800 8288
rect 1761 8258 1827 8261
rect 200 8256 1827 8258
rect 200 8200 1766 8256
rect 1822 8200 1827 8256
rect 200 8198 1827 8200
rect 200 8168 800 8198
rect 1761 8195 1827 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 20345 8122 20411 8125
rect 22461 8122 22527 8125
rect 23197 8122 23263 8125
rect 20345 8120 23263 8122
rect 20345 8064 20350 8120
rect 20406 8064 22466 8120
rect 22522 8064 23202 8120
rect 23258 8064 23263 8120
rect 20345 8062 23263 8064
rect 20345 8059 20411 8062
rect 22461 8059 22527 8062
rect 23197 8059 23263 8062
rect 19977 7986 20043 7989
rect 20662 7986 20668 7988
rect 19977 7984 20668 7986
rect 19977 7928 19982 7984
rect 20038 7928 20668 7984
rect 19977 7926 20668 7928
rect 19977 7923 20043 7926
rect 20662 7924 20668 7926
rect 20732 7924 20738 7988
rect 20846 7924 20852 7988
rect 20916 7986 20922 7988
rect 26233 7986 26299 7989
rect 20916 7984 26299 7986
rect 20916 7928 26238 7984
rect 26294 7928 26299 7984
rect 20916 7926 26299 7928
rect 20916 7924 20922 7926
rect 26233 7923 26299 7926
rect 20621 7850 20687 7853
rect 22277 7850 22343 7853
rect 20621 7848 22343 7850
rect 20621 7792 20626 7848
rect 20682 7792 22282 7848
rect 22338 7792 22343 7848
rect 20621 7790 22343 7792
rect 20621 7787 20687 7790
rect 22277 7787 22343 7790
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 29200 7578 29800 7608
rect 29913 7578 29979 7581
rect 29200 7576 29979 7578
rect 29200 7520 29918 7576
rect 29974 7520 29979 7576
rect 29200 7518 29979 7520
rect 29200 7488 29800 7518
rect 29913 7515 29979 7518
rect 17677 7442 17743 7445
rect 20529 7442 20595 7445
rect 21357 7442 21423 7445
rect 17677 7440 21423 7442
rect 17677 7384 17682 7440
rect 17738 7384 20534 7440
rect 20590 7384 21362 7440
rect 21418 7384 21423 7440
rect 17677 7382 21423 7384
rect 17677 7379 17743 7382
rect 20529 7379 20595 7382
rect 21357 7379 21423 7382
rect 17401 7306 17467 7309
rect 20846 7306 20852 7308
rect 17401 7304 20852 7306
rect 17401 7248 17406 7304
rect 17462 7248 20852 7304
rect 17401 7246 20852 7248
rect 17401 7243 17467 7246
rect 20846 7244 20852 7246
rect 20916 7244 20922 7308
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 200 6898 800 6928
rect 1761 6898 1827 6901
rect 200 6896 1827 6898
rect 200 6840 1766 6896
rect 1822 6840 1827 6896
rect 200 6838 1827 6840
rect 200 6808 800 6838
rect 1761 6835 1827 6838
rect 23749 6900 23815 6901
rect 23749 6896 23796 6900
rect 23860 6898 23866 6900
rect 25405 6898 25471 6901
rect 26877 6898 26943 6901
rect 23749 6840 23754 6896
rect 23749 6836 23796 6840
rect 23860 6838 23906 6898
rect 25405 6896 26943 6898
rect 25405 6840 25410 6896
rect 25466 6840 26882 6896
rect 26938 6840 26943 6896
rect 25405 6838 26943 6840
rect 23860 6836 23866 6838
rect 23749 6835 23815 6836
rect 25405 6835 25471 6838
rect 26877 6835 26943 6838
rect 14549 6762 14615 6765
rect 19609 6762 19675 6765
rect 14549 6760 19675 6762
rect 14549 6704 14554 6760
rect 14610 6704 19614 6760
rect 19670 6704 19675 6760
rect 14549 6702 19675 6704
rect 14549 6699 14615 6702
rect 19609 6699 19675 6702
rect 19977 6762 20043 6765
rect 22369 6762 22435 6765
rect 19977 6760 22435 6762
rect 19977 6704 19982 6760
rect 20038 6704 22374 6760
rect 22430 6704 22435 6760
rect 19977 6702 22435 6704
rect 19977 6699 20043 6702
rect 22369 6699 22435 6702
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 200 6218 800 6248
rect 1761 6218 1827 6221
rect 200 6216 1827 6218
rect 200 6160 1766 6216
rect 1822 6160 1827 6216
rect 200 6158 1827 6160
rect 200 6128 800 6158
rect 1761 6155 1827 6158
rect 19885 6218 19951 6221
rect 26509 6218 26575 6221
rect 19885 6216 26575 6218
rect 19885 6160 19890 6216
rect 19946 6160 26514 6216
rect 26570 6160 26575 6216
rect 19885 6158 26575 6160
rect 19885 6155 19951 6158
rect 26509 6155 26575 6158
rect 28257 6218 28323 6221
rect 29200 6218 29800 6248
rect 28257 6216 29800 6218
rect 28257 6160 28262 6216
rect 28318 6160 29800 6216
rect 28257 6158 29800 6160
rect 28257 6155 28323 6158
rect 29200 6128 29800 6158
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 20069 5946 20135 5949
rect 24669 5946 24735 5949
rect 20069 5944 24735 5946
rect 20069 5888 20074 5944
rect 20130 5888 24674 5944
rect 24730 5888 24735 5944
rect 20069 5886 24735 5888
rect 20069 5883 20135 5886
rect 24669 5883 24735 5886
rect 23105 5810 23171 5813
rect 24209 5810 24275 5813
rect 23105 5808 24275 5810
rect 23105 5752 23110 5808
rect 23166 5752 24214 5808
rect 24270 5752 24275 5808
rect 23105 5750 24275 5752
rect 23105 5747 23171 5750
rect 24209 5747 24275 5750
rect 11973 5674 12039 5677
rect 16389 5674 16455 5677
rect 11973 5672 16455 5674
rect 11973 5616 11978 5672
rect 12034 5616 16394 5672
rect 16450 5616 16455 5672
rect 11973 5614 16455 5616
rect 11973 5611 12039 5614
rect 16389 5611 16455 5614
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 20846 5204 20852 5268
rect 20916 5266 20922 5268
rect 22553 5266 22619 5269
rect 20916 5264 22619 5266
rect 20916 5208 22558 5264
rect 22614 5208 22619 5264
rect 20916 5206 22619 5208
rect 20916 5204 20922 5206
rect 22553 5203 22619 5206
rect 4419 4928 4735 4929
rect 200 4858 800 4888
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 1761 4858 1827 4861
rect 200 4856 1827 4858
rect 200 4800 1766 4856
rect 1822 4800 1827 4856
rect 200 4798 1827 4800
rect 200 4768 800 4798
rect 1761 4795 1827 4798
rect 28257 4858 28323 4861
rect 29200 4858 29800 4888
rect 28257 4856 29800 4858
rect 28257 4800 28262 4856
rect 28318 4800 29800 4856
rect 28257 4798 29800 4800
rect 28257 4795 28323 4798
rect 29200 4768 29800 4798
rect 12985 4724 13051 4725
rect 12934 4660 12940 4724
rect 13004 4722 13051 4724
rect 13004 4720 13096 4722
rect 13046 4664 13096 4720
rect 13004 4662 13096 4664
rect 13004 4660 13051 4662
rect 12985 4659 13051 4660
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 18045 4180 18111 4181
rect 18045 4178 18092 4180
rect 18000 4176 18092 4178
rect 18000 4120 18050 4176
rect 18000 4118 18092 4120
rect 18045 4116 18092 4118
rect 18156 4116 18162 4180
rect 18229 4178 18295 4181
rect 22645 4178 22711 4181
rect 18229 4176 22711 4178
rect 18229 4120 18234 4176
rect 18290 4120 22650 4176
rect 22706 4120 22711 4176
rect 18229 4118 22711 4120
rect 18045 4115 18111 4116
rect 18229 4115 18295 4118
rect 22645 4115 22711 4118
rect 17718 3980 17724 4044
rect 17788 4042 17794 4044
rect 25037 4042 25103 4045
rect 17788 4040 25103 4042
rect 17788 3984 25042 4040
rect 25098 3984 25103 4040
rect 17788 3982 25103 3984
rect 17788 3980 17794 3982
rect 25037 3979 25103 3982
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 19333 3770 19399 3773
rect 20897 3770 20963 3773
rect 19333 3768 20963 3770
rect 19333 3712 19338 3768
rect 19394 3712 20902 3768
rect 20958 3712 20963 3768
rect 19333 3710 20963 3712
rect 19333 3707 19399 3710
rect 20897 3707 20963 3710
rect 200 3498 800 3528
rect 1761 3498 1827 3501
rect 200 3496 1827 3498
rect 200 3440 1766 3496
rect 1822 3440 1827 3496
rect 200 3438 1827 3440
rect 200 3408 800 3438
rect 1761 3435 1827 3438
rect 26969 3498 27035 3501
rect 29200 3498 29800 3528
rect 26969 3496 29800 3498
rect 26969 3440 26974 3496
rect 27030 3440 29800 3496
rect 26969 3438 29800 3440
rect 26969 3435 27035 3438
rect 29200 3408 29800 3438
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 20662 3028 20668 3092
rect 20732 3090 20738 3092
rect 20805 3090 20871 3093
rect 20732 3088 20871 3090
rect 20732 3032 20810 3088
rect 20866 3032 20871 3088
rect 20732 3030 20871 3032
rect 20732 3028 20738 3030
rect 20805 3027 20871 3030
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 7892 2208 8208 2209
rect 200 2138 800 2168
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 3141 2138 3207 2141
rect 200 2136 3207 2138
rect 200 2080 3146 2136
rect 3202 2080 3207 2136
rect 200 2078 3207 2080
rect 200 2048 800 2078
rect 3141 2075 3207 2078
rect 29200 2138 29800 2168
rect 29913 2138 29979 2141
rect 29200 2136 29979 2138
rect 29200 2080 29918 2136
rect 29974 2080 29979 2136
rect 29200 2078 29979 2080
rect 29200 2048 29800 2078
rect 29913 2075 29979 2078
rect 25405 1458 25471 1461
rect 29200 1458 29800 1488
rect 25405 1456 29800 1458
rect 25405 1400 25410 1456
rect 25466 1400 29800 1456
rect 25405 1398 29800 1400
rect 25405 1395 25471 1398
rect 29200 1368 29800 1398
rect 200 778 800 808
rect 2773 778 2839 781
rect 200 776 2839 778
rect 200 720 2778 776
rect 2834 720 2839 776
rect 200 718 2839 720
rect 200 688 800 718
rect 2773 715 2839 718
rect 28349 98 28415 101
rect 29200 98 29800 128
rect 28349 96 29800 98
rect 28349 40 28354 96
rect 28410 40 29800 96
rect 28349 38 29800 40
rect 28349 35 28415 38
rect 29200 8 29800 38
<< via3 >>
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 17356 25332 17420 25396
rect 23428 25196 23492 25260
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 23796 23700 23860 23764
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 20852 23488 20916 23492
rect 20852 23432 20866 23488
rect 20866 23432 20916 23488
rect 20852 23428 20916 23432
rect 22508 23428 22572 23492
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 23612 22536 23676 22540
rect 23612 22480 23662 22536
rect 23662 22480 23676 22536
rect 23612 22476 23676 22480
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 20668 20708 20732 20772
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 23428 19348 23492 19412
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 20668 16628 20732 16692
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 22508 16008 22572 16012
rect 22508 15952 22522 16008
rect 22522 15952 22572 16008
rect 22508 15948 22572 15952
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 20852 14996 20916 15060
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 16436 13832 16500 13836
rect 16436 13776 16486 13832
rect 16486 13776 16500 13832
rect 16436 13772 16500 13776
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 17908 12548 17972 12612
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 17356 12276 17420 12340
rect 17724 12276 17788 12340
rect 23612 12276 23676 12340
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 16436 11596 16500 11660
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 17724 11188 17788 11252
rect 20852 11052 20916 11116
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 18092 10644 18156 10708
rect 17908 10508 17972 10572
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 20668 9828 20732 9892
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 20668 8528 20732 8532
rect 20668 8472 20718 8528
rect 20718 8472 20732 8528
rect 20668 8468 20732 8472
rect 12940 8332 13004 8396
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 20668 7924 20732 7988
rect 20852 7924 20916 7988
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 20852 7244 20916 7308
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 23796 6896 23860 6900
rect 23796 6840 23810 6896
rect 23810 6840 23860 6896
rect 23796 6836 23860 6840
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 20852 5204 20916 5268
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 12940 4720 13004 4724
rect 12940 4664 12990 4720
rect 12990 4664 13004 4720
rect 12940 4660 13004 4664
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 18092 4176 18156 4180
rect 18092 4120 18106 4176
rect 18106 4120 18156 4176
rect 18092 4116 18156 4120
rect 17724 3980 17788 4044
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 20668 3028 20732 3092
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 27776 4737 27792
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 27232 8210 27792
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 27776 11683 27792
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 14836 27232 15156 27792
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 18309 27776 18629 27792
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 17355 25396 17421 25397
rect 17355 25332 17356 25396
rect 17420 25332 17421 25396
rect 17355 25331 17421 25332
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 16435 13836 16501 13837
rect 16435 13772 16436 13836
rect 16500 13772 16501 13836
rect 16435 13771 16501 13772
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 16438 11661 16498 13771
rect 17358 12341 17418 25331
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 21782 27232 22102 27792
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 25255 27776 25575 27792
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 23427 25260 23493 25261
rect 23427 25196 23428 25260
rect 23492 25196 23493 25260
rect 23427 25195 23493 25196
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 20851 23492 20917 23493
rect 20851 23428 20852 23492
rect 20916 23428 20917 23492
rect 20851 23427 20917 23428
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 20667 20772 20733 20773
rect 20667 20708 20668 20772
rect 20732 20708 20733 20772
rect 20667 20707 20733 20708
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 20670 16693 20730 20707
rect 20667 16692 20733 16693
rect 20667 16628 20668 16692
rect 20732 16628 20733 16692
rect 20667 16627 20733 16628
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 20854 15061 20914 23427
rect 21782 22880 22102 23904
rect 22507 23492 22573 23493
rect 22507 23428 22508 23492
rect 22572 23428 22573 23492
rect 22507 23427 22573 23428
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 22510 16013 22570 23427
rect 23430 19413 23490 25195
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 23795 23764 23861 23765
rect 23795 23700 23796 23764
rect 23860 23700 23861 23764
rect 23795 23699 23861 23700
rect 23611 22540 23677 22541
rect 23611 22476 23612 22540
rect 23676 22476 23677 22540
rect 23611 22475 23677 22476
rect 23427 19412 23493 19413
rect 23427 19348 23428 19412
rect 23492 19348 23493 19412
rect 23427 19347 23493 19348
rect 22507 16012 22573 16013
rect 22507 15948 22508 16012
rect 22572 15948 22573 16012
rect 22507 15947 22573 15948
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 20851 15060 20917 15061
rect 20851 14996 20852 15060
rect 20916 14996 20917 15060
rect 20851 14995 20917 14996
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 17907 12612 17973 12613
rect 17907 12548 17908 12612
rect 17972 12548 17973 12612
rect 17907 12547 17973 12548
rect 17355 12340 17421 12341
rect 17355 12276 17356 12340
rect 17420 12276 17421 12340
rect 17355 12275 17421 12276
rect 17723 12340 17789 12341
rect 17723 12276 17724 12340
rect 17788 12276 17789 12340
rect 17723 12275 17789 12276
rect 16435 11660 16501 11661
rect 16435 11596 16436 11660
rect 16500 11596 16501 11660
rect 16435 11595 16501 11596
rect 17726 11253 17786 12275
rect 17723 11252 17789 11253
rect 17723 11188 17724 11252
rect 17788 11188 17789 11252
rect 17723 11187 17789 11188
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 12939 8396 13005 8397
rect 12939 8332 12940 8396
rect 13004 8332 13005 8396
rect 12939 8331 13005 8332
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 12942 4725 13002 8331
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 12939 4724 13005 4725
rect 12939 4660 12940 4724
rect 13004 4660 13005 4724
rect 12939 4659 13005 4660
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 17726 4045 17786 11187
rect 17910 10573 17970 12547
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18091 10708 18157 10709
rect 18091 10644 18092 10708
rect 18156 10644 18157 10708
rect 18091 10643 18157 10644
rect 17907 10572 17973 10573
rect 17907 10508 17908 10572
rect 17972 10508 17973 10572
rect 17907 10507 17973 10508
rect 18094 4181 18154 10643
rect 18309 10368 18629 11392
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 23614 12341 23674 22475
rect 23611 12340 23677 12341
rect 23611 12276 23612 12340
rect 23676 12276 23677 12340
rect 23611 12275 23677 12276
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 20851 11116 20917 11117
rect 20851 11052 20852 11116
rect 20916 11052 20917 11116
rect 20851 11051 20917 11052
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 20667 9892 20733 9893
rect 20667 9828 20668 9892
rect 20732 9828 20733 9892
rect 20667 9827 20733 9828
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 20670 8533 20730 9827
rect 20667 8532 20733 8533
rect 20667 8468 20668 8532
rect 20732 8468 20733 8532
rect 20667 8467 20733 8468
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 20854 7989 20914 11051
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 20667 7988 20733 7989
rect 20667 7924 20668 7988
rect 20732 7924 20733 7988
rect 20667 7923 20733 7924
rect 20851 7988 20917 7989
rect 20851 7924 20852 7988
rect 20916 7924 20917 7988
rect 20851 7923 20917 7924
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18091 4180 18157 4181
rect 18091 4116 18092 4180
rect 18156 4116 18157 4180
rect 18091 4115 18157 4116
rect 17723 4044 17789 4045
rect 17723 3980 17724 4044
rect 17788 3980 17789 4044
rect 17723 3979 17789 3980
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 20670 3093 20730 7923
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 20851 7308 20917 7309
rect 20851 7244 20852 7308
rect 20916 7244 20917 7308
rect 20851 7243 20917 7244
rect 20854 5269 20914 7243
rect 21782 6560 22102 7584
rect 23798 6901 23858 23699
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 23795 6900 23861 6901
rect 23795 6836 23796 6900
rect 23860 6836 23861 6900
rect 23795 6835 23861 6836
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 20851 5268 20917 5269
rect 20851 5204 20852 5268
rect 20916 5204 20917 5268
rect 20851 5203 20917 5204
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 20667 3092 20733 3093
rect 20667 3028 20668 3092
rect 20732 3028 20733 3092
rect 20667 3027 20733 3028
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 27232 29048 27792
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24932 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 25208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 24380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1667941163
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76
timestamp 1667941163
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1667941163
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130
timestamp 1667941163
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1667941163
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1667941163
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1667941163
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1667941163
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1667941163
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1667941163
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1667941163
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_23
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_35
timestamp 1667941163
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1667941163
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1667941163
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1667941163
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_106
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1667941163
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_121
timestamp 1667941163
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1667941163
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_139
timestamp 1667941163
transform 1 0 13892 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_150
timestamp 1667941163
transform 1 0 14904 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1667941163
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1667941163
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1667941163
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1667941163
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1667941163
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1667941163
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1667941163
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1667941163
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_244
timestamp 1667941163
transform 1 0 23552 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_250
timestamp 1667941163
transform 1 0 24104 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1667941163
transform 1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1667941163
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_272
timestamp 1667941163
transform 1 0 26128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1667941163
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1667941163
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1667941163
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1667941163
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1667941163
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_115
timestamp 1667941163
transform 1 0 11684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1667941163
transform 1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_126
timestamp 1667941163
transform 1 0 12696 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1667941163
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1667941163
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1667941163
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_159
timestamp 1667941163
transform 1 0 15732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_174
timestamp 1667941163
transform 1 0 17112 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1667941163
transform 1 0 17848 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1667941163
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_210
timestamp 1667941163
transform 1 0 20424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_220
timestamp 1667941163
transform 1 0 21344 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_234
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_242
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1667941163
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_261
timestamp 1667941163
transform 1 0 25116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_264
timestamp 1667941163
transform 1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_274
timestamp 1667941163
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_278
timestamp 1667941163
transform 1 0 26680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_282
timestamp 1667941163
transform 1 0 27048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1667941163
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_73
timestamp 1667941163
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1667941163
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1667941163
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1667941163
transform 1 0 10212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1667941163
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_123
timestamp 1667941163
transform 1 0 12420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1667941163
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1667941163
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1667941163
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1667941163
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1667941163
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1667941163
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_190
timestamp 1667941163
transform 1 0 18584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_198
timestamp 1667941163
transform 1 0 19320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1667941163
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_209
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_232
timestamp 1667941163
transform 1 0 22448 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_240
timestamp 1667941163
transform 1 0 23184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1667941163
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_258
timestamp 1667941163
transform 1 0 24840 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp 1667941163
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_56
timestamp 1667941163
transform 1 0 6256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_68
timestamp 1667941163
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1667941163
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_90
timestamp 1667941163
transform 1 0 9384 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_98
timestamp 1667941163
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1667941163
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1667941163
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_122
timestamp 1667941163
transform 1 0 12328 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_131
timestamp 1667941163
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1667941163
transform 1 0 14536 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1667941163
transform 1 0 15088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_156
timestamp 1667941163
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_163
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_183
timestamp 1667941163
transform 1 0 17940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1667941163
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1667941163
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1667941163
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_222
timestamp 1667941163
transform 1 0 21528 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1667941163
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1667941163
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_263
timestamp 1667941163
transform 1 0 25300 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_270
timestamp 1667941163
transform 1 0 25944 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1667941163
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_286
timestamp 1667941163
transform 1 0 27416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_290
timestamp 1667941163
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_29
timestamp 1667941163
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_34
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1667941163
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_85
timestamp 1667941163
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_92
timestamp 1667941163
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_99
timestamp 1667941163
transform 1 0 10212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1667941163
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1667941163
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1667941163
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1667941163
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1667941163
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_159
timestamp 1667941163
transform 1 0 15732 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1667941163
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1667941163
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1667941163
transform 1 0 18032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_188
timestamp 1667941163
transform 1 0 18400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1667941163
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_241
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_262
timestamp 1667941163
transform 1 0 25208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_268
timestamp 1667941163
transform 1 0 25760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1667941163
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1667941163
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_47
timestamp 1667941163
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_59
timestamp 1667941163
transform 1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1667941163
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1667941163
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_92
timestamp 1667941163
transform 1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1667941163
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_106
timestamp 1667941163
transform 1 0 10856 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_118
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1667941163
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1667941163
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_159
timestamp 1667941163
transform 1 0 15732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_169
timestamp 1667941163
transform 1 0 16652 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1667941163
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_190
timestamp 1667941163
transform 1 0 18584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_213
timestamp 1667941163
transform 1 0 20700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_225
timestamp 1667941163
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_229
timestamp 1667941163
transform 1 0 22172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_240
timestamp 1667941163
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1667941163
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_272
timestamp 1667941163
transform 1 0 26128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_279
timestamp 1667941163
transform 1 0 26772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_286
timestamp 1667941163
transform 1 0 27416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_293
timestamp 1667941163
transform 1 0 28060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_21
timestamp 1667941163
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_37
timestamp 1667941163
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1667941163
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_65
timestamp 1667941163
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1667941163
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1667941163
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_89
timestamp 1667941163
transform 1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1667941163
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1667941163
transform 1 0 10580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_120
timestamp 1667941163
transform 1 0 12144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1667941163
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1667941163
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_156
timestamp 1667941163
transform 1 0 15456 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_162
timestamp 1667941163
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_175
timestamp 1667941163
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1667941163
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_197
timestamp 1667941163
transform 1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1667941163
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1667941163
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_243
timestamp 1667941163
transform 1 0 23460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_253
timestamp 1667941163
transform 1 0 24380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_271
timestamp 1667941163
transform 1 0 26036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_292
timestamp 1667941163
transform 1 0 27968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1667941163
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1667941163
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_75
timestamp 1667941163
transform 1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1667941163
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_98
timestamp 1667941163
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_102
timestamp 1667941163
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_106
timestamp 1667941163
transform 1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_114
timestamp 1667941163
transform 1 0 11592 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1667941163
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1667941163
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_147
timestamp 1667941163
transform 1 0 14628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1667941163
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1667941163
transform 1 0 15640 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1667941163
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1667941163
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1667941163
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_210
timestamp 1667941163
transform 1 0 20424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_220
timestamp 1667941163
transform 1 0 21344 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_237
timestamp 1667941163
transform 1 0 22908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1667941163
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_278
timestamp 1667941163
transform 1 0 26680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_285
timestamp 1667941163
transform 1 0 27324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_293
timestamp 1667941163
transform 1 0 28060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1667941163
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1667941163
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_87
timestamp 1667941163
transform 1 0 9108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_91
timestamp 1667941163
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1667941163
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1667941163
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_123
timestamp 1667941163
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_151
timestamp 1667941163
transform 1 0 14996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1667941163
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_191
timestamp 1667941163
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_195
timestamp 1667941163
transform 1 0 19044 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1667941163
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_236
timestamp 1667941163
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_243
timestamp 1667941163
transform 1 0 23460 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1667941163
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_290
timestamp 1667941163
transform 1 0 27784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 1667941163
transform 1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1667941163
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1667941163
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp 1667941163
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1667941163
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1667941163
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_75
timestamp 1667941163
transform 1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1667941163
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1667941163
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_111
timestamp 1667941163
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1667941163
transform 1 0 11684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_119
timestamp 1667941163
transform 1 0 12052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_126
timestamp 1667941163
transform 1 0 12696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_134
timestamp 1667941163
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_157
timestamp 1667941163
transform 1 0 15548 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1667941163
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1667941163
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_270
timestamp 1667941163
transform 1 0 25944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1667941163
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_8
timestamp 1667941163
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_20
timestamp 1667941163
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1667941163
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_72
timestamp 1667941163
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1667941163
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1667941163
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1667941163
transform 1 0 10120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_124
timestamp 1667941163
transform 1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_133
timestamp 1667941163
transform 1 0 13340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1667941163
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_153
timestamp 1667941163
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1667941163
transform 1 0 15732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_175
timestamp 1667941163
transform 1 0 17204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1667941163
transform 1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_208
timestamp 1667941163
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1667941163
transform 1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_254
timestamp 1667941163
transform 1 0 24472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_296
timestamp 1667941163
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1667941163
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1667941163
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_49
timestamp 1667941163
transform 1 0 5612 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_71
timestamp 1667941163
transform 1 0 7636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1667941163
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1667941163
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_104
timestamp 1667941163
transform 1 0 10672 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_113
timestamp 1667941163
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_125
timestamp 1667941163
transform 1 0 12604 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_159
timestamp 1667941163
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1667941163
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_215
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1667941163
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_294
timestamp 1667941163
transform 1 0 28152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1667941163
transform 1 0 28520 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_30
timestamp 1667941163
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1667941163
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_63
timestamp 1667941163
transform 1 0 6900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1667941163
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1667941163
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_89
timestamp 1667941163
transform 1 0 9292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1667941163
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1667941163
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1667941163
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1667941163
transform 1 0 12420 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1667941163
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1667941163
transform 1 0 13892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1667941163
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1667941163
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1667941163
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1667941163
transform 1 0 17572 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_203
timestamp 1667941163
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1667941163
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1667941163
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1667941163
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1667941163
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1667941163
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_37
timestamp 1667941163
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_43
timestamp 1667941163
transform 1 0 5060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_55
timestamp 1667941163
transform 1 0 6164 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_67
timestamp 1667941163
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1667941163
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_94
timestamp 1667941163
transform 1 0 9752 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_102
timestamp 1667941163
transform 1 0 10488 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1667941163
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_118
timestamp 1667941163
transform 1 0 11960 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1667941163
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1667941163
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_161
timestamp 1667941163
transform 1 0 15916 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_176
timestamp 1667941163
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_226
timestamp 1667941163
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_282
timestamp 1667941163
transform 1 0 27048 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1667941163
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_64
timestamp 1667941163
transform 1 0 6992 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1667941163
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1667941163
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_94
timestamp 1667941163
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1667941163
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1667941163
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1667941163
transform 1 0 12420 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_130
timestamp 1667941163
transform 1 0 13064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_134
timestamp 1667941163
transform 1 0 13432 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1667941163
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1667941163
transform 1 0 14996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1667941163
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1667941163
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1667941163
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_209
timestamp 1667941163
transform 1 0 20332 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_251
timestamp 1667941163
transform 1 0 24196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_255
timestamp 1667941163
transform 1 0 24564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1667941163
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1667941163
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1667941163
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_61
timestamp 1667941163
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1667941163
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_74
timestamp 1667941163
transform 1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_78
timestamp 1667941163
transform 1 0 8280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_96
timestamp 1667941163
transform 1 0 9936 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_102
timestamp 1667941163
transform 1 0 10488 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1667941163
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1667941163
transform 1 0 12052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_126
timestamp 1667941163
transform 1 0 12696 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 1667941163
transform 1 0 13432 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1667941163
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1667941163
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1667941163
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_217
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_240
timestamp 1667941163
transform 1 0 23184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_262
timestamp 1667941163
transform 1 0 25208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1667941163
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_273
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_47
timestamp 1667941163
transform 1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1667941163
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_63
timestamp 1667941163
transform 1 0 6900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1667941163
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1667941163
transform 1 0 7912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1667941163
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1667941163
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1667941163
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_148
timestamp 1667941163
transform 1 0 14720 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_157
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1667941163
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_208
timestamp 1667941163
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1667941163
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_247
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1667941163
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1667941163
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_63
timestamp 1667941163
transform 1 0 6900 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp 1667941163
transform 1 0 7452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_73
timestamp 1667941163
transform 1 0 7820 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1667941163
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1667941163
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1667941163
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1667941163
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1667941163
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_154
timestamp 1667941163
transform 1 0 15272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1667941163
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_176
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1667941163
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_229
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1667941163
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1667941163
transform 1 0 28520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1667941163
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_20
timestamp 1667941163
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1667941163
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_49
timestamp 1667941163
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_67
timestamp 1667941163
transform 1 0 7268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1667941163
transform 1 0 8280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_91
timestamp 1667941163
transform 1 0 9476 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1667941163
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1667941163
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1667941163
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1667941163
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_141
timestamp 1667941163
transform 1 0 14076 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1667941163
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_178
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_182
timestamp 1667941163
transform 1 0 17848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_198
timestamp 1667941163
transform 1 0 19320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_48
timestamp 1667941163
transform 1 0 5520 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1667941163
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1667941163
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_95
timestamp 1667941163
transform 1 0 9844 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1667941163
transform 1 0 10488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1667941163
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1667941163
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_161
timestamp 1667941163
transform 1 0 15916 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_167
timestamp 1667941163
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_258
timestamp 1667941163
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_266
timestamp 1667941163
transform 1 0 25576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1667941163
transform 1 0 25944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1667941163
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1667941163
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_32
timestamp 1667941163
transform 1 0 4048 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_38
timestamp 1667941163
transform 1 0 4600 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_47
timestamp 1667941163
transform 1 0 5428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_67
timestamp 1667941163
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp 1667941163
transform 1 0 8372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1667941163
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_101
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_124
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1667941163
transform 1 0 13248 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_141
timestamp 1667941163
transform 1 0 14076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1667941163
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1667941163
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1667941163
transform 1 0 18032 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_212
timestamp 1667941163
transform 1 0 20608 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1667941163
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_247
timestamp 1667941163
transform 1 0 23828 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1667941163
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1667941163
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1667941163
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_42
timestamp 1667941163
transform 1 0 4968 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_54
timestamp 1667941163
transform 1 0 6072 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_66
timestamp 1667941163
transform 1 0 7176 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1667941163
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1667941163
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1667941163
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1667941163
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_106
timestamp 1667941163
transform 1 0 10856 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_129
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1667941163
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1667941163
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_185
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1667941163
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_217
timestamp 1667941163
transform 1 0 21068 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_239
timestamp 1667941163
transform 1 0 23092 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1667941163
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_278
timestamp 1667941163
transform 1 0 26680 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_290
timestamp 1667941163
transform 1 0 27784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1667941163
transform 1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1667941163
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_102
timestamp 1667941163
transform 1 0 10488 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1667941163
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1667941163
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_130
timestamp 1667941163
transform 1 0 13064 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1667941163
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_152
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_158
timestamp 1667941163
transform 1 0 15640 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1667941163
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_185
timestamp 1667941163
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_206
timestamp 1667941163
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_213
timestamp 1667941163
transform 1 0 20700 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1667941163
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1667941163
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_64
timestamp 1667941163
transform 1 0 6992 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_72
timestamp 1667941163
transform 1 0 7728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1667941163
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_122
timestamp 1667941163
transform 1 0 12328 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1667941163
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_155
timestamp 1667941163
transform 1 0 15364 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1667941163
transform 1 0 16468 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_179
timestamp 1667941163
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1667941163
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1667941163
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1667941163
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_264
timestamp 1667941163
transform 1 0 25392 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_272
timestamp 1667941163
transform 1 0 26128 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1667941163
transform 1 0 28336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1667941163
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1667941163
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_32
timestamp 1667941163
transform 1 0 4048 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_40
timestamp 1667941163
transform 1 0 4784 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1667941163
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1667941163
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 1667941163
transform 1 0 8648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1667941163
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1667941163
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1667941163
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_131
timestamp 1667941163
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1667941163
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1667941163
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1667941163
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1667941163
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_190
timestamp 1667941163
transform 1 0 18584 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_211
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1667941163
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_50
timestamp 1667941163
transform 1 0 5704 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1667941163
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_63
timestamp 1667941163
transform 1 0 6900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1667941163
transform 1 0 7268 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1667941163
transform 1 0 7636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1667941163
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_101
timestamp 1667941163
transform 1 0 10396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_114
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1667941163
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1667941163
transform 1 0 14536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1667941163
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1667941163
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1667941163
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_273
timestamp 1667941163
transform 1 0 26220 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1667941163
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1667941163
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_45
timestamp 1667941163
transform 1 0 5244 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_63
timestamp 1667941163
transform 1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1667941163
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_89
timestamp 1667941163
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp 1667941163
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_101
timestamp 1667941163
transform 1 0 10396 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1667941163
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_138
timestamp 1667941163
transform 1 0 13800 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1667941163
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_157
timestamp 1667941163
transform 1 0 15548 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_177
timestamp 1667941163
transform 1 0 17388 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_183
timestamp 1667941163
transform 1 0 17940 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_211
timestamp 1667941163
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1667941163
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1667941163
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1667941163
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_54
timestamp 1667941163
transform 1 0 6072 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_66
timestamp 1667941163
transform 1 0 7176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1667941163
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_91
timestamp 1667941163
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_103
timestamp 1667941163
transform 1 0 10580 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1667941163
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_119
timestamp 1667941163
transform 1 0 12052 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1667941163
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1667941163
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_164
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1667941163
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1667941163
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1667941163
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1667941163
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_261
timestamp 1667941163
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_284
timestamp 1667941163
transform 1 0 27232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1667941163
transform 1 0 28336 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_37
timestamp 1667941163
transform 1 0 4508 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1667941163
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_79
timestamp 1667941163
transform 1 0 8372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_85
timestamp 1667941163
transform 1 0 8924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_103
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_129
timestamp 1667941163
transform 1 0 12972 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_135
timestamp 1667941163
transform 1 0 13524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1667941163
transform 1 0 13892 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1667941163
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1667941163
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1667941163
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1667941163
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_267
timestamp 1667941163
transform 1 0 25668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_9
timestamp 1667941163
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1667941163
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_71
timestamp 1667941163
transform 1 0 7636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1667941163
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1667941163
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_122
timestamp 1667941163
transform 1 0 12328 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_130
timestamp 1667941163
transform 1 0 13064 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1667941163
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1667941163
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_169
timestamp 1667941163
transform 1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1667941163
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1667941163
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1667941163
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_278
timestamp 1667941163
transform 1 0 26680 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1667941163
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1667941163
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_62
timestamp 1667941163
transform 1 0 6808 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_71
timestamp 1667941163
transform 1 0 7636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp 1667941163
transform 1 0 8740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1667941163
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_121
timestamp 1667941163
transform 1 0 12236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_133
timestamp 1667941163
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1667941163
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_152
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1667941163
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1667941163
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_212
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_251
timestamp 1667941163
transform 1 0 24196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1667941163
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1667941163
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_47
timestamp 1667941163
transform 1 0 5428 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_57
timestamp 1667941163
transform 1 0 6348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_69
timestamp 1667941163
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1667941163
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_98
timestamp 1667941163
transform 1 0 10120 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_103
timestamp 1667941163
transform 1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1667941163
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1667941163
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1667941163
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_131
timestamp 1667941163
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1667941163
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_162
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1667941163
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_220
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_279
timestamp 1667941163
transform 1 0 26772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_291
timestamp 1667941163
transform 1 0 27876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1667941163
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_35
timestamp 1667941163
transform 1 0 4324 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_86
timestamp 1667941163
transform 1 0 9016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_94
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1667941163
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1667941163
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_130
timestamp 1667941163
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1667941163
transform 1 0 14168 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_154
timestamp 1667941163
transform 1 0 15272 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1667941163
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_174
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_182
timestamp 1667941163
transform 1 0 17848 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_204
timestamp 1667941163
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1667941163
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_238
timestamp 1667941163
transform 1 0 23000 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_263
timestamp 1667941163
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1667941163
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_289
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1667941163
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1667941163
transform 1 0 28520 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_57
timestamp 1667941163
transform 1 0 6348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_69
timestamp 1667941163
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1667941163
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1667941163
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_95
timestamp 1667941163
transform 1 0 9844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_102
timestamp 1667941163
transform 1 0 10488 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_111
timestamp 1667941163
transform 1 0 11316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_117
timestamp 1667941163
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_126
timestamp 1667941163
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_154
timestamp 1667941163
transform 1 0 15272 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1667941163
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1667941163
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_202
timestamp 1667941163
transform 1 0 19688 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_240
timestamp 1667941163
transform 1 0 23184 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1667941163
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_273
timestamp 1667941163
transform 1 0 26220 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1667941163
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_70
timestamp 1667941163
transform 1 0 7544 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_82
timestamp 1667941163
transform 1 0 8648 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_99
timestamp 1667941163
transform 1 0 10212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_131
timestamp 1667941163
transform 1 0 13156 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_141
timestamp 1667941163
transform 1 0 14076 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_148
timestamp 1667941163
transform 1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1667941163
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_174
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_203
timestamp 1667941163
transform 1 0 19780 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1667941163
transform 1 0 20424 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_234
timestamp 1667941163
transform 1 0 22632 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_255
timestamp 1667941163
transform 1 0 24564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_267
timestamp 1667941163
transform 1 0 25668 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_286
timestamp 1667941163
transform 1 0 27416 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_292
timestamp 1667941163
transform 1 0 27968 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1667941163
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_8
timestamp 1667941163
transform 1 0 1840 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1667941163
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_92
timestamp 1667941163
transform 1 0 9568 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_98
timestamp 1667941163
transform 1 0 10120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_102
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_114
timestamp 1667941163
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1667941163
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_162
timestamp 1667941163
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_174
timestamp 1667941163
transform 1 0 17112 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_187
timestamp 1667941163
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_202
timestamp 1667941163
transform 1 0 19688 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_219
timestamp 1667941163
transform 1 0 21252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_232
timestamp 1667941163
transform 1 0 22448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1667941163
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_258
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_293
timestamp 1667941163
transform 1 0 28060 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_80
timestamp 1667941163
transform 1 0 8464 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1667941163
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_94
timestamp 1667941163
transform 1 0 9752 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_103
timestamp 1667941163
transform 1 0 10580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1667941163
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_126
timestamp 1667941163
transform 1 0 12696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_136
timestamp 1667941163
transform 1 0 13616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_152
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_156
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_174
timestamp 1667941163
transform 1 0 17112 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_189
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_199
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_211
timestamp 1667941163
transform 1 0 20516 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_230
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_236
timestamp 1667941163
transform 1 0 22816 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1667941163
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1667941163
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_297
timestamp 1667941163
transform 1 0 28428 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1667941163
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_95
timestamp 1667941163
transform 1 0 9844 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1667941163
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_119
timestamp 1667941163
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1667941163
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_151
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1667941163
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_162
timestamp 1667941163
transform 1 0 16008 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1667941163
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_179
timestamp 1667941163
transform 1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1667941163
transform 1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_215
timestamp 1667941163
transform 1 0 20884 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1667941163
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1667941163
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_258
timestamp 1667941163
transform 1 0 24840 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_266
timestamp 1667941163
transform 1 0 25576 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_270
timestamp 1667941163
transform 1 0 25944 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1667941163
transform 1 0 28244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1667941163
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1667941163
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_32
timestamp 1667941163
transform 1 0 4048 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_44
timestamp 1667941163
transform 1 0 5152 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_78
timestamp 1667941163
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1667941163
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_99
timestamp 1667941163
transform 1 0 10212 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_117
timestamp 1667941163
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_121
timestamp 1667941163
transform 1 0 12236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_128
timestamp 1667941163
transform 1 0 12880 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1667941163
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_155
timestamp 1667941163
transform 1 0 15364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_159
timestamp 1667941163
transform 1 0 15732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_190
timestamp 1667941163
transform 1 0 18584 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_203
timestamp 1667941163
transform 1 0 19780 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_210
timestamp 1667941163
transform 1 0 20424 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_229
timestamp 1667941163
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_233
timestamp 1667941163
transform 1 0 22540 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_239
timestamp 1667941163
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1667941163
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1667941163
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_270
timestamp 1667941163
transform 1 0 25944 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1667941163
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_96
timestamp 1667941163
transform 1 0 9936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_104
timestamp 1667941163
transform 1 0 10672 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_115
timestamp 1667941163
transform 1 0 11684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_119
timestamp 1667941163
transform 1 0 12052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_123
timestamp 1667941163
transform 1 0 12420 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1667941163
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1667941163
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1667941163
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_151
timestamp 1667941163
transform 1 0 14996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1667941163
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_162
timestamp 1667941163
transform 1 0 16008 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1667941163
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1667941163
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1667941163
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_206
timestamp 1667941163
transform 1 0 20056 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1667941163
transform 1 0 20424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1667941163
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_224
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_230
timestamp 1667941163
transform 1 0 22264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_239
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1667941163
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_263
timestamp 1667941163
transform 1 0 25300 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_279
timestamp 1667941163
transform 1 0 26772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1667941163
transform 1 0 27416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_293
timestamp 1667941163
transform 1 0 28060 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1667941163
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1667941163
transform 1 0 8924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_89
timestamp 1667941163
transform 1 0 9292 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_96
timestamp 1667941163
transform 1 0 9936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_103
timestamp 1667941163
transform 1 0 10580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_118
timestamp 1667941163
transform 1 0 11960 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_126
timestamp 1667941163
transform 1 0 12696 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1667941163
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_147
timestamp 1667941163
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_159
timestamp 1667941163
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1667941163
transform 1 0 18400 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1667941163
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1667941163
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_209
timestamp 1667941163
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_235
timestamp 1667941163
transform 1 0 22724 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1667941163
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_252
timestamp 1667941163
transform 1 0 24288 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_260
timestamp 1667941163
transform 1 0 25024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_265
timestamp 1667941163
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1667941163
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_287
timestamp 1667941163
transform 1 0 27508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_291
timestamp 1667941163
transform 1 0 27876 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1667941163
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_103
timestamp 1667941163
transform 1 0 10580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_110
timestamp 1667941163
transform 1 0 11224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_117
timestamp 1667941163
transform 1 0 11868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_124
timestamp 1667941163
transform 1 0 12512 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_131
timestamp 1667941163
transform 1 0 13156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1667941163
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_160
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_166
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1667941163
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_206
timestamp 1667941163
transform 1 0 20056 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_213
timestamp 1667941163
transform 1 0 20700 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_217
timestamp 1667941163
transform 1 0 21068 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_226
timestamp 1667941163
transform 1 0 21896 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_234
timestamp 1667941163
transform 1 0 22632 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_238
timestamp 1667941163
transform 1 0 23000 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1667941163
transform 1 0 24840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_272
timestamp 1667941163
transform 1 0 26128 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_279
timestamp 1667941163
transform 1 0 26772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_287
timestamp 1667941163
transform 1 0 27508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_293
timestamp 1667941163
transform 1 0 28060 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_44
timestamp 1667941163
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_79
timestamp 1667941163
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_91
timestamp 1667941163
transform 1 0 9476 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_99
timestamp 1667941163
transform 1 0 10212 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1667941163
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_124
timestamp 1667941163
transform 1 0 12512 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_130
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_140
timestamp 1667941163
transform 1 0 13984 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_147
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_154
timestamp 1667941163
transform 1 0 15272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_176
timestamp 1667941163
transform 1 0 17296 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_185
timestamp 1667941163
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1667941163
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_204
timestamp 1667941163
transform 1 0 19872 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_212
timestamp 1667941163
transform 1 0 20608 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_230
timestamp 1667941163
transform 1 0 22264 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_242
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_250
timestamp 1667941163
transform 1 0 24104 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_254
timestamp 1667941163
transform 1 0 24472 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1667941163
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_290
timestamp 1667941163
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1667941163
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_36
timestamp 1667941163
transform 1 0 4416 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_40
timestamp 1667941163
transform 1 0 4784 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_44
timestamp 1667941163
transform 1 0 5152 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_56
timestamp 1667941163
transform 1 0 6256 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_68
timestamp 1667941163
transform 1 0 7360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1667941163
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_103
timestamp 1667941163
transform 1 0 10580 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_107
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1667941163
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_125
timestamp 1667941163
transform 1 0 12604 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_129
timestamp 1667941163
transform 1 0 12972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1667941163
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_147
timestamp 1667941163
transform 1 0 14628 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_159
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_175
timestamp 1667941163
transform 1 0 17204 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_183
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_187
timestamp 1667941163
transform 1 0 18308 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_202
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_216
timestamp 1667941163
transform 1 0 20976 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_223
timestamp 1667941163
transform 1 0 21620 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1667941163
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_237
timestamp 1667941163
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1667941163
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_262
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_270
timestamp 1667941163
transform 1 0 25944 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_274
timestamp 1667941163
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_281
timestamp 1667941163
transform 1 0 26956 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1667941163
transform 1 0 27600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_292
timestamp 1667941163
transform 1 0 27968 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1667941163
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_16
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_23
timestamp 1667941163
transform 1 0 3220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_29
timestamp 1667941163
transform 1 0 3772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1667941163
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1667941163
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_118
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_130
timestamp 1667941163
transform 1 0 13064 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_134
timestamp 1667941163
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_141
timestamp 1667941163
transform 1 0 14076 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_148
timestamp 1667941163
transform 1 0 14720 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1667941163
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1667941163
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_184
timestamp 1667941163
transform 1 0 18032 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_191
timestamp 1667941163
transform 1 0 18676 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_198
timestamp 1667941163
transform 1 0 19320 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_214
timestamp 1667941163
transform 1 0 20792 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1667941163
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1667941163
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_242
timestamp 1667941163
transform 1 0 23368 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_256
timestamp 1667941163
transform 1 0 24656 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_262
timestamp 1667941163
transform 1 0 25208 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_266
timestamp 1667941163
transform 1 0 25576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_289
timestamp 1667941163
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1667941163
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_17
timestamp 1667941163
transform 1 0 2668 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_34
timestamp 1667941163
transform 1 0 4232 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_42
timestamp 1667941163
transform 1 0 4968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_48
timestamp 1667941163
transform 1 0 5520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_57
timestamp 1667941163
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_62
timestamp 1667941163
transform 1 0 6808 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_70
timestamp 1667941163
transform 1 0 7544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1667941163
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_90
timestamp 1667941163
transform 1 0 9384 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_98
timestamp 1667941163
transform 1 0 10120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_105
timestamp 1667941163
transform 1 0 10764 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_111
timestamp 1667941163
transform 1 0 11316 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1667941163
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_118
timestamp 1667941163
transform 1 0 11960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_125
timestamp 1667941163
transform 1 0 12604 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1667941163
transform 1 0 14536 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_154
timestamp 1667941163
transform 1 0 15272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_161
timestamp 1667941163
transform 1 0 15916 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_167
timestamp 1667941163
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_169
timestamp 1667941163
transform 1 0 16652 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_175
timestamp 1667941163
transform 1 0 17204 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_183
timestamp 1667941163
transform 1 0 17940 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_217
timestamp 1667941163
transform 1 0 21068 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_223
timestamp 1667941163
transform 1 0 21620 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_225
timestamp 1667941163
transform 1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_230
timestamp 1667941163
transform 1 0 22264 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1667941163
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_272
timestamp 1667941163
transform 1 0 26128 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_281
timestamp 1667941163
transform 1 0 26956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1667941163
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp 1667941163
transform 1 0 28152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_298
timestamp 1667941163
transform 1 0 28520 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0416_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 14168 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 22724 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 11316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 11316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 18216 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 20700 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 15640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 13800 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1667941163
transform 1 0 12788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 19044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 26496 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 17480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 19780 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 20148 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 20792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 12144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 12880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 5244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 7544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 5704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 5704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 23276 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 15916 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 6624 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 10212 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 13432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 12420 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 10948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 10212 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 14720 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 15364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 18400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 26312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 25668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 23552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 23552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 14168 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1667941163
transform 1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1667941163
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0530_
timestamp 1667941163
transform 1 0 12144 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1667941163
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1667941163
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1667941163
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 9568 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1667941163
transform 1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 17756 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 14168 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 8004 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1667941163
transform 1 0 8648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 14720 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 15364 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 11776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1667941163
transform 1 0 9016 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 17940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 14260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 9752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1667941163
transform 1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 18124 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 18584 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 17296 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 13156 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1667941163
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 11776 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 13616 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1667941163
transform 1 0 11960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0607_
timestamp 1667941163
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 15824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 17572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0611_
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 8372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1667941163
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 6532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 6072 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1667941163
transform 1 0 4232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 23460 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 11040 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 9476 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1667941163
transform 1 0 8832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 24932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 24196 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 26312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1667941163
transform 1 0 23092 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 21988 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 20792 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 13064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 9568 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1667941163
transform 1 0 10212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 25024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1667941163
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 25668 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 25944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1667941163
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 12420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1667941163
transform 1 0 12144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 9476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 10120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1667941163
transform 1 0 10304 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1667941163
transform 1 0 11684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 11960 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1667941163
transform 1 0 10304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 21252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 13800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1667941163
transform 1 0 14536 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0692_
timestamp 1667941163
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1667941163
transform 1 0 9292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 14536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1667941163
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1667941163
transform 1 0 12328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1667941163
transform 1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1667941163
transform 1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1667941163
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1667941163
transform 1 0 10580 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0708_
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1667941163
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 6992 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 27784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 20608 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0716_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 20056 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 11592 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 12696 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 27140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 23736 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 27784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 8096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 7268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 27232 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0736_
timestamp 1667941163
transform 1 0 5060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0737_
timestamp 1667941163
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 27784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 27968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 14444 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 27048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 24932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0748_
timestamp 1667941163
transform 1 0 20516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 27140 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0750_
timestamp 1667941163
transform 1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 27784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 6072 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 26496 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 7636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 11592 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 27968 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 16100 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 10304 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 10212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 4876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 17020 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 27508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 4140 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 25576 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 20056 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 14996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 23276 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0795_
timestamp 1667941163
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 4876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 24380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0801_
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0803_
timestamp 1667941163
transform 1 0 11224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12144 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0807_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 20792 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 21988 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0818_
timestamp 1667941163
transform 1 0 15916 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 18216 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 20148 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 20424 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0829_
timestamp 1667941163
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 18492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 17480 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 20056 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0840_
timestamp 1667941163
transform 1 0 16560 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 17664 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 24104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0851_
timestamp 1667941163
transform 1 0 13064 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 21252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 18400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 20148 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 23460 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 20424 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0862_
timestamp 1667941163
transform 1 0 15824 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 21160 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 24932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 25576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 25208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 20884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0873_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 23552 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 25668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 25208 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1667941163
transform 1 0 22816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1667941163
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1667941163
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1667941163
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1667941163
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1667941163
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0890_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24840 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0891_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26312 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 22264 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0893_
timestamp 1667941163
transform 1 0 22080 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 22356 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0895_
timestamp 1667941163
transform 1 0 24564 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0896_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0897_
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0898_
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 26220 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 26220 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 24564 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 24564 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0904_
timestamp 1667941163
transform 1 0 22172 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 18216 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 22724 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform 1 0 23552 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0908_
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 24656 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 26312 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0912_
timestamp 1667941163
transform 1 0 25116 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0913_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0915_
timestamp 1667941163
transform 1 0 26036 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 18216 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0918_
timestamp 1667941163
transform 1 0 26496 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0919_
timestamp 1667941163
transform 1 0 24564 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 25300 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 26312 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0922_
timestamp 1667941163
transform 1 0 24748 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0923_
timestamp 1667941163
transform 1 0 24380 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0924_
timestamp 1667941163
transform 1 0 26220 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0925_
timestamp 1667941163
transform 1 0 26312 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 17112 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0927_
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 22540 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 17940 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0931_
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0932_
timestamp 1667941163
transform 1 0 20976 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0933_
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform 1 0 21620 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 21068 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 18676 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 22540 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0946_
timestamp 1667941163
transform 1 0 21712 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 18124 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 18216 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0951_
timestamp 1667941163
transform 1 0 21160 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 19504 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1667941163
transform 1 0 17940 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1667941163
transform 1 0 22356 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0956_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0957_
timestamp 1667941163
transform 1 0 21712 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform 1 0 18032 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1667941163
transform 1 0 21344 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1667941163
transform 1 0 21620 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1667941163
transform 1 0 19136 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1667941163
transform 1 0 24104 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 13156 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 6440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 25300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 25668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 14352 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 27508 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 3864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 14352 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 27968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 27416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 27324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 25208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19136 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1043_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1043__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1044_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 16192 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1047_
timestamp 1667941163
transform 1 0 22080 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1048_
timestamp 1667941163
transform 1 0 16836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1049__101
timestamp 1667941163
transform 1 0 14260 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 13432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1053_
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 17480 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 9844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1055__102
timestamp 1667941163
transform 1 0 9568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 14536 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1057_
timestamp 1667941163
transform 1 0 20424 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 9292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1059_
timestamp 1667941163
transform 1 0 15088 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 12788 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1061__103
timestamp 1667941163
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 13892 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1067__104
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1068_
timestamp 1667941163
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1069_
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1071_
timestamp 1667941163
transform 1 0 12788 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1072_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1073__105
timestamp 1667941163
transform 1 0 21988 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1074_
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1075_
timestamp 1667941163
transform 1 0 22632 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 23552 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1077_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1078_
timestamp 1667941163
transform 1 0 16468 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1079_
timestamp 1667941163
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1079__106
timestamp 1667941163
transform 1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 9384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1081_
timestamp 1667941163
transform 1 0 17296 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1082_
timestamp 1667941163
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 16008 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1084_
timestamp 1667941163
transform 1 0 12972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1085__107
timestamp 1667941163
transform 1 0 12420 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 9844 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1087_
timestamp 1667941163
transform 1 0 11500 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 20240 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1090_
timestamp 1667941163
transform 1 0 22356 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1091__108
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform 1 0 10856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1093_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1094_
timestamp 1667941163
transform 1 0 26036 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 11960 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 7268 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1097__109
timestamp 1667941163
transform 1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 7636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 8464 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 4600 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 6900 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 13340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1103__110
timestamp 1667941163
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1104_
timestamp 1667941163
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 11224 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 17204 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1107_
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 16560 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1109__111
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 16560 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 21620 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 17756 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 21712 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1114_
timestamp 1667941163
transform 1 0 14720 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1115__112
timestamp 1667941163
transform 1 0 12788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1116_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 14260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1119_
timestamp 1667941163
transform 1 0 11224 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1120_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1121__113
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1123_
timestamp 1667941163
transform 1 0 18952 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform 1 0 18216 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 17664 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1127__114
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 20516 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1130_
timestamp 1667941163
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 20700 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1133__115
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform 1 0 10212 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 15548 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 12420 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1137_
timestamp 1667941163
transform 1 0 9200 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 16560 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 15272 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1139__116
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 16928 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 23184 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1142_
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 23000 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 8280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1145__117
timestamp 1667941163
transform 1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 10396 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform 1 0 6256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1150_
timestamp 1667941163
transform 1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1151__118
timestamp 1667941163
transform 1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 12972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1153_
timestamp 1667941163
transform 1 0 13616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1154_
timestamp 1667941163
transform 1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform 1 0 19596 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 14720 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1157__119
timestamp 1667941163
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1158_
timestamp 1667941163
transform 1 0 10580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 15548 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1161_
timestamp 1667941163
transform 1 0 9936 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1163__120
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1163_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1164_
timestamp 1667941163
transform 1 0 17296 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 13524 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1166_
timestamp 1667941163
transform 1 0 12512 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 14720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1169__121
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1170_
timestamp 1667941163
transform 1 0 22540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 22632 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1172_
timestamp 1667941163
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1174__122
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1174_
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1176_
timestamp 1667941163
transform 1 0 15272 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 16376 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform 1 0 17756 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1178__123
timestamp 1667941163
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1182__124
timestamp 1667941163
transform 1 0 9568 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 12512 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 12420 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1186__125
timestamp 1667941163
transform 1 0 14444 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 11592 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 14444 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1190_
timestamp 1667941163
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1190__126
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 6532 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1192_
timestamp 1667941163
transform 1 0 6624 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 11500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1194__127
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1195_
timestamp 1667941163
transform 1 0 25852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1197_
timestamp 1667941163
transform 1 0 25208 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1198__128
timestamp 1667941163
transform 1 0 4232 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1198_
timestamp 1667941163
transform 1 0 4140 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1200_
timestamp 1667941163
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 7728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1202__129
timestamp 1667941163
transform 1 0 10304 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 21160 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 14996 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 15640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1206_
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1206__130
timestamp 1667941163
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16008 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1208_
timestamp 1667941163
transform 1 0 25576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1209_
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1210__131
timestamp 1667941163
transform 1 0 19596 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 18492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 17848 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 13432 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1214__132
timestamp 1667941163
transform 1 0 14352 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1214_
timestamp 1667941163
transform 1 0 14996 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 20056 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1216_
timestamp 1667941163
transform 1 0 16468 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1667941163
transform 1 0 15088 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1218_
timestamp 1667941163
transform 1 0 8280 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1218__133
timestamp 1667941163
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1219_
timestamp 1667941163
transform 1 0 14260 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 10212 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1221_
timestamp 1667941163
transform 1 0 14352 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1222__134
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1222_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1223_
timestamp 1667941163
transform 1 0 16468 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1224_
timestamp 1667941163
transform 1 0 13156 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1225_
timestamp 1667941163
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1226__135
timestamp 1667941163
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1226_
timestamp 1667941163
transform 1 0 11684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1228_
timestamp 1667941163
transform 1 0 15456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1230__136
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform 1 0 11868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1232_
timestamp 1667941163
transform 1 0 15364 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1234__137
timestamp 1667941163
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1234_
timestamp 1667941163
transform 1 0 20516 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1667941163
transform 1 0 12512 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1236_
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1237_
timestamp 1667941163
transform 1 0 11776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 5244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 3220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 28152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 18400 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 26680 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 11684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 12328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 26036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 28152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 7820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 27140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 3956 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 28152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 25208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 2300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 13432 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 16836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 10396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 28060 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 27324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 5704 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 5170 29200 5226 29800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 3238 29200 3294 29800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 2 nsew signal input
flabel metal3 s 29200 8848 29800 8968 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 3 nsew signal input
flabel metal3 s 29200 18368 29800 18488 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 16762 29200 16818 29800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 5 nsew signal input
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 6 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 8 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 9 nsew signal input
flabel metal3 s 29200 23128 29800 23248 0 FreeSans 480 0 0 0 ccff_head
port 10 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 12 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 13 nsew signal input
flabel metal2 s 25134 29200 25190 29800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 14 nsew signal input
flabel metal3 s 29200 14968 29800 15088 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 15 nsew signal input
flabel metal2 s 9034 29200 9090 29800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 16 nsew signal input
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 17 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 18 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 19 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 20 nsew signal input
flabel metal3 s 29200 25848 29800 25968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 21 nsew signal input
flabel metal3 s 29200 3408 29800 3528 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 22 nsew signal input
flabel metal2 s 19338 29200 19394 29800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 23 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 24 nsew signal input
flabel metal2 s 10966 29200 11022 29800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 25 nsew signal input
flabel metal2 s 12254 29200 12310 29800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 26 nsew signal input
flabel metal2 s 21914 29200 21970 29800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 27 nsew signal input
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 28 nsew signal input
flabel metal3 s 29200 28568 29800 28688 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 29 nsew signal input
flabel metal3 s 29200 24488 29800 24608 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 30 nsew signal input
flabel metal3 s 29200 27208 29800 27328 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 31 nsew signal tristate
flabel metal3 s 29200 6128 29800 6248 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 32 nsew signal tristate
flabel metal2 s 18050 29200 18106 29800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 33 nsew signal tristate
flabel metal2 s 13542 29200 13598 29800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 34 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 35 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 36 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 37 nsew signal tristate
flabel metal3 s 29200 21088 29800 21208 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 38 nsew signal tristate
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 39 nsew signal tristate
flabel metal3 s 29200 10888 29800 11008 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 40 nsew signal tristate
flabel metal2 s 16118 29200 16174 29800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 41 nsew signal tristate
flabel metal2 s 10322 29200 10378 29800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 42 nsew signal tristate
flabel metal3 s 29200 8 29800 128 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 43 nsew signal tristate
flabel metal3 s 29200 22448 29800 22568 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 44 nsew signal tristate
flabel metal2 s 28998 29200 29054 29800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 45 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 46 nsew signal tristate
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 47 nsew signal tristate
flabel metal3 s 29200 4768 29800 4888 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 48 nsew signal tristate
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 49 nsew signal tristate
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal2 s 7746 29200 7802 29800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal2 s 26422 29200 26478 29800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal3 s 29200 12248 29800 12368 0 FreeSans 480 0 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal3 s 29200 7488 29800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal3 s 29200 1368 29800 1488 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal2 s 3882 29200 3938 29800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 29200 9528 29800 9648 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal3 s 29200 19728 29800 19848 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 14830 29200 14886 29800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 662 29200 718 29800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 27710 29200 27766 29800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal2 s 20626 29200 20682 29800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 29642 29200 29698 29800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal3 s 29200 2048 29800 2168 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 29200 15648 29800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 88 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 89 nsew signal input
flabel metal3 s 29200 17008 29800 17128 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 90 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 91 nsew signal input
flabel metal2 s 23846 29200 23902 29800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 23202 29200 23258 29800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 1950 29200 2006 29800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 6458 29200 6514 29800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 96 nsew signal input
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 97 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 pReset
port 98 nsew signal input
flabel metal3 s 29200 13608 29800 13728 0 FreeSans 480 0 0 0 prog_clk
port 99 nsew signal input
flabel metal4 s 4417 2128 4737 27792 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 11363 2128 11683 27792 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 18309 2128 18629 27792 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 25255 2128 25575 27792 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew power bidirectional
flabel metal4 s 7890 2128 8210 27792 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 27792 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 27792 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 27792 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vccd1
rlabel via1 15076 27200 15076 27200 0 vssd1
rlabel metal2 19918 22338 19918 22338 0 _0000_
rlabel metal2 18998 10846 18998 10846 0 _0001_
rlabel metal1 20102 6834 20102 6834 0 _0002_
rlabel metal2 19734 15861 19734 15861 0 _0003_
rlabel metal3 23690 12716 23690 12716 0 _0004_
rlabel metal1 18807 15062 18807 15062 0 _0005_
rlabel metal2 19090 19550 19090 19550 0 _0006_
rlabel metal1 25990 6324 25990 6324 0 _0007_
rlabel metal2 21942 16167 21942 16167 0 _0008_
rlabel metal1 22678 18904 22678 18904 0 _0009_
rlabel metal1 21298 14484 21298 14484 0 _0010_
rlabel via2 21850 15419 21850 15419 0 _0011_
rlabel metal2 23138 17544 23138 17544 0 _0012_
rlabel metal1 20240 8602 20240 8602 0 _0013_
rlabel metal1 19826 13702 19826 13702 0 _0014_
rlabel metal1 19925 8874 19925 8874 0 _0015_
rlabel via2 22310 12869 22310 12869 0 _0016_
rlabel metal1 20654 6188 20654 6188 0 _0017_
rlabel metal1 25208 5882 25208 5882 0 _0018_
rlabel metal2 20286 6188 20286 6188 0 _0019_
rlabel metal1 21206 4794 21206 4794 0 _0020_
rlabel via2 20010 6715 20010 6715 0 _0021_
rlabel metal1 19504 5338 19504 5338 0 _0022_
rlabel metal2 19182 19329 19182 19329 0 _0023_
rlabel metal2 20286 19261 20286 19261 0 _0024_
rlabel metal1 21121 17578 21121 17578 0 _0025_
rlabel metal1 19964 21862 19964 21862 0 _0026_
rlabel metal2 19458 21257 19458 21257 0 _0027_
rlabel metal1 20562 15096 20562 15096 0 _0028_
rlabel metal1 20569 16082 20569 16082 0 _0029_
rlabel metal2 21298 15266 21298 15266 0 _0030_
rlabel metal1 24334 8806 24334 8806 0 _0031_
rlabel metal1 24019 13974 24019 13974 0 _0032_
rlabel metal1 24978 10982 24978 10982 0 _0033_
rlabel metal2 21390 12223 21390 12223 0 _0034_
rlabel metal1 24702 9112 24702 9112 0 _0035_
rlabel metal1 23966 12410 23966 12410 0 _0036_
rlabel metal2 20976 20740 20976 20740 0 _0037_
rlabel metal1 18209 18326 18209 18326 0 _0038_
rlabel metal2 23690 11764 23690 11764 0 _0039_
rlabel metal1 25300 13498 25300 13498 0 _0040_
rlabel metal1 21121 19822 21121 19822 0 _0041_
rlabel metal2 25530 23851 25530 23851 0 _0042_
rlabel metal1 20845 21590 20845 21590 0 _0043_
rlabel metal2 23782 20655 23782 20655 0 _0044_
rlabel metal1 21121 13226 21121 13226 0 _0045_
rlabel metal2 22494 19618 22494 19618 0 _0046_
rlabel metal1 19458 17129 19458 17129 0 _0047_
rlabel metal1 19826 17272 19826 17272 0 _0048_
rlabel metal1 19688 4114 19688 4114 0 _0049_
rlabel metal2 22402 15266 22402 15266 0 _0050_
rlabel metal1 16284 6426 16284 6426 0 _0051_
rlabel metal1 17664 5270 17664 5270 0 _0052_
rlabel metal1 18492 3638 18492 3638 0 _0053_
rlabel metal2 17250 7412 17250 7412 0 _0054_
rlabel metal3 17457 12580 17457 12580 0 _0055_
rlabel metal2 20470 18768 20470 18768 0 _0056_
rlabel metal1 20608 13838 20608 13838 0 _0057_
rlabel metal1 20447 12070 20447 12070 0 _0058_
rlabel via3 20861 23460 20861 23460 0 _0059_
rlabel metal2 22586 16796 22586 16796 0 _0060_
rlabel metal1 25339 19414 25339 19414 0 _0061_
rlabel metal2 23414 20604 23414 20604 0 _0062_
rlabel metal1 24833 10710 24833 10710 0 _0063_
rlabel metal3 25599 19380 25599 19380 0 _0064_
rlabel metal2 19550 24429 19550 24429 0 _0065_
rlabel metal2 20102 9129 20102 9129 0 _0066_
rlabel metal4 20884 9520 20884 9520 0 _0067_
rlabel metal1 16284 18258 16284 18258 0 _0068_
rlabel metal2 20378 16473 20378 16473 0 _0069_
rlabel metal2 19642 10914 19642 10914 0 _0070_
rlabel metal1 21896 23562 21896 23562 0 _0071_
rlabel metal2 19918 18496 19918 18496 0 _0072_
rlabel metal2 19550 18054 19550 18054 0 _0073_
rlabel metal1 21942 25160 21942 25160 0 _0074_
rlabel metal2 20378 4862 20378 4862 0 _0075_
rlabel metal1 11270 6902 11270 6902 0 _0076_
rlabel metal1 19412 3638 19412 3638 0 _0077_
rlabel metal2 10810 6970 10810 6970 0 _0078_
rlabel metal1 14950 16082 14950 16082 0 _0079_
rlabel metal1 19780 3162 19780 3162 0 _0080_
rlabel metal1 14214 3026 14214 3026 0 _0081_
rlabel metal1 21666 24208 21666 24208 0 _0082_
rlabel metal1 11132 26350 11132 26350 0 _0083_
rlabel metal1 11408 16558 11408 16558 0 _0084_
rlabel metal1 7912 6426 7912 6426 0 _0085_
rlabel metal1 19228 25126 19228 25126 0 _0086_
rlabel metal1 14030 26996 14030 26996 0 _0087_
rlabel metal1 12466 25228 12466 25228 0 _0088_
rlabel metal1 18538 4080 18538 4080 0 _0089_
rlabel metal2 19458 26758 19458 26758 0 _0090_
rlabel metal2 17802 11322 17802 11322 0 _0091_
rlabel metal1 25990 3026 25990 3026 0 _0092_
rlabel metal1 20608 24378 20608 24378 0 _0093_
rlabel metal2 13110 24820 13110 24820 0 _0094_
rlabel metal2 5842 14212 5842 14212 0 _0095_
rlabel metal1 5842 11866 5842 11866 0 _0096_
rlabel metal2 26082 6698 26082 6698 0 _0097_
rlabel metal1 15548 16422 15548 16422 0 _0098_
rlabel metal2 9614 11900 9614 11900 0 _0099_
rlabel metal2 7222 11322 7222 11322 0 _0100_
rlabel metal2 11178 17340 11178 17340 0 _0101_
rlabel metal2 12650 8602 12650 8602 0 _0102_
rlabel metal1 10488 21998 10488 21998 0 _0103_
rlabel metal1 9982 14858 9982 14858 0 _0104_
rlabel metal2 15686 18972 15686 18972 0 _0105_
rlabel metal1 15594 6732 15594 6732 0 _0106_
rlabel metal1 26082 23086 26082 23086 0 _0107_
rlabel metal2 10994 19958 10994 19958 0 _0108_
rlabel metal2 22402 3910 22402 3910 0 _0109_
rlabel metal2 14306 4998 14306 4998 0 _0110_
rlabel metal1 13616 3706 13616 3706 0 _0111_
rlabel metal1 16514 5338 16514 5338 0 _0112_
rlabel metal2 12834 11424 12834 11424 0 _0113_
rlabel metal1 11684 9690 11684 9690 0 _0114_
rlabel metal1 8510 6970 8510 6970 0 _0115_
rlabel metal1 10396 6154 10396 6154 0 _0116_
rlabel metal2 12374 5508 12374 5508 0 _0117_
rlabel metal1 9614 5338 9614 5338 0 _0118_
rlabel metal2 12098 4250 12098 4250 0 _0119_
rlabel metal1 9062 4080 9062 4080 0 _0120_
rlabel metal1 11178 14416 11178 14416 0 _0121_
rlabel metal2 9246 9724 9246 9724 0 _0122_
rlabel metal1 7038 10778 7038 10778 0 _0123_
rlabel metal1 14306 19346 14306 19346 0 _0124_
rlabel metal1 17434 21114 17434 21114 0 _0125_
rlabel metal1 13570 14382 13570 14382 0 _0126_
rlabel metal1 8878 23732 8878 23732 0 _0127_
rlabel metal1 15594 24140 15594 24140 0 _0128_
rlabel metal1 9430 24650 9430 24650 0 _0129_
rlabel metal2 15686 16014 15686 16014 0 _0130_
rlabel metal2 17158 8908 17158 8908 0 _0131_
rlabel metal1 10488 12410 10488 12410 0 _0132_
rlabel metal1 19596 21998 19596 21998 0 _0133_
rlabel metal1 18722 24786 18722 24786 0 _0134_
rlabel metal2 17526 23290 17526 23290 0 _0135_
rlabel metal2 13754 8942 13754 8942 0 _0136_
rlabel metal2 12006 17850 12006 17850 0 _0137_
rlabel metal2 12006 19652 12006 19652 0 _0138_
rlabel metal1 19136 11254 19136 11254 0 _0139_
rlabel metal1 15870 20434 15870 20434 0 _0140_
rlabel metal1 15916 12410 15916 12410 0 _0141_
rlabel metal2 8418 18054 8418 18054 0 _0142_
rlabel metal1 13340 4794 13340 4794 0 _0143_
rlabel metal2 12006 3706 12006 3706 0 _0144_
rlabel metal1 7590 19380 7590 19380 0 _0145_
rlabel metal1 7498 16762 7498 16762 0 _0146_
rlabel metal1 5290 18224 5290 18224 0 _0147_
rlabel metal1 9292 22610 9292 22610 0 _0148_
rlabel metal1 24702 25874 24702 25874 0 _0149_
rlabel metal1 22494 26350 22494 26350 0 _0150_
rlabel metal2 9890 18700 9890 18700 0 _0151_
rlabel metal2 11086 15470 11086 15470 0 _0152_
rlabel metal1 10534 21488 10534 21488 0 _0153_
rlabel metal1 9016 4590 9016 4590 0 _0154_
rlabel metal1 13340 8330 13340 8330 0 _0155_
rlabel metal1 9936 13906 9936 13906 0 _0156_
rlabel metal1 17710 10610 17710 10610 0 _0157_
rlabel metal1 25530 23698 25530 23698 0 _0158_
rlabel metal1 23092 26350 23092 26350 0 _0159_
rlabel metal1 12328 10642 12328 10642 0 _0160_
rlabel metal1 9936 13838 9936 13838 0 _0161_
rlabel metal2 10534 19516 10534 19516 0 _0162_
rlabel metal2 11914 17646 11914 17646 0 _0163_
rlabel metal1 12190 23664 12190 23664 0 _0164_
rlabel metal1 10764 24650 10764 24650 0 _0165_
rlabel metal1 14904 22610 14904 22610 0 _0166_
rlabel metal1 14628 21862 14628 21862 0 _0167_
rlabel metal1 9154 21998 9154 21998 0 _0168_
rlabel metal1 13478 12886 13478 12886 0 _0169_
rlabel metal2 12374 17476 12374 17476 0 _0170_
rlabel metal1 13754 16048 13754 16048 0 _0171_
rlabel metal1 10902 9690 10902 9690 0 _0172_
rlabel metal1 18630 2414 18630 2414 0 _0173_
rlabel metal1 15916 15470 15916 15470 0 _0174_
rlabel metal1 20930 19346 20930 19346 0 _0175_
rlabel metal1 17388 21522 17388 21522 0 _0176_
rlabel metal1 17204 20434 17204 20434 0 _0177_
rlabel metal1 18952 14382 18952 14382 0 _0178_
rlabel metal2 18722 21454 18722 21454 0 _0179_
rlabel metal1 17342 18734 17342 18734 0 _0180_
rlabel metal1 17572 19346 17572 19346 0 _0181_
rlabel metal1 18860 3978 18860 3978 0 _0182_
rlabel metal1 18492 2618 18492 2618 0 _0183_
rlabel metal1 13846 10166 13846 10166 0 _0184_
rlabel metal2 16422 8296 16422 8296 0 _0185_
rlabel metal2 14306 14076 14306 14076 0 _0186_
rlabel metal1 23690 3706 23690 3706 0 _0187_
rlabel metal1 15318 15538 15318 15538 0 _0188_
rlabel metal1 15042 17612 15042 17612 0 _0189_
rlabel metal1 14306 12682 14306 12682 0 _0190_
rlabel metal1 14950 13498 14950 13498 0 _0191_
rlabel metal2 13570 20944 13570 20944 0 _0192_
rlabel metal1 15226 12954 15226 12954 0 _0193_
rlabel metal1 16284 21114 16284 21114 0 _0194_
rlabel metal1 9706 21862 9706 21862 0 _0195_
rlabel metal1 14812 22406 14812 22406 0 _0196_
rlabel metal1 20746 21930 20746 21930 0 _0197_
rlabel metal1 9384 18802 9384 18802 0 _0198_
rlabel metal1 15272 21454 15272 21454 0 _0199_
rlabel metal1 13754 23664 13754 23664 0 _0200_
rlabel metal2 11822 24956 11822 24956 0 _0201_
rlabel metal1 12374 17034 12374 17034 0 _0202_
rlabel metal1 15272 23630 15272 23630 0 _0203_
rlabel metal2 14122 24956 14122 24956 0 _0204_
rlabel metal1 13800 22066 13800 22066 0 _0205_
rlabel metal1 11914 14008 11914 14008 0 _0206_
rlabel metal2 11086 18802 11086 18802 0 _0207_
rlabel metal2 12926 11356 12926 11356 0 _0208_
rlabel metal2 14122 12070 14122 12070 0 _0209_
rlabel metal1 11638 20026 11638 20026 0 _0210_
rlabel metal1 12788 11322 12788 11322 0 _0211_
rlabel metal2 25714 24004 25714 24004 0 _0212_
rlabel metal2 22678 26724 22678 26724 0 _0213_
rlabel metal2 17526 11458 17526 11458 0 _0214_
rlabel metal1 24656 23834 24656 23834 0 _0215_
rlabel metal1 24932 24718 24932 24718 0 _0216_
rlabel metal1 15594 11866 15594 11866 0 _0217_
rlabel metal1 14858 9690 14858 9690 0 _0218_
rlabel metal1 9154 12886 9154 12886 0 _0219_
rlabel metal1 9384 4794 9384 4794 0 _0220_
rlabel metal2 14398 6120 14398 6120 0 _0221_
rlabel metal1 9062 14586 9062 14586 0 _0222_
rlabel metal2 16514 6222 16514 6222 0 _0223_
rlabel metal2 10902 15759 10902 15759 0 _0224_
rlabel metal2 10350 21148 10350 21148 0 _0225_
rlabel metal1 9890 17714 9890 17714 0 _0226_
rlabel metal1 11224 15402 11224 15402 0 _0227_
rlabel metal1 20700 24038 20700 24038 0 _0228_
rlabel metal2 10626 15810 10626 15810 0 _0229_
rlabel metal1 23000 24242 23000 24242 0 _0230_
rlabel metal1 22770 20978 22770 20978 0 _0231_
rlabel metal1 10718 22066 10718 22066 0 _0232_
rlabel metal1 22908 24378 22908 24378 0 _0233_
rlabel metal2 26450 23732 26450 23732 0 _0234_
rlabel metal1 11684 21114 11684 21114 0 _0235_
rlabel metal1 7084 17238 7084 17238 0 _0236_
rlabel metal2 5566 17612 5566 17612 0 _0237_
rlabel metal1 7636 18258 7636 18258 0 _0238_
rlabel metal1 6670 16422 6670 16422 0 _0239_
rlabel metal1 6164 20026 6164 20026 0 _0240_
rlabel metal1 7820 18802 7820 18802 0 _0241_
rlabel metal2 13570 4590 13570 4590 0 _0242_
rlabel metal1 13455 3570 13455 3570 0 _0243_
rlabel metal2 9890 17374 9890 17374 0 _0244_
rlabel metal2 10442 10302 10442 10302 0 _0245_
rlabel metal1 18216 3162 18216 3162 0 _0246_
rlabel via1 10534 15997 10534 15997 0 _0247_
rlabel metal2 16790 19992 16790 19992 0 _0248_
rlabel metal1 16422 15130 16422 15130 0 _0249_
rlabel metal1 16836 13226 16836 13226 0 _0250_
rlabel metal1 21965 21930 21965 21930 0 _0251_
rlabel metal1 17940 12954 17940 12954 0 _0252_
rlabel metal2 22310 7208 22310 7208 0 _0253_
rlabel metal2 13662 18258 13662 18258 0 _0254_
rlabel metal1 13846 20026 13846 20026 0 _0255_
rlabel metal2 13662 10302 13662 10302 0 _0256_
rlabel metal2 14490 18462 14490 18462 0 _0257_
rlabel metal1 13846 18394 13846 18394 0 _0258_
rlabel metal1 13018 6698 13018 6698 0 _0259_
rlabel metal1 19642 22984 19642 22984 0 _0260_
rlabel metal1 18952 22610 18952 22610 0 _0261_
rlabel metal2 19458 22372 19458 22372 0 _0262_
rlabel metal2 19182 23902 19182 23902 0 _0263_
rlabel metal1 18446 23290 18446 23290 0 _0264_
rlabel metal1 18308 12818 18308 12818 0 _0265_
rlabel metal2 16974 9248 16974 9248 0 _0266_
rlabel metal1 12857 13294 12857 13294 0 _0267_
rlabel metal2 21758 15640 21758 15640 0 _0268_
rlabel metal1 20792 6698 20792 6698 0 _0269_
rlabel metal1 13386 15062 13386 15062 0 _0270_
rlabel metal2 23046 5032 23046 5032 0 _0271_
rlabel metal2 16330 23664 16330 23664 0 _0272_
rlabel metal1 11408 23086 11408 23086 0 _0273_
rlabel metal2 10442 23324 10442 23324 0 _0274_
rlabel metal2 15778 22814 15778 22814 0 _0275_
rlabel metal1 12466 23084 12466 23084 0 _0276_
rlabel metal1 8970 24242 8970 24242 0 _0277_
rlabel metal1 16836 22406 16836 22406 0 _0278_
rlabel metal1 15502 14518 15502 14518 0 _0279_
rlabel metal1 14720 19482 14720 19482 0 _0280_
rlabel metal2 24702 23528 24702 23528 0 _0281_
rlabel metal1 14444 14042 14444 14042 0 _0282_
rlabel metal2 23414 5406 23414 5406 0 _0283_
rlabel metal1 9200 9418 9200 9418 0 _0284_
rlabel metal1 8096 11322 8096 11322 0 _0285_
rlabel metal1 12466 14484 12466 14484 0 _0286_
rlabel metal1 8510 11220 8510 11220 0 _0287_
rlabel metal1 8418 8058 8418 8058 0 _0288_
rlabel metal1 8418 15130 8418 15130 0 _0289_
rlabel metal1 12696 3706 12696 3706 0 _0290_
rlabel metal1 9292 3978 9292 3978 0 _0291_
rlabel metal1 13202 7276 13202 7276 0 _0292_
rlabel metal2 13754 5780 13754 5780 0 _0293_
rlabel metal1 10764 5338 10764 5338 0 _0294_
rlabel metal1 20240 6290 20240 6290 0 _0295_
rlabel metal1 13662 7752 13662 7752 0 _0296_
rlabel metal1 12972 5066 12972 5066 0 _0297_
rlabel metal1 9614 7854 9614 7854 0 _0298_
rlabel metal2 15778 6766 15778 6766 0 _0299_
rlabel metal1 10580 8466 10580 8466 0 _0300_
rlabel metal1 8280 8602 8280 8602 0 _0301_
rlabel metal1 12328 12886 12328 12886 0 _0302_
rlabel metal1 11454 10778 11454 10778 0 _0303_
rlabel metal1 18354 6970 18354 6970 0 _0304_
rlabel metal2 13754 10846 13754 10846 0 _0305_
rlabel metal1 11546 9146 11546 9146 0 _0306_
rlabel metal1 20286 5678 20286 5678 0 _0307_
rlabel metal1 14260 5338 14260 5338 0 _0308_
rlabel metal1 13892 4726 13892 4726 0 _0309_
rlabel metal1 22494 4250 22494 4250 0 _0310_
rlabel metal1 23460 4794 23460 4794 0 _0311_
rlabel metal2 12190 7548 12190 7548 0 _0312_
rlabel metal1 23874 5202 23874 5202 0 _0313_
rlabel metal1 11362 20230 11362 20230 0 _0314_
rlabel metal1 23138 22678 23138 22678 0 _0315_
rlabel metal2 16054 19652 16054 19652 0 _0316_
rlabel metal1 18308 19686 18308 19686 0 _0317_
rlabel metal1 16008 6630 16008 6630 0 _0318_
rlabel metal1 15548 18394 15548 18394 0 _0319_
rlabel metal1 16054 8602 16054 8602 0 _0320_
rlabel metal1 15824 16626 15824 16626 0 _0321_
rlabel metal1 9936 12954 9936 12954 0 _0322_
rlabel metal1 10672 21862 10672 21862 0 _0323_
rlabel metal1 12558 16456 12558 16456 0 _0324_
rlabel metal1 12650 21420 12650 21420 0 _0325_
rlabel metal1 13892 8058 13892 8058 0 _0326_
rlabel metal1 11408 17306 11408 17306 0 _0327_
rlabel metal1 14674 12104 14674 12104 0 _0328_
rlabel metal1 13340 14042 13340 14042 0 _0329_
rlabel metal1 6394 11322 6394 11322 0 _0330_
rlabel metal1 7636 13838 7636 13838 0 _0331_
rlabel metal1 6808 12410 6808 12410 0 _0332_
rlabel metal1 11040 13362 11040 13362 0 _0333_
rlabel metal1 16514 17782 16514 17782 0 _0334_
rlabel metal2 26082 5406 26082 5406 0 _0335_
rlabel metal1 18078 14314 18078 14314 0 _0336_
rlabel metal1 25300 6358 25300 6358 0 _0337_
rlabel metal1 5060 12954 5060 12954 0 _0338_
rlabel metal2 4922 14076 4922 14076 0 _0339_
rlabel metal2 6762 12988 6762 12988 0 _0340_
rlabel metal1 7820 13362 7820 13362 0 _0341_
rlabel metal2 12650 24582 12650 24582 0 _0342_
rlabel metal2 21390 25500 21390 25500 0 _0343_
rlabel metal1 14030 24378 14030 24378 0 _0344_
rlabel metal1 19090 25466 19090 25466 0 _0345_
rlabel metal1 25346 3162 25346 3162 0 _0346_
rlabel metal1 16606 11050 16606 11050 0 _0347_
rlabel metal2 25806 3740 25806 3740 0 _0348_
rlabel metal1 23138 23018 23138 23018 0 _0349_
rlabel metal2 18722 26282 18722 26282 0 _0350_
rlabel metal2 13938 24310 13938 24310 0 _0351_
rlabel metal1 18032 23698 18032 23698 0 _0352_
rlabel metal1 13294 23698 13294 23698 0 _0353_
rlabel metal1 14536 26418 14536 26418 0 _0354_
rlabel metal2 20746 26724 20746 26724 0 _0355_
rlabel metal2 16698 26588 16698 26588 0 _0356_
rlabel metal1 17894 26554 17894 26554 0 _0357_
rlabel metal1 7774 6664 7774 6664 0 _0358_
rlabel metal2 12466 16320 12466 16320 0 _0359_
rlabel metal1 8096 6358 8096 6358 0 _0360_
rlabel metal1 13846 8534 13846 8534 0 _0361_
rlabel metal2 11914 26248 11914 26248 0 _0362_
rlabel metal1 20654 24310 20654 24310 0 _0363_
rlabel metal2 13386 26078 13386 26078 0 _0364_
rlabel metal1 23230 25330 23230 25330 0 _0365_
rlabel metal2 11914 3604 11914 3604 0 _0366_
rlabel metal1 19182 3706 19182 3706 0 _0367_
rlabel metal2 15594 3876 15594 3876 0 _0368_
rlabel metal1 20562 2958 20562 2958 0 _0369_
rlabel metal2 14214 16728 14214 16728 0 _0370_
rlabel metal2 10626 7820 10626 7820 0 _0371_
rlabel metal1 15226 10710 15226 10710 0 _0372_
rlabel metal1 10764 6426 10764 6426 0 _0373_
rlabel metal1 20596 3434 20596 3434 0 _0374_
rlabel metal2 12742 7140 12742 7140 0 _0375_
rlabel metal1 17618 5576 17618 5576 0 _0376_
rlabel metal1 12006 8364 12006 8364 0 _0377_
rlabel metal2 5474 28373 5474 28373 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 3450 28373 3450 28373 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 1234 20468 1234 20468 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 28428 9554 28428 9554 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 29164 18734 29164 18734 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 18630 26996 18630 26996 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 7774 1588 7774 1588 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 11638 1588 11638 1588 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 24518 1588 24518 1588 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1740 748 1740 748 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 28382 23443 28382 23443 0 ccff_head
rlabel metal2 3266 1520 3266 1520 0 ccff_tail
rlabel metal2 25806 1588 25806 1588 0 chanx_left_in[0]
rlabel metal3 1234 24548 1234 24548 0 chanx_left_in[10]
rlabel metal1 26082 27472 26082 27472 0 chanx_left_in[11]
rlabel metal2 28382 14705 28382 14705 0 chanx_left_in[12]
rlabel metal1 9200 27438 9200 27438 0 chanx_left_in[13]
rlabel metal2 3174 27455 3174 27455 0 chanx_left_in[14]
rlabel metal3 1234 19788 1234 19788 0 chanx_left_in[15]
rlabel metal2 29026 1027 29026 1027 0 chanx_left_in[16]
rlabel metal3 1234 13668 1234 13668 0 chanx_left_in[17]
rlabel metal2 26910 26129 26910 26129 0 chanx_left_in[18]
rlabel via2 27002 3485 27002 3485 0 chanx_left_in[1]
rlabel metal1 20562 26962 20562 26962 0 chanx_left_in[2]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_in[3]
rlabel metal1 11500 27438 11500 27438 0 chanx_left_in[4]
rlabel metal1 12512 27438 12512 27438 0 chanx_left_in[5]
rlabel metal2 21942 28366 21942 28366 0 chanx_left_in[6]
rlabel metal3 1234 21828 1234 21828 0 chanx_left_in[7]
rlabel metal2 26266 27489 26266 27489 0 chanx_left_in[8]
rlabel metal1 28382 25840 28382 25840 0 chanx_left_in[9]
rlabel metal1 29118 27098 29118 27098 0 chanx_left_out[0]
rlabel via2 28290 6171 28290 6171 0 chanx_left_out[10]
rlabel metal1 18216 27574 18216 27574 0 chanx_left_out[11]
rlabel metal1 13616 27574 13616 27574 0 chanx_left_out[12]
rlabel metal3 1234 3468 1234 3468 0 chanx_left_out[13]
rlabel metal2 2806 28203 2806 28203 0 chanx_left_out[14]
rlabel metal2 6486 1520 6486 1520 0 chanx_left_out[15]
rlabel metal2 28290 21233 28290 21233 0 chanx_left_out[16]
rlabel metal2 27738 1520 27738 1520 0 chanx_left_out[17]
rlabel metal1 29118 10778 29118 10778 0 chanx_left_out[18]
rlabel metal1 16606 27574 16606 27574 0 chanx_left_out[1]
rlabel metal1 10488 27574 10488 27574 0 chanx_left_out[2]
rlabel metal3 28850 68 28850 68 0 chanx_left_out[3]
rlabel via2 28290 22491 28290 22491 0 chanx_left_out[4]
rlabel metal1 28474 26554 28474 26554 0 chanx_left_out[5]
rlabel metal3 1234 4828 1234 4828 0 chanx_left_out[6]
rlabel metal2 10350 1520 10350 1520 0 chanx_left_out[7]
rlabel metal2 28290 4913 28290 4913 0 chanx_left_out[8]
rlabel metal3 1234 17068 1234 17068 0 chanx_left_out[9]
rlabel metal3 1924 2108 1924 2108 0 chany_bottom_in[0]
rlabel metal3 1234 23188 1234 23188 0 chany_bottom_in[10]
rlabel metal2 8050 28373 8050 28373 0 chany_bottom_in[11]
rlabel metal2 21942 1095 21942 1095 0 chany_bottom_in[12]
rlabel metal1 26910 27438 26910 27438 0 chany_bottom_in[13]
rlabel metal2 18722 1078 18722 1078 0 chany_bottom_in[14]
rlabel metal2 1978 1588 1978 1588 0 chany_bottom_in[15]
rlabel metal3 1234 14348 1234 14348 0 chany_bottom_in[16]
rlabel metal2 26450 1588 26450 1588 0 chany_bottom_in[17]
rlabel metal3 28850 12308 28850 12308 0 chany_bottom_in[18]
rlabel metal1 29164 6766 29164 6766 0 chany_bottom_in[1]
rlabel metal1 20654 3060 20654 3060 0 chany_bottom_in[2]
rlabel metal3 1234 25908 1234 25908 0 chany_bottom_in[3]
rlabel metal2 25438 1921 25438 1921 0 chany_bottom_in[4]
rlabel metal2 4140 27438 4140 27438 0 chany_bottom_in[5]
rlabel metal2 28382 9809 28382 9809 0 chany_bottom_in[6]
rlabel metal3 1234 12308 1234 12308 0 chany_bottom_in[7]
rlabel metal2 23230 1588 23230 1588 0 chany_bottom_in[8]
rlabel via2 28382 19805 28382 19805 0 chany_bottom_in[9]
rlabel metal2 13570 1520 13570 1520 0 chany_bottom_out[0]
rlabel metal3 1234 18428 1234 18428 0 chany_bottom_out[10]
rlabel metal2 14858 1027 14858 1027 0 chany_bottom_out[11]
rlabel metal2 46 1520 46 1520 0 chany_bottom_out[12]
rlabel metal2 17434 1520 17434 1520 0 chany_bottom_out[13]
rlabel metal3 1234 6188 1234 6188 0 chany_bottom_out[14]
rlabel metal2 15134 28441 15134 28441 0 chany_bottom_out[15]
rlabel metal3 1234 9588 1234 9588 0 chany_bottom_out[16]
rlabel metal1 1794 27574 1794 27574 0 chany_bottom_out[17]
rlabel metal2 4554 1520 4554 1520 0 chany_bottom_out[18]
rlabel metal2 690 1792 690 1792 0 chany_bottom_out[1]
rlabel metal1 27876 27574 27876 27574 0 chany_bottom_out[2]
rlabel metal1 20838 27574 20838 27574 0 chany_bottom_out[3]
rlabel metal2 12926 1520 12926 1520 0 chany_bottom_out[4]
rlabel metal2 27554 27370 27554 27370 0 chany_bottom_out[5]
rlabel metal1 29118 3366 29118 3366 0 chany_bottom_out[6]
rlabel metal3 1234 6868 1234 6868 0 chany_bottom_out[7]
rlabel metal2 28290 15793 28290 15793 0 chany_bottom_out[8]
rlabel metal2 5842 1520 5842 1520 0 chany_bottom_out[9]
rlabel metal2 9062 1588 9062 1588 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal3 1234 10948 1234 10948 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 28382 17119 28382 17119 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 16146 1588 16146 1588 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 25438 27404 25438 27404 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24748 27438 24748 27438 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 2254 26962 2254 26962 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 6762 28373 6762 28373 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 20424 2890 20424 2890 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 8228 1234 8228 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 18998 3060 18998 3060 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 13524 8942 13524 8942 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 12742 10336 12742 10336 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal2 21206 10387 21206 10387 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal2 24978 20468 24978 20468 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal2 10442 14433 10442 14433 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal1 14398 5678 14398 5678 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal2 21482 23817 21482 23817 0 mem_bottom_track_15.DFFR_0_.Q
rlabel via2 21574 15691 21574 15691 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal2 14398 21794 14398 21794 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 24058 21454 24058 21454 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 17986 18326 17986 18326 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal2 21482 17034 21482 17034 0 mem_bottom_track_19.DFFR_1_.Q
rlabel metal1 21988 17578 21988 17578 0 mem_bottom_track_21.DFFR_0_.Q
rlabel metal1 20368 21114 20368 21114 0 mem_bottom_track_21.DFFR_1_.Q
rlabel metal1 19872 17578 19872 17578 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal2 21206 16048 21206 16048 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal2 20746 19686 20746 19686 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 19642 16626 19642 16626 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 20838 16422 20838 16422 0 mem_bottom_track_27.DFFR_0_.Q
rlabel via1 20470 15861 20470 15861 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal1 19596 13838 19596 13838 0 mem_bottom_track_29.DFFR_0_.Q
rlabel metal1 18344 13702 18344 13702 0 mem_bottom_track_29.DFFR_1_.Q
rlabel metal1 15226 12818 15226 12818 0 mem_bottom_track_3.DFFR_0_.Q
rlabel metal1 14582 13362 14582 13362 0 mem_bottom_track_3.DFFR_1_.Q
rlabel metal1 20286 14042 20286 14042 0 mem_bottom_track_31.DFFR_0_.Q
rlabel metal1 19688 15402 19688 15402 0 mem_bottom_track_31.DFFR_1_.Q
rlabel metal1 21804 13226 21804 13226 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal2 18170 13549 18170 13549 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal1 19228 19278 19228 19278 0 mem_bottom_track_35.DFFR_0_.Q
rlabel metal2 19918 19261 19918 19261 0 mem_bottom_track_35.DFFR_1_.Q
rlabel metal1 13754 17782 13754 17782 0 mem_bottom_track_37.DFFR_0_.Q
rlabel metal1 13064 4590 13064 4590 0 mem_bottom_track_37.DFFR_1_.Q
rlabel metal1 14168 21522 14168 21522 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal1 23828 15130 23828 15130 0 mem_bottom_track_5.DFFR_1_.Q
rlabel metal1 13570 18190 13570 18190 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal1 19274 23800 19274 23800 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal1 12742 11118 12742 11118 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal1 17710 12818 17710 12818 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 26358 10234 26358 10234 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 15410 23120 15410 23120 0 mem_left_track_11.DFFR_0_.D
rlabel metal2 14858 14654 14858 14654 0 mem_left_track_11.DFFR_0_.Q
rlabel metal1 17986 20978 17986 20978 0 mem_left_track_11.DFFR_1_.Q
rlabel metal1 13570 11220 13570 11220 0 mem_left_track_13.DFFR_0_.Q
rlabel metal1 13846 11696 13846 11696 0 mem_left_track_13.DFFR_1_.Q
rlabel metal1 20838 12716 20838 12716 0 mem_left_track_15.DFFR_0_.Q
rlabel metal2 20562 9180 20562 9180 0 mem_left_track_15.DFFR_1_.Q
rlabel metal2 9338 8721 9338 8721 0 mem_left_track_17.DFFR_0_.Q
rlabel metal1 19642 8398 19642 8398 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 21206 11526 21206 11526 0 mem_left_track_19.DFFR_0_.Q
rlabel metal1 20562 9486 20562 9486 0 mem_left_track_19.DFFR_1_.Q
rlabel metal2 18078 11526 18078 11526 0 mem_left_track_21.DFFR_0_.Q
rlabel metal2 23782 17204 23782 17204 0 mem_left_track_21.DFFR_1_.Q
rlabel via2 18170 20587 18170 20587 0 mem_left_track_23.DFFR_0_.Q
rlabel metal1 21436 19958 21436 19958 0 mem_left_track_23.DFFR_1_.Q
rlabel metal2 18262 21012 18262 21012 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 17802 26928 17802 26928 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 19734 13379 19734 13379 0 mem_left_track_27.DFFR_0_.Q
rlabel metal2 12466 7038 12466 7038 0 mem_left_track_27.DFFR_1_.Q
rlabel metal2 21942 16830 21942 16830 0 mem_left_track_29.DFFR_0_.Q
rlabel metal1 19872 16966 19872 16966 0 mem_left_track_29.DFFR_1_.Q
rlabel metal2 13938 8636 13938 8636 0 mem_left_track_3.DFFR_0_.Q
rlabel metal1 13892 18734 13892 18734 0 mem_left_track_3.DFFR_1_.Q
rlabel metal2 19734 7871 19734 7871 0 mem_left_track_31.DFFR_0_.Q
rlabel metal1 15502 3536 15502 3536 0 mem_left_track_31.DFFR_1_.Q
rlabel metal2 19366 8126 19366 8126 0 mem_left_track_33.DFFR_0_.Q
rlabel metal1 23092 11186 23092 11186 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 12604 6766 12604 6766 0 mem_left_track_35.DFFR_0_.Q
rlabel metal2 20930 8602 20930 8602 0 mem_left_track_35.DFFR_1_.Q
rlabel metal2 13478 5712 13478 5712 0 mem_left_track_37.DFFR_0_.Q
rlabel metal1 18354 14926 18354 14926 0 mem_left_track_5.DFFR_0_.Q
rlabel metal1 20240 15130 20240 15130 0 mem_left_track_5.DFFR_1_.Q
rlabel metal2 26818 6222 26818 6222 0 mem_left_track_7.DFFR_0_.Q
rlabel metal2 17802 9044 17802 9044 0 mem_left_track_7.DFFR_1_.Q
rlabel metal2 12328 20332 12328 20332 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 13662 15062 13662 15062 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 15502 13362 15502 13362 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 27600 4046 27600 4046 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 16928 13770 16928 13770 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 19182 6800 19182 6800 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16836 7786 16836 7786 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 14858 2992 14858 2992 0 mux_bottom_track_1.out
rlabel metal1 14398 12750 14398 12750 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal1 16054 6732 16054 6732 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal1 23736 24786 23736 24786 0 mux_bottom_track_11.INVTX1_2_.out
rlabel metal1 16468 12750 16468 12750 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23276 24582 23276 24582 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24886 24378 24886 24378 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 27278 25364 27278 25364 0 mux_bottom_track_11.out
rlabel metal1 8050 13294 8050 13294 0 mux_bottom_track_13.INVTX1_1_.out
rlabel metal1 7866 15538 7866 15538 0 mux_bottom_track_13.INVTX1_2_.out
rlabel metal2 17434 6528 17434 6528 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13202 12648 13202 12648 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18078 6154 18078 6154 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 27784 3502 27784 3502 0 mux_bottom_track_13.out
rlabel metal1 14030 25704 14030 25704 0 mux_bottom_track_15.INVTX1_1_.out
rlabel metal1 20286 20332 20286 20332 0 mux_bottom_track_15.INVTX1_2_.out
rlabel metal1 11132 15674 11132 15674 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13432 21046 13432 21046 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 1610 9010 1610 9010 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 1794 8636 1794 8636 0 mux_bottom_track_15.out
rlabel metal2 7406 21794 7406 21794 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal2 26082 24412 26082 24412 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal2 12650 21726 12650 21726 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 22770 24174 22770 24174 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24104 24650 24104 24650 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 28198 24990 28198 24990 0 mux_bottom_track_17.out
rlabel metal2 5106 20162 5106 20162 0 mux_bottom_track_19.INVTX1_2_.out
rlabel metal2 8326 18496 8326 18496 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 5750 18632 5750 18632 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 7590 17102 7590 17102 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 5750 3468 5750 3468 0 mux_bottom_track_19.out
rlabel metal2 22954 23052 22954 23052 0 mux_bottom_track_21.INVTX1_1_.out
rlabel metal1 16100 19890 16100 19890 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 13294 19618 13294 19618 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 7958 17578 7958 17578 0 mux_bottom_track_21.out
rlabel metal2 15134 21182 15134 21182 0 mux_bottom_track_23.INVTX1_0_.out
rlabel via2 15962 18819 15962 18819 0 mux_bottom_track_23.INVTX1_1_.out
rlabel metal1 16422 18598 16422 18598 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18078 7922 18078 7922 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17066 3468 17066 3468 0 mux_bottom_track_23.out
rlabel metal1 13892 21998 13892 21998 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 11086 22474 11086 22474 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal2 12466 18428 12466 18428 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12926 16660 12926 16660 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4738 5712 4738 5712 0 mux_bottom_track_25.out
rlabel metal1 12834 15470 12834 15470 0 mux_bottom_track_27.INVTX1_0_.out
rlabel metal1 10994 18802 10994 18802 0 mux_bottom_track_27.INVTX1_1_.out
rlabel metal1 13432 15334 13432 15334 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15916 9962 15916 9962 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 17618 3264 17618 3264 0 mux_bottom_track_27.out
rlabel metal2 6578 14892 6578 14892 0 mux_bottom_track_29.INVTX1_1_.out
rlabel metal1 8188 13702 8188 13702 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 6854 13430 6854 13430 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 5934 9146 5934 9146 0 mux_bottom_track_29.out
rlabel metal2 21160 21964 21160 21964 0 mux_bottom_track_3.INVTX1_2_.out
rlabel metal2 16974 14722 16974 14722 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15226 19040 15226 19040 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17618 14008 17618 14008 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6578 4590 6578 4590 0 mux_bottom_track_3.out
rlabel metal2 27646 4964 27646 4964 0 mux_bottom_track_31.INVTX1_1_.out
rlabel via3 16491 13804 16491 13804 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17250 16320 17250 16320 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14582 25296 14582 25296 0 mux_bottom_track_31.out
rlabel metal1 3772 13498 3772 13498 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal1 6532 12818 6532 12818 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 5888 12682 5888 12682 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4370 9554 4370 9554 0 mux_bottom_track_33.out
rlabel metal1 21206 25364 21206 25364 0 mux_bottom_track_35.INVTX1_1_.out
rlabel metal1 18952 25738 18952 25738 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15778 25058 15778 25058 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 4278 26758 4278 26758 0 mux_bottom_track_35.out
rlabel metal2 19274 3944 19274 3944 0 mux_bottom_track_37.INVTX1_2_.out
rlabel metal2 10994 15385 10994 15385 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 14766 4216 14766 4216 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12466 3383 12466 3383 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 9292 3026 9292 3026 0 mux_bottom_track_37.out
rlabel metal2 9338 18292 9338 18292 0 mux_bottom_track_5.INVTX1_2_.out
rlabel metal1 16790 21590 16790 21590 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15594 21386 15594 21386 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21022 22287 21022 22287 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 25438 25058 25438 25058 0 mux_bottom_track_5.out
rlabel metal2 13202 25092 13202 25092 0 mux_bottom_track_7.INVTX1_2_.out
rlabel metal1 15180 22066 15180 22066 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13892 24582 13892 24582 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15640 23766 15640 23766 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 21574 26826 21574 26826 0 mux_bottom_track_7.out
rlabel metal1 12098 21318 12098 21318 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal2 13478 11968 13478 11968 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12834 15946 12834 15946 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 13984 13838 13984 13838 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 11086 4318 11086 4318 0 mux_bottom_track_9.out
rlabel metal1 21850 6664 21850 6664 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 18538 13226 18538 13226 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 16836 13362 16836 13362 0 mux_left_track_1.INVTX1_2_.out
rlabel metal3 19941 16660 19941 16660 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17526 17918 17526 17918 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21942 19839 21942 19839 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 27830 24378 27830 24378 0 mux_left_track_1.out
rlabel metal1 26634 4726 26634 4726 0 mux_left_track_11.INVTX1_0_.out
rlabel metal2 12466 24684 12466 24684 0 mux_left_track_11.INVTX1_1_.out
rlabel metal1 16974 14926 16974 14926 0 mux_left_track_11.INVTX1_2_.out
rlabel via3 23805 6868 23805 6868 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17066 14790 17066 14790 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 19642 21250 19642 21250 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 27922 26180 27922 26180 0 mux_left_track_11.out
rlabel metal1 6256 15538 6256 15538 0 mux_left_track_13.INVTX1_0_.out
rlabel metal1 11960 8942 11960 8942 0 mux_left_track_13.INVTX1_2_.out
rlabel metal2 9982 15130 9982 15130 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9338 11186 9338 11186 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 9706 11390 9706 11390 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6808 7854 6808 7854 0 mux_left_track_13.out
rlabel metal2 19642 6052 19642 6052 0 mux_left_track_15.INVTX1_0_.out
rlabel metal2 12558 5984 12558 5984 0 mux_left_track_15.INVTX1_2_.out
rlabel metal1 13800 6290 13800 6290 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12190 5236 12190 5236 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 13110 4420 13110 4420 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 10442 3060 10442 3060 0 mux_left_track_15.out
rlabel metal1 8924 9010 8924 9010 0 mux_left_track_17.INVTX1_0_.out
rlabel metal1 12926 10030 12926 10030 0 mux_left_track_17.INVTX1_2_.out
rlabel metal2 11270 8364 11270 8364 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14444 9078 14444 9078 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17434 7446 17434 7446 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 26634 6086 26634 6086 0 mux_left_track_17.out
rlabel metal2 22402 4896 22402 4896 0 mux_left_track_19.INVTX1_0_.out
rlabel metal1 18354 7378 18354 7378 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12788 12750 12788 12750 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 13018 12954 13018 12954 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 5658 16524 5658 16524 0 mux_left_track_19.out
rlabel metal1 25714 21658 25714 21658 0 mux_left_track_21.INVTX1_0_.out
rlabel metal4 17756 8160 17756 8160 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 26220 4794 26220 4794 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27278 6086 27278 6086 0 mux_left_track_21.out
rlabel metal2 13018 24106 13018 24106 0 mux_left_track_23.INVTX1_0_.out
rlabel metal1 13708 19278 13708 19278 0 mux_left_track_23.INVTX1_1_.out
rlabel metal2 14950 23392 14950 23392 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 18906 24718 18906 24718 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 19918 26554 19918 26554 0 mux_left_track_23.out
rlabel metal1 14950 26962 14950 26962 0 mux_left_track_25.INVTX1_0_.out
rlabel metal1 23092 15538 23092 15538 0 mux_left_track_25.INVTX1_1_.out
rlabel metal1 17112 26350 17112 26350 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16284 26486 16284 26486 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14536 26010 14536 26010 0 mux_left_track_25.out
rlabel metal2 20194 6222 20194 6222 0 mux_left_track_27.INVTX1_0_.out
rlabel metal1 13202 14960 13202 14960 0 mux_left_track_27.INVTX1_1_.out
rlabel metal1 14582 14926 14582 14926 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 8694 7276 8694 7276 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 4186 5644 4186 5644 0 mux_left_track_27.out
rlabel metal1 23966 25262 23966 25262 0 mux_left_track_29.INVTX1_0_.out
rlabel metal1 18814 25398 18814 25398 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13570 25772 13570 25772 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5060 26010 5060 26010 0 mux_left_track_29.out
rlabel metal1 9706 9146 9706 9146 0 mux_left_track_3.INVTX1_0_.out
rlabel metal1 14628 11322 14628 11322 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 14398 19856 14398 19856 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 19044 21318 19044 21318 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 17986 25262 17986 25262 0 mux_left_track_3.out
rlabel metal1 19642 2618 19642 2618 0 mux_left_track_31.INVTX1_0_.out
rlabel metal1 19780 4726 19780 4726 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14145 3978 14145 3978 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 11178 2992 11178 2992 0 mux_left_track_31.out
rlabel metal1 11592 6970 11592 6970 0 mux_left_track_33.INVTX1_0_.out
rlabel metal1 12972 9146 12972 9146 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15502 17272 15502 17272 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23736 21046 23736 21046 0 mux_left_track_33.out
rlabel metal1 9752 13974 9752 13974 0 mux_left_track_35.INVTX1_0_.out
rlabel metal2 13202 6018 13202 6018 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 21206 4590 21206 4590 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24702 3026 24702 3026 0 mux_left_track_35.out
rlabel metal2 24702 4692 24702 4692 0 mux_left_track_37.INVTX1_0_.out
rlabel metal2 22954 5644 22954 5644 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15088 6426 15088 6426 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 20378 6120 20378 6120 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 27968 7514 27968 7514 0 mux_left_track_37.out
rlabel metal1 18262 12716 18262 12716 0 mux_left_track_5.INVTX1_0_.out
rlabel metal1 19366 12750 19366 12750 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel via1 19550 23035 19550 23035 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 19550 23681 19550 23681 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 14582 26316 14582 26316 0 mux_left_track_5.out
rlabel metal1 20792 4794 20792 4794 0 mux_left_track_7.INVTX1_0_.out
rlabel metal1 20562 6698 20562 6698 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13800 13498 13800 13498 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21298 8262 21298 8262 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 25898 4794 25898 4794 0 mux_left_track_7.out
rlabel metal2 9246 24004 9246 24004 0 mux_left_track_9.INVTX1_0_.out
rlabel metal2 14030 22916 14030 22916 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14674 23018 14674 23018 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 16882 22848 16882 22848 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 28106 20876 28106 20876 0 mux_left_track_9.out
rlabel metal1 7314 25874 7314 25874 0 net1
rlabel metal2 3910 4386 3910 4386 0 net10
rlabel metal1 18400 4658 18400 4658 0 net100
rlabel metal2 14306 17136 14306 17136 0 net101
rlabel metal2 9890 20604 9890 20604 0 net102
rlabel metal1 11914 24718 11914 24718 0 net103
rlabel metal2 12282 18428 12282 18428 0 net104
rlabel metal1 21850 26962 21850 26962 0 net105
rlabel metal1 8418 12750 8418 12750 0 net106
rlabel metal1 12834 20910 12834 20910 0 net107
rlabel metal1 21850 20570 21850 20570 0 net108
rlabel metal2 5382 17340 5382 17340 0 net109
rlabel metal1 27416 23494 27416 23494 0 net11
rlabel metal1 14766 3502 14766 3502 0 net110
rlabel metal1 16514 16014 16514 16014 0 net111
rlabel metal1 13708 20434 13708 20434 0 net112
rlabel metal1 20792 21658 20792 21658 0 net113
rlabel metal2 11822 13668 11822 13668 0 net114
rlabel metal1 11224 23154 11224 23154 0 net115
rlabel metal1 15640 14042 15640 14042 0 net116
rlabel metal2 8326 11220 8326 11220 0 net117
rlabel metal1 11316 4590 11316 4590 0 net118
rlabel metal1 13938 7922 13938 7922 0 net119
rlabel metal1 24610 3094 24610 3094 0 net12
rlabel metal2 11730 11900 11730 11900 0 net120
rlabel metal1 14812 5338 14812 5338 0 net121
rlabel metal2 12650 19516 12650 19516 0 net122
rlabel metal1 18170 7514 18170 7514 0 net123
rlabel metal1 10074 12886 10074 12886 0 net124
rlabel metal1 14858 9962 14858 9962 0 net125
rlabel metal1 5244 12206 5244 12206 0 net126
rlabel metal2 16974 18802 16974 18802 0 net127
rlabel metal2 4278 13124 4278 13124 0 net128
rlabel metal1 10672 24242 10672 24242 0 net129
rlabel metal1 4600 19822 4600 19822 0 net13
rlabel metal2 23966 4420 23966 4420 0 net130
rlabel metal1 19090 25874 19090 25874 0 net131
rlabel metal1 14720 26350 14720 26350 0 net132
rlabel metal1 8050 7310 8050 7310 0 net133
rlabel metal2 11822 26418 11822 26418 0 net134
rlabel metal2 11730 4284 11730 4284 0 net135
rlabel metal1 14812 16218 14812 16218 0 net136
rlabel metal1 21206 3570 21206 3570 0 net137
rlabel metal1 24656 23698 24656 23698 0 net14
rlabel metal1 28336 14586 28336 14586 0 net15
rlabel metal1 10074 22610 10074 22610 0 net16
rlabel metal1 6624 26758 6624 26758 0 net17
rlabel metal2 3726 17884 3726 17884 0 net18
rlabel metal1 27508 3162 27508 3162 0 net19
rlabel metal1 5290 27506 5290 27506 0 net2
rlabel metal2 3266 13668 3266 13668 0 net20
rlabel metal1 26174 25874 26174 25874 0 net21
rlabel metal1 27324 3706 27324 3706 0 net22
rlabel metal1 20930 23086 20930 23086 0 net23
rlabel metal1 2185 15946 2185 15946 0 net24
rlabel metal1 11684 25262 11684 25262 0 net25
rlabel metal2 12742 26826 12742 26826 0 net26
rlabel metal1 23782 26996 23782 26996 0 net27
rlabel metal2 8786 21148 8786 21148 0 net28
rlabel metal2 25898 25636 25898 25636 0 net29
rlabel metal2 4002 18734 4002 18734 0 net3
rlabel metal1 27324 24786 27324 24786 0 net30
rlabel metal1 2990 2924 2990 2924 0 net31
rlabel metal2 10718 24174 10718 24174 0 net32
rlabel metal1 14306 27472 14306 27472 0 net33
rlabel metal1 20102 4080 20102 4080 0 net34
rlabel metal1 24426 26996 24426 26996 0 net35
rlabel metal1 19918 2448 19918 2448 0 net36
rlabel metal1 2346 2312 2346 2312 0 net37
rlabel metal1 1610 14280 1610 14280 0 net38
rlabel metal1 26588 2618 26588 2618 0 net39
rlabel metal1 26266 13158 26266 13158 0 net4
rlabel metal2 28198 9996 28198 9996 0 net40
rlabel metal1 27646 6766 27646 6766 0 net41
rlabel metal1 20746 4590 20746 4590 0 net42
rlabel metal1 2185 26554 2185 26554 0 net43
rlabel metal1 26266 2550 26266 2550 0 net44
rlabel metal1 5060 27574 5060 27574 0 net45
rlabel metal1 23046 5678 23046 5678 0 net46
rlabel metal1 2852 12614 2852 12614 0 net47
rlabel metal1 22816 2550 22816 2550 0 net48
rlabel metal2 28198 20740 28198 20740 0 net49
rlabel metal1 28106 18938 28106 18938 0 net5
rlabel metal1 9246 2618 9246 2618 0 net50
rlabel metal2 1610 11492 1610 11492 0 net51
rlabel metal2 28014 15980 28014 15980 0 net52
rlabel metal1 16514 5202 16514 5202 0 net53
rlabel metal1 22310 23664 22310 23664 0 net54
rlabel metal1 23966 27438 23966 27438 0 net55
rlabel metal2 8326 24956 8326 24956 0 net56
rlabel metal2 12006 26860 12006 26860 0 net57
rlabel metal1 20470 2380 20470 2380 0 net58
rlabel metal2 8372 7990 8372 7990 0 net59
rlabel metal2 16146 25500 16146 25500 0 net6
rlabel metal2 1886 25024 1886 25024 0 net60
rlabel metal1 3174 2448 3174 2448 0 net61
rlabel metal2 27554 26486 27554 26486 0 net62
rlabel metal1 28106 6324 28106 6324 0 net63
rlabel metal1 18814 27438 18814 27438 0 net64
rlabel metal2 13202 27268 13202 27268 0 net65
rlabel metal2 4002 4250 4002 4250 0 net66
rlabel metal1 1610 26928 1610 26928 0 net67
rlabel metal1 7130 2414 7130 2414 0 net68
rlabel metal2 24610 21726 24610 21726 0 net69
rlabel metal1 8464 2618 8464 2618 0 net7
rlabel metal1 26358 2822 26358 2822 0 net70
rlabel metal2 28106 9622 28106 9622 0 net71
rlabel metal1 17250 25466 17250 25466 0 net72
rlabel metal1 14352 25670 14352 25670 0 net73
rlabel metal2 28106 3740 28106 3740 0 net74
rlabel metal1 28014 22610 28014 22610 0 net75
rlabel metal1 28106 26384 28106 26384 0 net76
rlabel metal1 1610 5236 1610 5236 0 net77
rlabel metal1 10350 2822 10350 2822 0 net78
rlabel metal2 28106 5644 28106 5644 0 net79
rlabel metal1 11454 2618 11454 2618 0 net8
rlabel metal1 5336 16762 5336 16762 0 net80
rlabel metal1 14076 2414 14076 2414 0 net81
rlabel metal1 7314 17850 7314 17850 0 net82
rlabel metal1 15364 2414 15364 2414 0 net83
rlabel metal1 1610 2482 1610 2482 0 net84
rlabel metal1 17204 3366 17204 3366 0 net85
rlabel metal1 1610 6324 1610 6324 0 net86
rlabel metal2 14398 26452 14398 26452 0 net87
rlabel metal2 3634 9860 3634 9860 0 net88
rlabel metal1 3588 27098 3588 27098 0 net89
rlabel metal2 24610 4148 24610 4148 0 net9
rlabel metal1 5106 2414 5106 2414 0 net90
rlabel metal1 1610 3060 1610 3060 0 net91
rlabel metal1 26358 25466 26358 25466 0 net92
rlabel metal2 21390 26996 21390 26996 0 net93
rlabel metal1 12512 2414 12512 2414 0 net94
rlabel metal2 27370 26758 27370 26758 0 net95
rlabel metal1 28106 3468 28106 3468 0 net96
rlabel metal2 1610 7820 1610 7820 0 net97
rlabel metal1 28336 16082 28336 16082 0 net98
rlabel metal1 5658 2822 5658 2822 0 net99
rlabel metal3 1188 27268 1188 27268 0 pReset
rlabel metal1 18032 20434 18032 20434 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
