VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2810.000 BY 2950.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 2946.000 1024.330 2950.000 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 0.000 2241.490 4.000 ;
    END
  END clk
  PIN gfpga_pad_GPIO_PAD_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.150 0.000 2489.430 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[0]
  PIN gfpga_pad_GPIO_PAD_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[10]
  PIN gfpga_pad_GPIO_PAD_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 2946.000 1272.270 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[11]
  PIN gfpga_pad_GPIO_PAD_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 98.640 2810.000 99.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[12]
  PIN gfpga_pad_GPIO_PAD_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2553.440 2810.000 2554.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[13]
  PIN gfpga_pad_GPIO_PAD_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2769.290 2946.000 2769.570 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[14]
  PIN gfpga_pad_GPIO_PAD_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 2946.000 1687.650 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[15]
  PIN gfpga_pad_GPIO_PAD_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[16]
  PIN gfpga_pad_GPIO_PAD_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[17]
  PIN gfpga_pad_GPIO_PAD_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[18]
  PIN gfpga_pad_GPIO_PAD_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[19]
  PIN gfpga_pad_GPIO_PAD_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 2946.000 1439.710 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[1]
  PIN gfpga_pad_GPIO_PAD_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 2946.000 277.290 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[20]
  PIN gfpga_pad_GPIO_PAD_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2291.640 2810.000 2292.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[21]
  PIN gfpga_pad_GPIO_PAD_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2104.640 4.000 2105.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[22]
  PIN gfpga_pad_GPIO_PAD_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2380.040 2810.000 2380.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[23]
  PIN gfpga_pad_GPIO_PAD_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[24]
  PIN gfpga_pad_GPIO_PAD_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.850 2946.000 2602.130 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[25]
  PIN gfpga_pad_GPIO_PAD_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 2946.000 1855.090 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[26]
  PIN gfpga_pad_GPIO_PAD_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 2946.000 361.010 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[27]
  PIN gfpga_pad_GPIO_PAD_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 2946.000 1355.990 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[28]
  PIN gfpga_pad_GPIO_PAD_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2366.440 4.000 2367.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[29]
  PIN gfpga_pad_GPIO_PAD_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1152.640 2810.000 1153.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[2]
  PIN gfpga_pad_GPIO_PAD_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[30]
  PIN gfpga_pad_GPIO_PAD_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 10.240 2810.000 10.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[31]
  PIN gfpga_pad_GPIO_PAD_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 2946.000 109.850 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[32]
  PIN gfpga_pad_GPIO_PAD_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[33]
  PIN gfpga_pad_GPIO_PAD_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1241.040 2810.000 1241.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[34]
  PIN gfpga_pad_GPIO_PAD_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[35]
  PIN gfpga_pad_GPIO_PAD_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[36]
  PIN gfpga_pad_GPIO_PAD_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 2946.000 441.510 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[37]
  PIN gfpga_pad_GPIO_PAD_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 2946.000 1523.430 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[38]
  PIN gfpga_pad_GPIO_PAD_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 2946.000 2354.190 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[39]
  PIN gfpga_pad_GPIO_PAD_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1764.640 2810.000 1765.240 ;
    END
  END gfpga_pad_GPIO_PAD_in[3]
  PIN gfpga_pad_GPIO_PAD_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1853.040 2810.000 1853.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[40]
  PIN gfpga_pad_GPIO_PAD_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 2946.000 608.950 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[41]
  PIN gfpga_pad_GPIO_PAD_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 2946.000 2270.470 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[42]
  PIN gfpga_pad_GPIO_PAD_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 0.000 1742.390 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[43]
  PIN gfpga_pad_GPIO_PAD_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[44]
  PIN gfpga_pad_GPIO_PAD_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2029.840 2810.000 2030.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[45]
  PIN gfpga_pad_GPIO_PAD_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2740.310 0.000 2740.590 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[46]
  PIN gfpga_pad_GPIO_PAD_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.430 0.000 2405.710 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[47]
  PIN gfpga_pad_GPIO_PAD_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1326.040 2810.000 1326.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[48]
  PIN gfpga_pad_GPIO_PAD_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.410 2946.000 2434.690 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[49]
  PIN gfpga_pad_GPIO_PAD_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[4]
  PIN gfpga_pad_GPIO_PAD_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 887.440 2810.000 888.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[50]
  PIN gfpga_pad_GPIO_PAD_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[51]
  PIN gfpga_pad_GPIO_PAD_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[52]
  PIN gfpga_pad_GPIO_PAD_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 802.440 2810.000 803.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[53]
  PIN gfpga_pad_GPIO_PAD_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 2946.000 940.610 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[54]
  PIN gfpga_pad_GPIO_PAD_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[55]
  PIN gfpga_pad_GPIO_PAD_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[56]
  PIN gfpga_pad_GPIO_PAD_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 363.840 2810.000 364.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[57]
  PIN gfpga_pad_GPIO_PAD_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.770 0.000 2074.050 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[58]
  PIN gfpga_pad_GPIO_PAD_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2203.240 2810.000 2203.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[59]
  PIN gfpga_pad_GPIO_PAD_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END gfpga_pad_GPIO_PAD_in[5]
  PIN gfpga_pad_GPIO_PAD_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[60]
  PIN gfpga_pad_GPIO_PAD_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[61]
  PIN gfpga_pad_GPIO_PAD_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.570 2946.000 2685.850 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[62]
  PIN gfpga_pad_GPIO_PAD_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END gfpga_pad_GPIO_PAD_in[63]
  PIN gfpga_pad_GPIO_PAD_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[6]
  PIN gfpga_pad_GPIO_PAD_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1591.240 2810.000 1591.840 ;
    END
  END gfpga_pad_GPIO_PAD_in[7]
  PIN gfpga_pad_GPIO_PAD_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 2946.000 692.670 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_in[8]
  PIN gfpga_pad_GPIO_PAD_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2907.040 2810.000 2907.640 ;
    END
  END gfpga_pad_GPIO_PAD_in[9]
  PIN gfpga_pad_GPIO_PAD_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2016.240 4.000 2016.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[0]
  PIN gfpga_pad_GPIO_PAD_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[10]
  PIN gfpga_pad_GPIO_PAD_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 2946.000 193.570 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[11]
  PIN gfpga_pad_GPIO_PAD_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 2946.000 856.890 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[12]
  PIN gfpga_pad_GPIO_PAD_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 2946.000 1108.050 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[13]
  PIN gfpga_pad_GPIO_PAD_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2189.640 4.000 2190.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[14]
  PIN gfpga_pad_GPIO_PAD_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[15]
  PIN gfpga_pad_GPIO_PAD_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 975.840 2810.000 976.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[16]
  PIN gfpga_pad_GPIO_PAD_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2730.240 2810.000 2730.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[17]
  PIN gfpga_pad_GPIO_PAD_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[18]
  PIN gfpga_pad_GPIO_PAD_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 187.040 2810.000 187.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[19]
  PIN gfpga_pad_GPIO_PAD_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1064.240 2810.000 1064.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[1]
  PIN gfpga_pad_GPIO_PAD_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 2946.000 1938.810 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[20]
  PIN gfpga_pad_GPIO_PAD_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 625.640 2810.000 626.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[21]
  PIN gfpga_pad_GPIO_PAD_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2893.440 4.000 2894.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[22]
  PIN gfpga_pad_GPIO_PAD_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[23]
  PIN gfpga_pad_GPIO_PAD_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1502.840 2810.000 1503.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[24]
  PIN gfpga_pad_GPIO_PAD_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2818.640 2810.000 2819.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[25]
  PIN gfpga_pad_GPIO_PAD_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[26]
  PIN gfpga_pad_GPIO_PAD_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 448.840 2810.000 449.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[27]
  PIN gfpga_pad_GPIO_PAD_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[28]
  PIN gfpga_pad_GPIO_PAD_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.590 0.000 2656.870 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[29]
  PIN gfpga_pad_GPIO_PAD_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 2946.000 1191.770 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[2]
  PIN gfpga_pad_GPIO_PAD_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.490 0.000 2157.770 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[30]
  PIN gfpga_pad_GPIO_PAD_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[31]
  PIN gfpga_pad_GPIO_PAD_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[32]
  PIN gfpga_pad_GPIO_PAD_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 275.440 2810.000 276.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[33]
  PIN gfpga_pad_GPIO_PAD_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2114.840 2810.000 2115.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[34]
  PIN gfpga_pad_GPIO_PAD_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[35]
  PIN gfpga_pad_GPIO_PAD_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.930 0.000 2325.210 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[36]
  PIN gfpga_pad_GPIO_PAD_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1839.440 4.000 1840.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[37]
  PIN gfpga_pad_GPIO_PAD_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 714.040 2810.000 714.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[38]
  PIN gfpga_pad_GPIO_PAD_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 4.000 2455.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[39]
  PIN gfpga_pad_GPIO_PAD_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1679.640 2810.000 1680.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[3]
  PIN gfpga_pad_GPIO_PAD_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2468.440 2810.000 2469.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[40]
  PIN gfpga_pad_GPIO_PAD_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2572.870 0.000 2573.150 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[41]
  PIN gfpga_pad_GPIO_PAD_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 2641.840 2810.000 2642.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[42]
  PIN gfpga_pad_GPIO_PAD_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[43]
  PIN gfpga_pad_GPIO_PAD_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2628.240 4.000 2628.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[44]
  PIN gfpga_pad_GPIO_PAD_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[45]
  PIN gfpga_pad_GPIO_PAD_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[46]
  PIN gfpga_pad_GPIO_PAD_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[47]
  PIN gfpga_pad_GPIO_PAD_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2805.040 4.000 2805.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[48]
  PIN gfpga_pad_GPIO_PAD_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 2946.000 776.390 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[49]
  PIN gfpga_pad_GPIO_PAD_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 2946.000 1771.370 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[4]
  PIN gfpga_pad_GPIO_PAD_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2278.040 4.000 2278.640 ;
    END
  END gfpga_pad_GPIO_PAD_out[50]
  PIN gfpga_pad_GPIO_PAD_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[51]
  PIN gfpga_pad_GPIO_PAD_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[52]
  PIN gfpga_pad_GPIO_PAD_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 2946.000 2186.750 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[53]
  PIN gfpga_pad_GPIO_PAD_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 2946.000 1607.150 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[54]
  PIN gfpga_pad_GPIO_PAD_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[55]
  PIN gfpga_pad_GPIO_PAD_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.130 2946.000 2518.410 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[56]
  PIN gfpga_pad_GPIO_PAD_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 537.240 2810.000 537.840 ;
    END
  END gfpga_pad_GPIO_PAD_out[57]
  PIN gfpga_pad_GPIO_PAD_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2716.640 4.000 2717.240 ;
    END
  END gfpga_pad_GPIO_PAD_out[58]
  PIN gfpga_pad_GPIO_PAD_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[59]
  PIN gfpga_pad_GPIO_PAD_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[5]
  PIN gfpga_pad_GPIO_PAD_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[60]
  PIN gfpga_pad_GPIO_PAD_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END gfpga_pad_GPIO_PAD_out[61]
  PIN gfpga_pad_GPIO_PAD_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1941.440 2810.000 1942.040 ;
    END
  END gfpga_pad_GPIO_PAD_out[62]
  PIN gfpga_pad_GPIO_PAD_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 0.000 1578.170 4.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[63]
  PIN gfpga_pad_GPIO_PAD_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 2946.000 2103.030 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[6]
  PIN gfpga_pad_GPIO_PAD_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 2946.000 2019.310 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[7]
  PIN gfpga_pad_GPIO_PAD_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 2946.000 26.130 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[8]
  PIN gfpga_pad_GPIO_PAD_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 2946.000 525.230 2950.000 ;
    END
  END gfpga_pad_GPIO_PAD_out[9]
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.270 0.000 1993.550 4.000 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END prog_clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2539.840 4.000 2540.440 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2806.000 1414.440 2810.000 1415.040 ;
    END
  END set
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 41.720 10.640 43.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.720 10.640 113.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.720 10.640 183.320 157.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.720 348.725 183.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.720 10.640 253.320 155.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.720 353.220 253.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 10.640 323.320 555.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 747.125 323.320 810.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 893.765 323.320 1065.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 1257.125 323.320 1320.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 1403.765 323.320 1575.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 1767.125 323.320 1830.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 1913.765 323.320 2103.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 2249.925 323.320 2340.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.720 2423.765 323.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.720 10.640 393.320 555.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.720 747.125 393.320 1065.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.720 1257.125 393.320 1575.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.720 1767.125 393.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.720 10.640 463.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.720 10.640 533.320 800.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.720 1017.260 533.320 1310.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.720 1527.260 533.320 1820.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.720 2037.260 533.320 2330.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.720 2547.260 533.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 10.640 603.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 387.365 603.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 990.325 603.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 1500.325 603.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 2010.325 603.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 2270.325 603.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.720 2520.325 603.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 10.640 673.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 387.365 673.320 584.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 607.725 673.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 990.325 673.320 1094.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 1117.725 673.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 1500.325 673.320 1604.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 1627.725 673.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2010.325 673.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2270.325 673.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.720 2520.325 673.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.720 10.640 743.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 10.640 813.320 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 471.685 813.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 736.725 813.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 1246.725 813.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 1756.725 813.320 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 811.720 2287.125 813.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 10.640 883.320 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 471.685 883.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 736.725 883.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 1246.725 883.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 1756.725 883.320 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 881.720 2287.125 883.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.720 10.640 953.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.720 736.725 953.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.720 1246.725 953.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.720 1756.725 953.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 10.640 1023.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 990.325 1023.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 1500.325 1023.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 2010.325 1023.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.720 2520.325 1023.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 10.640 1093.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 990.325 1093.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 1500.325 1093.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2010.325 1093.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2270.325 1093.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1091.720 2520.325 1093.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 10.640 1163.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 387.365 1163.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 990.325 1163.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 1500.325 1163.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 2010.325 1163.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 2270.325 1163.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.720 2520.325 1163.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1231.720 10.640 1233.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 10.640 1303.320 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 471.685 1303.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 736.725 1303.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 1246.725 1303.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 1756.725 1303.320 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.720 2287.125 1303.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 10.640 1373.320 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 471.685 1373.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 736.725 1373.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 1246.725 1373.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 1756.725 1373.320 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.720 2287.125 1373.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 10.640 1443.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 736.725 1443.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 1246.725 1443.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1441.720 1756.725 1443.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1511.720 10.640 1513.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.720 10.640 1583.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.720 990.325 1583.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.720 1500.325 1583.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.720 2010.325 1583.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1581.720 2520.325 1583.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 10.640 1653.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 387.365 1653.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 990.325 1653.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 1500.325 1653.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 2010.325 1653.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 2270.325 1653.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.720 2520.325 1653.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 10.640 1723.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 387.365 1723.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 990.325 1723.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 1500.325 1723.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 2010.325 1723.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.720 2520.325 1723.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1791.720 10.640 1793.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 10.640 1863.320 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 471.685 1863.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 736.725 1863.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1246.725 1863.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 1756.725 1863.320 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1861.720 2287.125 1863.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.720 10.640 1933.320 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.720 736.725 1933.320 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.720 1246.725 1933.320 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.720 1756.725 1933.320 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1931.720 2287.125 1933.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2001.720 10.640 2003.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.720 10.640 2073.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.720 990.325 2073.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.720 1500.325 2073.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.720 2010.325 2073.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.720 2520.325 2073.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 10.640 2143.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 387.365 2143.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 990.325 2143.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 1500.325 2143.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 2010.325 2143.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 2270.325 2143.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2141.720 2520.325 2143.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 10.640 2213.320 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 387.365 2213.320 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 990.325 2213.320 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 1500.325 2213.320 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 2010.325 2213.320 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 2270.325 2213.320 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2211.720 2520.325 2213.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.720 10.640 2283.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 10.640 2353.320 289.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 473.045 2353.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 704.405 2353.320 777.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 863.525 2353.320 1022.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 1214.405 2353.320 1287.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 1373.525 2353.320 1532.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 1724.405 2353.320 1797.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 1883.525 2353.320 2307.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.720 2393.525 2353.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.720 10.640 2423.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.720 704.405 2423.320 1022.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.720 1214.405 2423.320 1532.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.720 1724.405 2423.320 2047.555 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.720 2171.845 2423.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2491.720 10.640 2493.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2561.720 10.640 2563.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2631.720 10.640 2633.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2701.720 10.640 2703.320 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2771.720 10.640 2773.320 2937.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 47.080 2804.400 48.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 122.080 2804.400 123.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 197.080 2804.400 198.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 272.080 2804.400 273.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 347.080 2804.400 348.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 422.080 2804.400 423.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 497.080 2804.400 498.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 572.080 2804.400 573.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 647.080 2804.400 648.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 722.080 2804.400 723.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 797.080 2804.400 798.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 872.080 2804.400 873.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 947.080 517.380 948.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1022.080 2804.400 1023.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1097.080 2804.400 1098.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1172.080 2804.400 1173.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1247.080 2804.400 1248.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1322.080 2804.400 1323.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1397.080 517.380 1398.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1472.080 517.380 1473.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1547.080 2357.380 1548.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1622.080 2804.400 1623.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1697.080 2804.400 1698.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1772.080 2804.400 1773.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1847.080 2804.400 1848.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1922.080 517.380 1923.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1997.080 2804.400 1998.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2072.080 2804.400 2073.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2147.080 2804.400 2148.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2222.080 2804.400 2223.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2297.080 2804.400 2298.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2372.080 2804.400 2373.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2447.080 517.380 2448.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2522.080 2804.400 2523.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2597.080 2804.400 2598.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2672.080 2804.400 2673.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2747.080 2804.400 2748.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2822.080 2804.400 2823.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2897.080 2804.400 2898.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 947.080 1027.380 948.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 1397.080 1027.380 1398.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 1472.080 1027.380 1473.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 1922.080 1027.380 1923.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 2447.080 1027.380 2448.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 947.080 1537.380 948.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 1397.080 1537.380 1398.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 1472.080 1537.380 1473.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 1922.080 1537.380 1923.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 2447.080 1537.380 2448.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 947.080 2047.380 948.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 1397.080 2047.380 1398.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 1472.080 2047.380 1473.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 1922.080 2047.380 1923.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 2447.080 2047.380 2448.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 947.080 2804.400 948.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 1397.080 2804.400 1398.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 1472.080 2804.400 1473.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 1922.080 2804.400 1923.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 2447.080 2804.400 2448.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 2487.060 1547.080 2804.400 1548.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.540 524.720 14.140 753.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 512.100 1046.960 513.700 1273.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.380 1569.200 1257.980 1781.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.140 2075.120 1766.740 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 785.840 2018.820 805.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.420 1275.440 2534.020 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2790.020 1786.800 2791.620 2013.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.540 1036.080 14.140 1265.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.740 535.600 506.340 764.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.860 785.840 999.460 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.540 269.040 1256.140 492.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.140 1566.480 1766.740 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 1294.480 2018.820 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.420 1786.800 2534.020 1999.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2790.020 2295.440 2791.620 2524.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.540 1544.720 14.140 1773.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.740 2066.960 506.340 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.540 1055.120 1256.140 1270.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.140 266.320 1766.740 495.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 805.660 2018.820 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.420 2295.440 2534.020 2508.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2790.020 1275.440 2791.620 1504.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.540 2056.080 14.140 2285.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.740 1555.600 506.340 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.540 546.480 1256.140 764.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.500 785.840 1774.100 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.580 266.320 2026.180 495.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.860 1294.480 999.460 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.540 2075.120 1256.140 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.140 546.480 1766.740 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.580 1055.120 2026.180 1278.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.820 785.840 1264.420 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.140 1055.120 1766.740 1273.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.580 546.480 2026.180 764.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.860 1805.840 999.460 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.820 1294.480 1264.420 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.500 2314.480 1774.100 2543.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.580 1566.480 2026.180 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2532.420 766.800 2534.020 979.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.820 1805.840 1264.420 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.500 1294.480 1774.100 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 2314.480 2018.820 2334.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2790.020 766.800 2791.620 993.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 997.860 2314.480 999.460 2543.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.500 1805.840 1774.100 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 1314.300 2018.820 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.820 2314.480 1264.420 2543.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 1805.840 2018.820 1825.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.720 1286.100 396.620 1287.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 1825.660 2018.820 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2024.580 2075.120 2026.180 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.220 2334.300 2018.820 2543.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 45.020 10.640 46.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.020 10.640 116.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.020 10.640 186.620 157.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.020 348.725 186.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 255.020 10.640 256.620 157.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 255.020 348.725 256.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 10.640 326.620 555.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 747.125 326.620 810.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 893.765 326.620 1065.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 1257.125 326.620 1320.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 1403.765 326.620 1575.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 1767.125 326.620 1830.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 1913.765 326.620 2103.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 2249.925 326.620 2340.275 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.020 2423.765 326.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 395.020 10.640 396.620 555.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 395.020 747.125 396.620 1065.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 395.020 1257.125 396.620 1575.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 395.020 1767.125 396.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 10.640 466.620 550.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 748.220 466.620 1060.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 1258.220 466.620 1570.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 1768.220 466.620 2080.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.020 2278.220 466.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.020 10.640 536.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.020 990.325 536.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.020 1500.325 536.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.020 2010.325 536.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.020 2520.325 536.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 10.640 606.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 387.365 606.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 990.325 606.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 1500.325 606.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 2010.325 606.620 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 2270.325 606.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 605.020 2520.325 606.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 10.640 676.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 387.365 676.620 584.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 607.725 676.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 990.325 676.620 1094.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 1117.725 676.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 1500.325 676.620 1604.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 1627.725 676.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2010.325 676.620 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2270.325 676.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.020 2520.325 676.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 745.020 10.640 746.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 10.640 816.620 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 471.685 816.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 736.725 816.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 1246.725 816.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 1756.725 816.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 815.020 2287.125 816.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 10.640 886.620 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 471.685 886.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 736.725 886.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 1246.725 886.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 1756.725 886.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 885.020 2287.125 886.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 10.640 956.620 280.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 478.220 956.620 560.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 758.220 956.620 800.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 998.220 956.620 1070.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 1268.220 956.620 1310.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 1508.220 956.620 1580.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 1778.220 956.620 1820.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 2018.220 956.620 2090.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 2288.220 956.620 2330.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.020 2528.220 956.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 10.640 1026.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 990.325 1026.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 1500.325 1026.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 2010.325 1026.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.020 2520.325 1026.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 10.640 1096.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 990.325 1096.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 1500.325 1096.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2010.325 1096.620 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2270.325 1096.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.020 2520.325 1096.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 10.640 1166.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 387.365 1166.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 990.325 1166.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 1500.325 1166.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 2010.325 1166.620 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 2270.325 1166.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1165.020 2520.325 1166.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1235.020 10.640 1236.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 10.640 1306.620 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 471.685 1306.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 736.725 1306.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 1246.725 1306.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 1756.725 1306.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.020 2287.125 1306.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 10.640 1376.620 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 471.685 1376.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 736.725 1376.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 1246.725 1376.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 1756.725 1376.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.020 2287.125 1376.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 10.640 1446.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 736.725 1446.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 1246.725 1446.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.020 1756.725 1446.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1515.020 10.640 1516.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 10.640 1586.620 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 228.220 1586.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 990.325 1586.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 1500.325 1586.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 2010.325 1586.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 2520.325 1586.620 2610.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1585.020 2808.220 1586.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 10.640 1656.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 387.365 1656.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 990.325 1656.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 1500.325 1656.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2010.325 1656.620 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2270.325 1656.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1655.020 2520.325 1656.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 10.640 1726.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 387.365 1726.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 990.325 1726.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 1500.325 1726.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 2010.325 1726.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.020 2520.325 1726.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1795.020 10.640 1796.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1795.020 2287.125 1796.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 10.640 1866.620 317.475 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 471.685 1866.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 736.725 1866.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 1246.725 1866.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 1756.725 1866.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1865.020 2287.125 1866.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.020 10.640 1936.620 562.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.020 736.725 1936.620 1072.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.020 1246.725 1936.620 1582.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.020 1756.725 1936.620 2092.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.020 2287.125 1936.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2005.020 10.640 2006.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 10.640 2076.620 280.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 478.220 2076.620 550.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 748.220 2076.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 990.325 2076.620 1063.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 1261.220 2076.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 1500.325 2076.620 1570.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 1768.220 2076.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 2010.325 2076.620 2080.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 2278.220 2076.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.020 2520.325 2076.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 10.640 2146.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 387.365 2146.620 801.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 990.325 2146.620 1311.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 1500.325 2146.620 1821.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 2010.325 2146.620 2085.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 2270.325 2146.620 2331.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.020 2520.325 2146.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.020 10.640 2216.620 282.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.020 387.365 2216.620 800.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.020 1017.260 2216.620 1310.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.020 1527.260 2216.620 1820.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.020 2037.260 2216.620 2330.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2215.020 2547.260 2216.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.020 10.640 2286.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 10.640 2356.620 289.595 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 473.045 2356.620 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 704.405 2356.620 777.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 863.525 2356.620 1022.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 1214.405 2356.620 1287.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 1373.525 2356.620 1532.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 1724.405 2356.620 1797.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 1883.525 2356.620 2307.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 2355.020 2393.525 2356.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.020 10.640 2426.620 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.020 704.405 2426.620 1022.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.020 1214.405 2426.620 1532.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.020 1724.405 2426.620 2040.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.020 2189.260 2426.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2495.020 10.640 2496.620 2040.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2495.020 2189.260 2496.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2565.020 10.640 2566.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2635.020 10.640 2636.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2705.020 10.640 2706.620 2937.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2775.020 10.640 2776.620 2937.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 50.380 2804.400 51.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 125.380 2804.400 126.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 200.380 2804.400 201.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 275.380 2804.400 276.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 350.380 2804.400 351.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 425.380 2804.400 426.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 500.380 2804.400 501.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 575.380 2804.400 576.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 650.380 2804.400 651.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 725.380 2804.400 726.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 800.380 2804.400 801.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 875.380 2804.400 876.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 950.380 517.380 951.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1025.380 2357.380 1026.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1100.380 2804.400 1101.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1175.380 2804.400 1176.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1250.380 2804.400 1251.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1325.380 2804.400 1326.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1400.380 517.380 1401.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1475.380 517.380 1476.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1550.380 2357.380 1551.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1625.380 2804.400 1626.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1700.380 2804.400 1701.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1775.380 2804.400 1776.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1850.380 2804.400 1851.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1925.380 517.380 1926.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2000.380 2804.400 2001.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2075.380 2804.400 2076.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2150.380 2804.400 2151.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2225.380 2804.400 2226.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2300.380 2804.400 2301.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2375.380 2804.400 2376.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2450.380 517.380 2451.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2525.380 2804.400 2526.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2600.380 2804.400 2601.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2675.380 2804.400 2676.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2750.380 2804.400 2751.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2825.380 2804.400 2826.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2900.380 2804.400 2901.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 950.380 1027.380 951.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 1400.380 1027.380 1401.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 1475.380 1027.380 1476.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 1925.380 1027.380 1926.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 633.260 2450.380 1027.380 2451.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 950.380 1537.380 951.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 1400.380 1537.380 1401.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 1475.380 1537.380 1476.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 1925.380 1537.380 1926.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1143.260 2450.380 1537.380 2451.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 950.380 2047.380 951.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 1400.380 2047.380 1401.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 1475.380 2047.380 1476.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 1925.380 2047.380 1926.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 1653.260 2450.380 2047.380 2451.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 950.380 2804.400 951.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 1400.380 2804.400 1401.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 1475.380 2804.400 1476.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 1925.380 2804.400 1926.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2163.260 2450.380 2804.400 2451.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2487.060 1025.380 2804.400 1026.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 2487.060 1550.380 2804.400 1551.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.220 524.720 17.820 753.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 515.780 1046.960 517.380 1273.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.060 266.320 1008.660 495.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.820 2075.120 1770.420 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 785.840 2022.500 805.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.100 1275.440 2537.700 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.700 1786.800 2795.300 2013.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.220 1036.080 17.820 1265.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.420 535.600 510.020 764.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.540 785.840 1003.140 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.220 269.040 1259.820 492.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.820 1566.480 1770.420 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 1294.480 2022.500 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.100 1786.800 2537.700 1999.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.700 2295.440 2795.300 2524.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.220 1544.720 17.820 1773.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.420 2066.960 510.020 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.060 549.200 1008.660 761.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.220 1055.120 1259.820 1270.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.820 266.320 1770.420 495.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 805.660 2022.500 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.100 2295.440 2537.700 2508.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.700 1275.440 2795.300 1504.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.220 2056.080 17.820 2285.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.420 1555.600 510.020 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.060 1055.120 1008.660 1273.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.220 546.480 1259.820 764.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.180 785.840 1777.780 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.260 266.320 2029.860 495.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.540 1294.480 1003.140 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.220 2075.120 1259.820 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.820 546.480 1770.420 775.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.260 1055.120 2029.860 1278.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.060 1566.480 1008.660 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.500 785.840 1268.100 1014.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.820 1055.120 1770.420 1273.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.260 546.480 2029.860 764.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.540 1805.840 1003.140 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.500 1294.480 1268.100 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.180 2314.480 1777.780 2543.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.260 1566.480 2029.860 1784.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2536.100 766.800 2537.700 979.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1007.060 2077.840 1008.660 2290.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.500 1805.840 1268.100 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.180 1294.480 1777.780 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 2314.480 2022.500 2334.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2793.700 766.800 2795.300 993.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.540 2314.480 1003.140 2543.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.180 1805.840 1777.780 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 1314.300 2022.500 1523.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1266.500 2314.480 1268.100 2543.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 1805.840 2022.500 1825.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 251.720 1289.500 396.620 1291.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 1825.660 2022.500 2034.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2028.260 2075.120 2029.860 2293.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.900 2334.300 2022.500 2543.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2804.160 2937.685 ;
      LAYER met1 ;
        RECT 0.070 8.880 2804.160 2937.840 ;
      LAYER met2 ;
        RECT 0.100 2945.720 25.570 2946.170 ;
        RECT 26.410 2945.720 109.290 2946.170 ;
        RECT 110.130 2945.720 193.010 2946.170 ;
        RECT 193.850 2945.720 276.730 2946.170 ;
        RECT 277.570 2945.720 360.450 2946.170 ;
        RECT 361.290 2945.720 440.950 2946.170 ;
        RECT 441.790 2945.720 524.670 2946.170 ;
        RECT 525.510 2945.720 608.390 2946.170 ;
        RECT 609.230 2945.720 692.110 2946.170 ;
        RECT 692.950 2945.720 775.830 2946.170 ;
        RECT 776.670 2945.720 856.330 2946.170 ;
        RECT 857.170 2945.720 940.050 2946.170 ;
        RECT 940.890 2945.720 1023.770 2946.170 ;
        RECT 1024.610 2945.720 1107.490 2946.170 ;
        RECT 1108.330 2945.720 1191.210 2946.170 ;
        RECT 1192.050 2945.720 1271.710 2946.170 ;
        RECT 1272.550 2945.720 1355.430 2946.170 ;
        RECT 1356.270 2945.720 1439.150 2946.170 ;
        RECT 1439.990 2945.720 1522.870 2946.170 ;
        RECT 1523.710 2945.720 1606.590 2946.170 ;
        RECT 1607.430 2945.720 1687.090 2946.170 ;
        RECT 1687.930 2945.720 1770.810 2946.170 ;
        RECT 1771.650 2945.720 1854.530 2946.170 ;
        RECT 1855.370 2945.720 1938.250 2946.170 ;
        RECT 1939.090 2945.720 2018.750 2946.170 ;
        RECT 2019.590 2945.720 2102.470 2946.170 ;
        RECT 2103.310 2945.720 2186.190 2946.170 ;
        RECT 2187.030 2945.720 2269.910 2946.170 ;
        RECT 2270.750 2945.720 2353.630 2946.170 ;
        RECT 2354.470 2945.720 2434.130 2946.170 ;
        RECT 2434.970 2945.720 2517.850 2946.170 ;
        RECT 2518.690 2945.720 2601.570 2946.170 ;
        RECT 2602.410 2945.720 2685.290 2946.170 ;
        RECT 2686.130 2945.720 2769.010 2946.170 ;
        RECT 2769.850 2945.720 2802.220 2946.170 ;
        RECT 0.100 4.280 2802.220 2945.720 ;
        RECT 0.650 3.670 80.310 4.280 ;
        RECT 81.150 3.670 164.030 4.280 ;
        RECT 164.870 3.670 247.750 4.280 ;
        RECT 248.590 3.670 331.470 4.280 ;
        RECT 332.310 3.670 411.970 4.280 ;
        RECT 412.810 3.670 495.690 4.280 ;
        RECT 496.530 3.670 579.410 4.280 ;
        RECT 580.250 3.670 663.130 4.280 ;
        RECT 663.970 3.670 746.850 4.280 ;
        RECT 747.690 3.670 827.350 4.280 ;
        RECT 828.190 3.670 911.070 4.280 ;
        RECT 911.910 3.670 994.790 4.280 ;
        RECT 995.630 3.670 1078.510 4.280 ;
        RECT 1079.350 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1242.730 4.280 ;
        RECT 1243.570 3.670 1326.450 4.280 ;
        RECT 1327.290 3.670 1410.170 4.280 ;
        RECT 1411.010 3.670 1493.890 4.280 ;
        RECT 1494.730 3.670 1577.610 4.280 ;
        RECT 1578.450 3.670 1658.110 4.280 ;
        RECT 1658.950 3.670 1741.830 4.280 ;
        RECT 1742.670 3.670 1825.550 4.280 ;
        RECT 1826.390 3.670 1909.270 4.280 ;
        RECT 1910.110 3.670 1992.990 4.280 ;
        RECT 1993.830 3.670 2073.490 4.280 ;
        RECT 2074.330 3.670 2157.210 4.280 ;
        RECT 2158.050 3.670 2240.930 4.280 ;
        RECT 2241.770 3.670 2324.650 4.280 ;
        RECT 2325.490 3.670 2405.150 4.280 ;
        RECT 2405.990 3.670 2488.870 4.280 ;
        RECT 2489.710 3.670 2572.590 4.280 ;
        RECT 2573.430 3.670 2656.310 4.280 ;
        RECT 2657.150 3.670 2740.030 4.280 ;
        RECT 2740.870 3.670 2802.220 4.280 ;
      LAYER met3 ;
        RECT 4.000 2908.040 2806.000 2937.765 ;
        RECT 4.000 2906.640 2805.600 2908.040 ;
        RECT 4.000 2894.440 2806.000 2906.640 ;
        RECT 4.400 2893.040 2806.000 2894.440 ;
        RECT 4.000 2819.640 2806.000 2893.040 ;
        RECT 4.000 2818.240 2805.600 2819.640 ;
        RECT 4.000 2806.040 2806.000 2818.240 ;
        RECT 4.400 2804.640 2806.000 2806.040 ;
        RECT 4.000 2731.240 2806.000 2804.640 ;
        RECT 4.000 2729.840 2805.600 2731.240 ;
        RECT 4.000 2717.640 2806.000 2729.840 ;
        RECT 4.400 2716.240 2806.000 2717.640 ;
        RECT 4.000 2642.840 2806.000 2716.240 ;
        RECT 4.000 2641.440 2805.600 2642.840 ;
        RECT 4.000 2629.240 2806.000 2641.440 ;
        RECT 4.400 2627.840 2806.000 2629.240 ;
        RECT 4.000 2554.440 2806.000 2627.840 ;
        RECT 4.000 2553.040 2805.600 2554.440 ;
        RECT 4.000 2540.840 2806.000 2553.040 ;
        RECT 4.400 2539.440 2806.000 2540.840 ;
        RECT 4.000 2469.440 2806.000 2539.440 ;
        RECT 4.000 2468.040 2805.600 2469.440 ;
        RECT 4.000 2455.840 2806.000 2468.040 ;
        RECT 4.400 2454.440 2806.000 2455.840 ;
        RECT 4.000 2381.040 2806.000 2454.440 ;
        RECT 4.000 2379.640 2805.600 2381.040 ;
        RECT 4.000 2367.440 2806.000 2379.640 ;
        RECT 4.400 2366.040 2806.000 2367.440 ;
        RECT 4.000 2292.640 2806.000 2366.040 ;
        RECT 4.000 2291.240 2805.600 2292.640 ;
        RECT 4.000 2279.040 2806.000 2291.240 ;
        RECT 4.400 2277.640 2806.000 2279.040 ;
        RECT 4.000 2204.240 2806.000 2277.640 ;
        RECT 4.000 2202.840 2805.600 2204.240 ;
        RECT 4.000 2190.640 2806.000 2202.840 ;
        RECT 4.400 2189.240 2806.000 2190.640 ;
        RECT 4.000 2115.840 2806.000 2189.240 ;
        RECT 4.000 2114.440 2805.600 2115.840 ;
        RECT 4.000 2105.640 2806.000 2114.440 ;
        RECT 4.400 2104.240 2806.000 2105.640 ;
        RECT 4.000 2030.840 2806.000 2104.240 ;
        RECT 4.000 2029.440 2805.600 2030.840 ;
        RECT 4.000 2017.240 2806.000 2029.440 ;
        RECT 4.400 2015.840 2806.000 2017.240 ;
        RECT 4.000 1942.440 2806.000 2015.840 ;
        RECT 4.000 1941.040 2805.600 1942.440 ;
        RECT 4.000 1928.840 2806.000 1941.040 ;
        RECT 4.400 1927.440 2806.000 1928.840 ;
        RECT 4.000 1854.040 2806.000 1927.440 ;
        RECT 4.000 1852.640 2805.600 1854.040 ;
        RECT 4.000 1840.440 2806.000 1852.640 ;
        RECT 4.400 1839.040 2806.000 1840.440 ;
        RECT 4.000 1765.640 2806.000 1839.040 ;
        RECT 4.000 1764.240 2805.600 1765.640 ;
        RECT 4.000 1752.040 2806.000 1764.240 ;
        RECT 4.400 1750.640 2806.000 1752.040 ;
        RECT 4.000 1680.640 2806.000 1750.640 ;
        RECT 4.000 1679.240 2805.600 1680.640 ;
        RECT 4.000 1667.040 2806.000 1679.240 ;
        RECT 4.400 1665.640 2806.000 1667.040 ;
        RECT 4.000 1592.240 2806.000 1665.640 ;
        RECT 4.000 1590.840 2805.600 1592.240 ;
        RECT 4.000 1578.640 2806.000 1590.840 ;
        RECT 4.400 1577.240 2806.000 1578.640 ;
        RECT 4.000 1503.840 2806.000 1577.240 ;
        RECT 4.000 1502.440 2805.600 1503.840 ;
        RECT 4.000 1490.240 2806.000 1502.440 ;
        RECT 4.400 1488.840 2806.000 1490.240 ;
        RECT 4.000 1415.440 2806.000 1488.840 ;
        RECT 4.000 1414.040 2805.600 1415.440 ;
        RECT 4.000 1401.840 2806.000 1414.040 ;
        RECT 4.400 1400.440 2806.000 1401.840 ;
        RECT 4.000 1327.040 2806.000 1400.440 ;
        RECT 4.000 1325.640 2805.600 1327.040 ;
        RECT 4.000 1313.440 2806.000 1325.640 ;
        RECT 4.400 1312.040 2806.000 1313.440 ;
        RECT 4.000 1242.040 2806.000 1312.040 ;
        RECT 4.000 1240.640 2805.600 1242.040 ;
        RECT 4.000 1228.440 2806.000 1240.640 ;
        RECT 4.400 1227.040 2806.000 1228.440 ;
        RECT 4.000 1153.640 2806.000 1227.040 ;
        RECT 4.000 1152.240 2805.600 1153.640 ;
        RECT 4.000 1140.040 2806.000 1152.240 ;
        RECT 4.400 1138.640 2806.000 1140.040 ;
        RECT 4.000 1065.240 2806.000 1138.640 ;
        RECT 4.000 1063.840 2805.600 1065.240 ;
        RECT 4.000 1051.640 2806.000 1063.840 ;
        RECT 4.400 1050.240 2806.000 1051.640 ;
        RECT 4.000 976.840 2806.000 1050.240 ;
        RECT 4.000 975.440 2805.600 976.840 ;
        RECT 4.000 963.240 2806.000 975.440 ;
        RECT 4.400 961.840 2806.000 963.240 ;
        RECT 4.000 888.440 2806.000 961.840 ;
        RECT 4.000 887.040 2805.600 888.440 ;
        RECT 4.000 874.840 2806.000 887.040 ;
        RECT 4.400 873.440 2806.000 874.840 ;
        RECT 4.000 803.440 2806.000 873.440 ;
        RECT 4.000 802.040 2805.600 803.440 ;
        RECT 4.000 789.840 2806.000 802.040 ;
        RECT 4.400 788.440 2806.000 789.840 ;
        RECT 4.000 715.040 2806.000 788.440 ;
        RECT 4.000 713.640 2805.600 715.040 ;
        RECT 4.000 701.440 2806.000 713.640 ;
        RECT 4.400 700.040 2806.000 701.440 ;
        RECT 4.000 626.640 2806.000 700.040 ;
        RECT 4.000 625.240 2805.600 626.640 ;
        RECT 4.000 613.040 2806.000 625.240 ;
        RECT 4.400 611.640 2806.000 613.040 ;
        RECT 4.000 538.240 2806.000 611.640 ;
        RECT 4.000 536.840 2805.600 538.240 ;
        RECT 4.000 524.640 2806.000 536.840 ;
        RECT 4.400 523.240 2806.000 524.640 ;
        RECT 4.000 449.840 2806.000 523.240 ;
        RECT 4.000 448.440 2805.600 449.840 ;
        RECT 4.000 436.240 2806.000 448.440 ;
        RECT 4.400 434.840 2806.000 436.240 ;
        RECT 4.000 364.840 2806.000 434.840 ;
        RECT 4.000 363.440 2805.600 364.840 ;
        RECT 4.000 351.240 2806.000 363.440 ;
        RECT 4.400 349.840 2806.000 351.240 ;
        RECT 4.000 276.440 2806.000 349.840 ;
        RECT 4.000 275.040 2805.600 276.440 ;
        RECT 4.000 262.840 2806.000 275.040 ;
        RECT 4.400 261.440 2806.000 262.840 ;
        RECT 4.000 188.040 2806.000 261.440 ;
        RECT 4.000 186.640 2805.600 188.040 ;
        RECT 4.000 174.440 2806.000 186.640 ;
        RECT 4.400 173.040 2806.000 174.440 ;
        RECT 4.000 99.640 2806.000 173.040 ;
        RECT 4.000 98.240 2805.600 99.640 ;
        RECT 4.000 86.040 2806.000 98.240 ;
        RECT 4.400 84.640 2806.000 86.040 ;
        RECT 4.000 11.240 2806.000 84.640 ;
        RECT 4.000 10.375 2805.600 11.240 ;
      LAYER met4 ;
        RECT 35.750 11.735 41.320 2936.745 ;
        RECT 43.720 11.735 44.620 2936.745 ;
        RECT 47.020 11.735 111.320 2936.745 ;
        RECT 113.720 11.735 114.620 2936.745 ;
        RECT 117.020 348.325 181.320 2936.745 ;
        RECT 183.720 348.325 184.620 2936.745 ;
        RECT 187.020 352.820 251.320 2936.745 ;
        RECT 253.720 352.820 254.620 2936.745 ;
        RECT 187.020 348.325 254.620 352.820 ;
        RECT 257.020 2423.365 321.320 2936.745 ;
        RECT 323.720 2423.365 324.620 2936.745 ;
        RECT 327.020 2423.365 391.320 2936.745 ;
        RECT 257.020 2340.675 391.320 2423.365 ;
        RECT 257.020 2249.525 321.320 2340.675 ;
        RECT 323.720 2249.525 324.620 2340.675 ;
        RECT 327.020 2249.525 391.320 2340.675 ;
        RECT 257.020 2104.275 391.320 2249.525 ;
        RECT 257.020 1913.365 321.320 2104.275 ;
        RECT 323.720 1913.365 324.620 2104.275 ;
        RECT 327.020 1913.365 391.320 2104.275 ;
        RECT 257.020 1830.675 391.320 1913.365 ;
        RECT 257.020 1766.725 321.320 1830.675 ;
        RECT 323.720 1766.725 324.620 1830.675 ;
        RECT 327.020 1766.725 391.320 1830.675 ;
        RECT 393.720 1766.725 394.620 2936.745 ;
        RECT 397.020 1766.725 461.320 2936.745 ;
        RECT 257.020 1575.915 461.320 1766.725 ;
        RECT 257.020 1403.365 321.320 1575.915 ;
        RECT 323.720 1403.365 324.620 1575.915 ;
        RECT 327.020 1403.365 391.320 1575.915 ;
        RECT 257.020 1320.675 391.320 1403.365 ;
        RECT 257.020 1256.725 321.320 1320.675 ;
        RECT 323.720 1256.725 324.620 1320.675 ;
        RECT 327.020 1256.725 391.320 1320.675 ;
        RECT 393.720 1256.725 394.620 1575.915 ;
        RECT 397.020 1256.725 461.320 1575.915 ;
        RECT 257.020 1065.915 461.320 1256.725 ;
        RECT 257.020 893.365 321.320 1065.915 ;
        RECT 323.720 893.365 324.620 1065.915 ;
        RECT 327.020 893.365 391.320 1065.915 ;
        RECT 257.020 810.675 391.320 893.365 ;
        RECT 257.020 746.725 321.320 810.675 ;
        RECT 323.720 746.725 324.620 810.675 ;
        RECT 327.020 746.725 391.320 810.675 ;
        RECT 393.720 746.725 394.620 1065.915 ;
        RECT 397.020 746.725 461.320 1065.915 ;
        RECT 257.020 555.915 461.320 746.725 ;
        RECT 257.020 348.325 321.320 555.915 ;
        RECT 117.020 158.195 321.320 348.325 ;
        RECT 117.020 11.735 181.320 158.195 ;
        RECT 183.720 11.735 184.620 158.195 ;
        RECT 187.020 155.740 254.620 158.195 ;
        RECT 187.020 11.735 251.320 155.740 ;
        RECT 253.720 11.735 254.620 155.740 ;
        RECT 257.020 11.735 321.320 158.195 ;
        RECT 323.720 11.735 324.620 555.915 ;
        RECT 327.020 11.735 391.320 555.915 ;
        RECT 393.720 11.735 394.620 555.915 ;
        RECT 397.020 11.735 461.320 555.915 ;
        RECT 463.720 2277.820 464.620 2936.745 ;
        RECT 467.020 2546.860 531.320 2936.745 ;
        RECT 533.720 2546.860 534.620 2936.745 ;
        RECT 467.020 2519.925 534.620 2546.860 ;
        RECT 537.020 2519.925 601.320 2936.745 ;
        RECT 603.720 2519.925 604.620 2936.745 ;
        RECT 607.020 2519.925 671.320 2936.745 ;
        RECT 673.720 2519.925 674.620 2936.745 ;
        RECT 677.020 2519.925 741.320 2936.745 ;
        RECT 467.020 2331.835 741.320 2519.925 ;
        RECT 467.020 2330.740 534.620 2331.835 ;
        RECT 467.020 2293.600 531.320 2330.740 ;
        RECT 467.020 2277.820 504.340 2293.600 ;
        RECT 463.720 2080.740 504.340 2277.820 ;
        RECT 463.720 1767.820 464.620 2080.740 ;
        RECT 467.020 2066.560 504.340 2080.740 ;
        RECT 506.740 2066.560 508.020 2293.600 ;
        RECT 510.420 2066.560 531.320 2293.600 ;
        RECT 467.020 2036.860 531.320 2066.560 ;
        RECT 533.720 2036.860 534.620 2330.740 ;
        RECT 467.020 2009.925 534.620 2036.860 ;
        RECT 537.020 2269.925 601.320 2331.835 ;
        RECT 603.720 2269.925 604.620 2331.835 ;
        RECT 607.020 2269.925 671.320 2331.835 ;
        RECT 673.720 2269.925 674.620 2331.835 ;
        RECT 677.020 2269.925 741.320 2331.835 ;
        RECT 537.020 2085.915 741.320 2269.925 ;
        RECT 537.020 2009.925 601.320 2085.915 ;
        RECT 603.720 2009.925 604.620 2085.915 ;
        RECT 607.020 2009.925 671.320 2085.915 ;
        RECT 673.720 2009.925 674.620 2085.915 ;
        RECT 677.020 2009.925 741.320 2085.915 ;
        RECT 467.020 1821.835 741.320 2009.925 ;
        RECT 467.020 1820.740 534.620 1821.835 ;
        RECT 467.020 1784.960 531.320 1820.740 ;
        RECT 467.020 1767.820 504.340 1784.960 ;
        RECT 463.720 1570.740 504.340 1767.820 ;
        RECT 463.720 1257.820 464.620 1570.740 ;
        RECT 467.020 1555.200 504.340 1570.740 ;
        RECT 506.740 1555.200 508.020 1784.960 ;
        RECT 510.420 1555.200 531.320 1784.960 ;
        RECT 467.020 1526.860 531.320 1555.200 ;
        RECT 533.720 1526.860 534.620 1820.740 ;
        RECT 467.020 1499.925 534.620 1526.860 ;
        RECT 537.020 1499.925 601.320 1821.835 ;
        RECT 603.720 1499.925 604.620 1821.835 ;
        RECT 607.020 1627.325 671.320 1821.835 ;
        RECT 673.720 1627.325 674.620 1821.835 ;
        RECT 677.020 1627.325 741.320 1821.835 ;
        RECT 607.020 1605.155 741.320 1627.325 ;
        RECT 607.020 1499.925 671.320 1605.155 ;
        RECT 673.720 1499.925 674.620 1605.155 ;
        RECT 677.020 1499.925 741.320 1605.155 ;
        RECT 467.020 1311.835 741.320 1499.925 ;
        RECT 467.020 1310.740 534.620 1311.835 ;
        RECT 467.020 1273.600 531.320 1310.740 ;
        RECT 467.020 1257.820 511.700 1273.600 ;
        RECT 463.720 1060.740 511.700 1257.820 ;
        RECT 463.720 747.820 464.620 1060.740 ;
        RECT 467.020 1046.560 511.700 1060.740 ;
        RECT 514.100 1046.560 515.380 1273.600 ;
        RECT 517.780 1046.560 531.320 1273.600 ;
        RECT 467.020 1016.860 531.320 1046.560 ;
        RECT 533.720 1016.860 534.620 1310.740 ;
        RECT 467.020 989.925 534.620 1016.860 ;
        RECT 537.020 989.925 601.320 1311.835 ;
        RECT 603.720 989.925 604.620 1311.835 ;
        RECT 607.020 1117.325 671.320 1311.835 ;
        RECT 673.720 1117.325 674.620 1311.835 ;
        RECT 677.020 1117.325 741.320 1311.835 ;
        RECT 607.020 1095.155 741.320 1117.325 ;
        RECT 607.020 989.925 671.320 1095.155 ;
        RECT 673.720 989.925 674.620 1095.155 ;
        RECT 677.020 989.925 741.320 1095.155 ;
        RECT 467.020 801.835 741.320 989.925 ;
        RECT 467.020 800.740 534.620 801.835 ;
        RECT 467.020 764.960 531.320 800.740 ;
        RECT 467.020 747.820 504.340 764.960 ;
        RECT 463.720 550.740 504.340 747.820 ;
        RECT 463.720 11.735 464.620 550.740 ;
        RECT 467.020 535.200 504.340 550.740 ;
        RECT 506.740 535.200 508.020 764.960 ;
        RECT 510.420 535.200 531.320 764.960 ;
        RECT 467.020 11.735 531.320 535.200 ;
        RECT 533.720 11.735 534.620 800.740 ;
        RECT 537.020 386.965 601.320 801.835 ;
        RECT 603.720 386.965 604.620 801.835 ;
        RECT 607.020 607.325 671.320 801.835 ;
        RECT 673.720 607.325 674.620 801.835 ;
        RECT 677.020 607.325 741.320 801.835 ;
        RECT 607.020 585.155 741.320 607.325 ;
        RECT 607.020 386.965 671.320 585.155 ;
        RECT 673.720 386.965 674.620 585.155 ;
        RECT 677.020 386.965 741.320 585.155 ;
        RECT 537.020 282.515 741.320 386.965 ;
        RECT 537.020 11.735 601.320 282.515 ;
        RECT 603.720 11.735 604.620 282.515 ;
        RECT 607.020 11.735 671.320 282.515 ;
        RECT 673.720 11.735 674.620 282.515 ;
        RECT 677.020 11.735 741.320 282.515 ;
        RECT 743.720 11.735 744.620 2936.745 ;
        RECT 747.020 2286.725 811.320 2936.745 ;
        RECT 813.720 2286.725 814.620 2936.745 ;
        RECT 817.020 2286.725 881.320 2936.745 ;
        RECT 883.720 2286.725 884.620 2936.745 ;
        RECT 887.020 2286.725 951.320 2936.745 ;
        RECT 747.020 2093.195 951.320 2286.725 ;
        RECT 747.020 1756.325 811.320 2093.195 ;
        RECT 813.720 1756.325 814.620 2093.195 ;
        RECT 817.020 1756.325 881.320 2093.195 ;
        RECT 883.720 1756.325 884.620 2093.195 ;
        RECT 887.020 1756.325 951.320 2093.195 ;
        RECT 953.720 2527.820 954.620 2936.745 ;
        RECT 957.020 2543.840 1021.320 2936.745 ;
        RECT 957.020 2527.820 997.460 2543.840 ;
        RECT 953.720 2330.740 997.460 2527.820 ;
        RECT 953.720 2287.820 954.620 2330.740 ;
        RECT 957.020 2314.080 997.460 2330.740 ;
        RECT 999.860 2314.080 1001.140 2543.840 ;
        RECT 1003.540 2519.925 1021.320 2543.840 ;
        RECT 1023.720 2519.925 1024.620 2936.745 ;
        RECT 1027.020 2519.925 1091.320 2936.745 ;
        RECT 1093.720 2519.925 1094.620 2936.745 ;
        RECT 1097.020 2519.925 1161.320 2936.745 ;
        RECT 1163.720 2519.925 1164.620 2936.745 ;
        RECT 1167.020 2519.925 1231.320 2936.745 ;
        RECT 1003.540 2331.835 1231.320 2519.925 ;
        RECT 1003.540 2314.080 1021.320 2331.835 ;
        RECT 957.020 2290.880 1021.320 2314.080 ;
        RECT 957.020 2287.820 1006.660 2290.880 ;
        RECT 953.720 2090.740 1006.660 2287.820 ;
        RECT 953.720 2017.820 954.620 2090.740 ;
        RECT 957.020 2077.440 1006.660 2090.740 ;
        RECT 1009.060 2077.440 1021.320 2290.880 ;
        RECT 957.020 2035.200 1021.320 2077.440 ;
        RECT 957.020 2017.820 997.460 2035.200 ;
        RECT 953.720 1820.740 997.460 2017.820 ;
        RECT 953.720 1777.820 954.620 1820.740 ;
        RECT 957.020 1805.440 997.460 1820.740 ;
        RECT 999.860 1805.440 1001.140 2035.200 ;
        RECT 1003.540 2009.925 1021.320 2035.200 ;
        RECT 1023.720 2009.925 1024.620 2331.835 ;
        RECT 1027.020 2269.925 1091.320 2331.835 ;
        RECT 1093.720 2269.925 1094.620 2331.835 ;
        RECT 1097.020 2269.925 1161.320 2331.835 ;
        RECT 1163.720 2269.925 1164.620 2331.835 ;
        RECT 1167.020 2269.925 1231.320 2331.835 ;
        RECT 1027.020 2085.915 1231.320 2269.925 ;
        RECT 1027.020 2009.925 1091.320 2085.915 ;
        RECT 1093.720 2009.925 1094.620 2085.915 ;
        RECT 1097.020 2009.925 1161.320 2085.915 ;
        RECT 1163.720 2009.925 1164.620 2085.915 ;
        RECT 1167.020 2009.925 1231.320 2085.915 ;
        RECT 1003.540 1821.835 1231.320 2009.925 ;
        RECT 1003.540 1805.440 1021.320 1821.835 ;
        RECT 957.020 1784.960 1021.320 1805.440 ;
        RECT 957.020 1777.820 1006.660 1784.960 ;
        RECT 953.720 1756.325 1006.660 1777.820 ;
        RECT 747.020 1582.515 1006.660 1756.325 ;
        RECT 747.020 1246.325 811.320 1582.515 ;
        RECT 813.720 1246.325 814.620 1582.515 ;
        RECT 817.020 1246.325 881.320 1582.515 ;
        RECT 883.720 1246.325 884.620 1582.515 ;
        RECT 887.020 1246.325 951.320 1582.515 ;
        RECT 953.720 1580.740 1006.660 1582.515 ;
        RECT 953.720 1507.820 954.620 1580.740 ;
        RECT 957.020 1566.080 1006.660 1580.740 ;
        RECT 1009.060 1566.080 1021.320 1784.960 ;
        RECT 957.020 1523.840 1021.320 1566.080 ;
        RECT 957.020 1507.820 997.460 1523.840 ;
        RECT 953.720 1310.740 997.460 1507.820 ;
        RECT 953.720 1267.820 954.620 1310.740 ;
        RECT 957.020 1294.080 997.460 1310.740 ;
        RECT 999.860 1294.080 1001.140 1523.840 ;
        RECT 1003.540 1499.925 1021.320 1523.840 ;
        RECT 1023.720 1499.925 1024.620 1821.835 ;
        RECT 1027.020 1499.925 1091.320 1821.835 ;
        RECT 1093.720 1499.925 1094.620 1821.835 ;
        RECT 1097.020 1499.925 1161.320 1821.835 ;
        RECT 1163.720 1499.925 1164.620 1821.835 ;
        RECT 1167.020 1499.925 1231.320 1821.835 ;
        RECT 1003.540 1311.835 1231.320 1499.925 ;
        RECT 1003.540 1294.080 1021.320 1311.835 ;
        RECT 957.020 1273.600 1021.320 1294.080 ;
        RECT 957.020 1267.820 1006.660 1273.600 ;
        RECT 953.720 1246.325 1006.660 1267.820 ;
        RECT 747.020 1072.515 1006.660 1246.325 ;
        RECT 747.020 736.325 811.320 1072.515 ;
        RECT 813.720 736.325 814.620 1072.515 ;
        RECT 817.020 736.325 881.320 1072.515 ;
        RECT 883.720 736.325 884.620 1072.515 ;
        RECT 887.020 736.325 951.320 1072.515 ;
        RECT 953.720 1070.740 1006.660 1072.515 ;
        RECT 953.720 997.820 954.620 1070.740 ;
        RECT 957.020 1054.720 1006.660 1070.740 ;
        RECT 1009.060 1054.720 1021.320 1273.600 ;
        RECT 957.020 1015.200 1021.320 1054.720 ;
        RECT 957.020 997.820 997.460 1015.200 ;
        RECT 953.720 800.740 997.460 997.820 ;
        RECT 953.720 757.820 954.620 800.740 ;
        RECT 957.020 785.440 997.460 800.740 ;
        RECT 999.860 785.440 1001.140 1015.200 ;
        RECT 1003.540 989.925 1021.320 1015.200 ;
        RECT 1023.720 989.925 1024.620 1311.835 ;
        RECT 1027.020 989.925 1091.320 1311.835 ;
        RECT 1093.720 989.925 1094.620 1311.835 ;
        RECT 1097.020 989.925 1161.320 1311.835 ;
        RECT 1163.720 989.925 1164.620 1311.835 ;
        RECT 1167.020 989.925 1231.320 1311.835 ;
        RECT 1003.540 801.835 1231.320 989.925 ;
        RECT 1003.540 785.440 1021.320 801.835 ;
        RECT 957.020 762.240 1021.320 785.440 ;
        RECT 957.020 757.820 1006.660 762.240 ;
        RECT 953.720 736.325 1006.660 757.820 ;
        RECT 747.020 562.515 1006.660 736.325 ;
        RECT 747.020 471.285 811.320 562.515 ;
        RECT 813.720 471.285 814.620 562.515 ;
        RECT 817.020 471.285 881.320 562.515 ;
        RECT 883.720 471.285 884.620 562.515 ;
        RECT 887.020 471.285 951.320 562.515 ;
        RECT 747.020 317.875 951.320 471.285 ;
        RECT 747.020 11.735 811.320 317.875 ;
        RECT 813.720 11.735 814.620 317.875 ;
        RECT 817.020 11.735 881.320 317.875 ;
        RECT 883.720 11.735 884.620 317.875 ;
        RECT 887.020 11.735 951.320 317.875 ;
        RECT 953.720 560.740 1006.660 562.515 ;
        RECT 953.720 477.820 954.620 560.740 ;
        RECT 957.020 548.800 1006.660 560.740 ;
        RECT 1009.060 548.800 1021.320 762.240 ;
        RECT 957.020 495.680 1021.320 548.800 ;
        RECT 957.020 477.820 1006.660 495.680 ;
        RECT 953.720 280.740 1006.660 477.820 ;
        RECT 953.720 11.735 954.620 280.740 ;
        RECT 957.020 265.920 1006.660 280.740 ;
        RECT 1009.060 265.920 1021.320 495.680 ;
        RECT 957.020 11.735 1021.320 265.920 ;
        RECT 1023.720 11.735 1024.620 801.835 ;
        RECT 1027.020 11.735 1091.320 801.835 ;
        RECT 1093.720 11.735 1094.620 801.835 ;
        RECT 1097.020 386.965 1161.320 801.835 ;
        RECT 1163.720 386.965 1164.620 801.835 ;
        RECT 1167.020 386.965 1231.320 801.835 ;
        RECT 1097.020 282.515 1231.320 386.965 ;
        RECT 1097.020 11.735 1161.320 282.515 ;
        RECT 1163.720 11.735 1164.620 282.515 ;
        RECT 1167.020 11.735 1231.320 282.515 ;
        RECT 1233.720 11.735 1234.620 2936.745 ;
        RECT 1237.020 2543.840 1301.320 2936.745 ;
        RECT 1237.020 2314.080 1262.420 2543.840 ;
        RECT 1264.820 2314.080 1266.100 2543.840 ;
        RECT 1268.500 2314.080 1301.320 2543.840 ;
        RECT 1237.020 2293.600 1301.320 2314.080 ;
        RECT 1237.020 2074.720 1254.140 2293.600 ;
        RECT 1256.540 2074.720 1257.820 2293.600 ;
        RECT 1260.220 2286.725 1301.320 2293.600 ;
        RECT 1303.720 2286.725 1304.620 2936.745 ;
        RECT 1307.020 2286.725 1371.320 2936.745 ;
        RECT 1373.720 2286.725 1374.620 2936.745 ;
        RECT 1377.020 2286.725 1441.320 2936.745 ;
        RECT 1260.220 2093.195 1441.320 2286.725 ;
        RECT 1260.220 2074.720 1301.320 2093.195 ;
        RECT 1237.020 2035.200 1301.320 2074.720 ;
        RECT 1237.020 1805.440 1262.420 2035.200 ;
        RECT 1264.820 1805.440 1266.100 2035.200 ;
        RECT 1268.500 1805.440 1301.320 2035.200 ;
        RECT 1237.020 1782.240 1301.320 1805.440 ;
        RECT 1237.020 1568.800 1255.980 1782.240 ;
        RECT 1258.380 1756.325 1301.320 1782.240 ;
        RECT 1303.720 1756.325 1304.620 2093.195 ;
        RECT 1307.020 1756.325 1371.320 2093.195 ;
        RECT 1373.720 1756.325 1374.620 2093.195 ;
        RECT 1377.020 1756.325 1441.320 2093.195 ;
        RECT 1443.720 1756.325 1444.620 2936.745 ;
        RECT 1447.020 1756.325 1511.320 2936.745 ;
        RECT 1258.380 1582.515 1511.320 1756.325 ;
        RECT 1258.380 1568.800 1301.320 1582.515 ;
        RECT 1237.020 1523.840 1301.320 1568.800 ;
        RECT 1237.020 1294.080 1262.420 1523.840 ;
        RECT 1264.820 1294.080 1266.100 1523.840 ;
        RECT 1268.500 1294.080 1301.320 1523.840 ;
        RECT 1237.020 1270.880 1301.320 1294.080 ;
        RECT 1237.020 1054.720 1254.140 1270.880 ;
        RECT 1256.540 1054.720 1257.820 1270.880 ;
        RECT 1260.220 1246.325 1301.320 1270.880 ;
        RECT 1303.720 1246.325 1304.620 1582.515 ;
        RECT 1307.020 1246.325 1371.320 1582.515 ;
        RECT 1373.720 1246.325 1374.620 1582.515 ;
        RECT 1377.020 1246.325 1441.320 1582.515 ;
        RECT 1443.720 1246.325 1444.620 1582.515 ;
        RECT 1447.020 1246.325 1511.320 1582.515 ;
        RECT 1260.220 1072.515 1511.320 1246.325 ;
        RECT 1260.220 1054.720 1301.320 1072.515 ;
        RECT 1237.020 1015.200 1301.320 1054.720 ;
        RECT 1237.020 785.440 1262.420 1015.200 ;
        RECT 1264.820 785.440 1266.100 1015.200 ;
        RECT 1268.500 785.440 1301.320 1015.200 ;
        RECT 1237.020 764.960 1301.320 785.440 ;
        RECT 1237.020 546.080 1254.140 764.960 ;
        RECT 1256.540 546.080 1257.820 764.960 ;
        RECT 1260.220 736.325 1301.320 764.960 ;
        RECT 1303.720 736.325 1304.620 1072.515 ;
        RECT 1307.020 736.325 1371.320 1072.515 ;
        RECT 1373.720 736.325 1374.620 1072.515 ;
        RECT 1377.020 736.325 1441.320 1072.515 ;
        RECT 1443.720 736.325 1444.620 1072.515 ;
        RECT 1447.020 736.325 1511.320 1072.515 ;
        RECT 1260.220 562.515 1511.320 736.325 ;
        RECT 1260.220 546.080 1301.320 562.515 ;
        RECT 1237.020 492.960 1301.320 546.080 ;
        RECT 1237.020 268.640 1254.140 492.960 ;
        RECT 1256.540 268.640 1257.820 492.960 ;
        RECT 1260.220 471.285 1301.320 492.960 ;
        RECT 1303.720 471.285 1304.620 562.515 ;
        RECT 1307.020 471.285 1371.320 562.515 ;
        RECT 1373.720 471.285 1374.620 562.515 ;
        RECT 1377.020 471.285 1441.320 562.515 ;
        RECT 1260.220 317.875 1441.320 471.285 ;
        RECT 1260.220 268.640 1301.320 317.875 ;
        RECT 1237.020 11.735 1301.320 268.640 ;
        RECT 1303.720 11.735 1304.620 317.875 ;
        RECT 1307.020 11.735 1371.320 317.875 ;
        RECT 1373.720 11.735 1374.620 317.875 ;
        RECT 1377.020 11.735 1441.320 317.875 ;
        RECT 1443.720 11.735 1444.620 562.515 ;
        RECT 1447.020 11.735 1511.320 562.515 ;
        RECT 1513.720 11.735 1514.620 2936.745 ;
        RECT 1517.020 2519.925 1581.320 2936.745 ;
        RECT 1583.720 2807.820 1584.620 2936.745 ;
        RECT 1587.020 2807.820 1651.320 2936.745 ;
        RECT 1583.720 2610.740 1651.320 2807.820 ;
        RECT 1583.720 2519.925 1584.620 2610.740 ;
        RECT 1587.020 2519.925 1651.320 2610.740 ;
        RECT 1653.720 2519.925 1654.620 2936.745 ;
        RECT 1657.020 2519.925 1721.320 2936.745 ;
        RECT 1723.720 2519.925 1724.620 2936.745 ;
        RECT 1727.020 2543.840 1791.320 2936.745 ;
        RECT 1727.020 2519.925 1772.100 2543.840 ;
        RECT 1517.020 2331.835 1772.100 2519.925 ;
        RECT 1517.020 2009.925 1581.320 2331.835 ;
        RECT 1583.720 2009.925 1584.620 2331.835 ;
        RECT 1587.020 2269.925 1651.320 2331.835 ;
        RECT 1653.720 2269.925 1654.620 2331.835 ;
        RECT 1657.020 2269.925 1721.320 2331.835 ;
        RECT 1587.020 2085.915 1721.320 2269.925 ;
        RECT 1587.020 2009.925 1651.320 2085.915 ;
        RECT 1653.720 2009.925 1654.620 2085.915 ;
        RECT 1657.020 2009.925 1721.320 2085.915 ;
        RECT 1723.720 2009.925 1724.620 2331.835 ;
        RECT 1727.020 2314.080 1772.100 2331.835 ;
        RECT 1774.500 2314.080 1775.780 2543.840 ;
        RECT 1778.180 2314.080 1791.320 2543.840 ;
        RECT 1727.020 2293.600 1791.320 2314.080 ;
        RECT 1727.020 2074.720 1764.740 2293.600 ;
        RECT 1767.140 2074.720 1768.420 2293.600 ;
        RECT 1770.820 2074.720 1791.320 2293.600 ;
        RECT 1727.020 2035.200 1791.320 2074.720 ;
        RECT 1727.020 2009.925 1772.100 2035.200 ;
        RECT 1517.020 1821.835 1772.100 2009.925 ;
        RECT 1517.020 1499.925 1581.320 1821.835 ;
        RECT 1583.720 1499.925 1584.620 1821.835 ;
        RECT 1587.020 1499.925 1651.320 1821.835 ;
        RECT 1653.720 1499.925 1654.620 1821.835 ;
        RECT 1657.020 1499.925 1721.320 1821.835 ;
        RECT 1723.720 1499.925 1724.620 1821.835 ;
        RECT 1727.020 1805.440 1772.100 1821.835 ;
        RECT 1774.500 1805.440 1775.780 2035.200 ;
        RECT 1778.180 1805.440 1791.320 2035.200 ;
        RECT 1727.020 1784.960 1791.320 1805.440 ;
        RECT 1727.020 1566.080 1764.740 1784.960 ;
        RECT 1767.140 1566.080 1768.420 1784.960 ;
        RECT 1770.820 1566.080 1791.320 1784.960 ;
        RECT 1727.020 1523.840 1791.320 1566.080 ;
        RECT 1727.020 1499.925 1772.100 1523.840 ;
        RECT 1517.020 1311.835 1772.100 1499.925 ;
        RECT 1517.020 989.925 1581.320 1311.835 ;
        RECT 1583.720 989.925 1584.620 1311.835 ;
        RECT 1587.020 989.925 1651.320 1311.835 ;
        RECT 1653.720 989.925 1654.620 1311.835 ;
        RECT 1657.020 989.925 1721.320 1311.835 ;
        RECT 1723.720 989.925 1724.620 1311.835 ;
        RECT 1727.020 1294.080 1772.100 1311.835 ;
        RECT 1774.500 1294.080 1775.780 1523.840 ;
        RECT 1778.180 1294.080 1791.320 1523.840 ;
        RECT 1727.020 1273.600 1791.320 1294.080 ;
        RECT 1727.020 1054.720 1764.740 1273.600 ;
        RECT 1767.140 1054.720 1768.420 1273.600 ;
        RECT 1770.820 1054.720 1791.320 1273.600 ;
        RECT 1727.020 1015.200 1791.320 1054.720 ;
        RECT 1727.020 989.925 1772.100 1015.200 ;
        RECT 1517.020 801.835 1772.100 989.925 ;
        RECT 1517.020 11.735 1581.320 801.835 ;
        RECT 1583.720 227.820 1584.620 801.835 ;
        RECT 1587.020 386.965 1651.320 801.835 ;
        RECT 1653.720 386.965 1654.620 801.835 ;
        RECT 1657.020 386.965 1721.320 801.835 ;
        RECT 1723.720 386.965 1724.620 801.835 ;
        RECT 1727.020 785.440 1772.100 801.835 ;
        RECT 1774.500 785.440 1775.780 1015.200 ;
        RECT 1778.180 785.440 1791.320 1015.200 ;
        RECT 1727.020 775.840 1791.320 785.440 ;
        RECT 1727.020 546.080 1764.740 775.840 ;
        RECT 1767.140 546.080 1768.420 775.840 ;
        RECT 1770.820 546.080 1791.320 775.840 ;
        RECT 1727.020 495.680 1791.320 546.080 ;
        RECT 1727.020 386.965 1764.740 495.680 ;
        RECT 1587.020 282.515 1764.740 386.965 ;
        RECT 1587.020 227.820 1651.320 282.515 ;
        RECT 1583.720 30.740 1651.320 227.820 ;
        RECT 1583.720 11.735 1584.620 30.740 ;
        RECT 1587.020 11.735 1651.320 30.740 ;
        RECT 1653.720 11.735 1654.620 282.515 ;
        RECT 1657.020 11.735 1721.320 282.515 ;
        RECT 1723.720 11.735 1724.620 282.515 ;
        RECT 1727.020 265.920 1764.740 282.515 ;
        RECT 1767.140 265.920 1768.420 495.680 ;
        RECT 1770.820 265.920 1791.320 495.680 ;
        RECT 1727.020 11.735 1791.320 265.920 ;
        RECT 1793.720 2286.725 1794.620 2936.745 ;
        RECT 1797.020 2286.725 1861.320 2936.745 ;
        RECT 1863.720 2286.725 1864.620 2936.745 ;
        RECT 1867.020 2286.725 1931.320 2936.745 ;
        RECT 1933.720 2286.725 1934.620 2936.745 ;
        RECT 1937.020 2286.725 2001.320 2936.745 ;
        RECT 1793.720 2093.195 2001.320 2286.725 ;
        RECT 1793.720 11.735 1794.620 2093.195 ;
        RECT 1797.020 1756.325 1861.320 2093.195 ;
        RECT 1863.720 1756.325 1864.620 2093.195 ;
        RECT 1867.020 1756.325 1931.320 2093.195 ;
        RECT 1933.720 1756.325 1934.620 2093.195 ;
        RECT 1937.020 1756.325 2001.320 2093.195 ;
        RECT 1797.020 1582.515 2001.320 1756.325 ;
        RECT 1797.020 1246.325 1861.320 1582.515 ;
        RECT 1863.720 1246.325 1864.620 1582.515 ;
        RECT 1867.020 1246.325 1931.320 1582.515 ;
        RECT 1933.720 1246.325 1934.620 1582.515 ;
        RECT 1937.020 1246.325 2001.320 1582.515 ;
        RECT 1797.020 1072.515 2001.320 1246.325 ;
        RECT 1797.020 736.325 1861.320 1072.515 ;
        RECT 1863.720 736.325 1864.620 1072.515 ;
        RECT 1867.020 736.325 1931.320 1072.515 ;
        RECT 1933.720 736.325 1934.620 1072.515 ;
        RECT 1937.020 736.325 2001.320 1072.515 ;
        RECT 1797.020 562.515 2001.320 736.325 ;
        RECT 1797.020 471.285 1861.320 562.515 ;
        RECT 1863.720 471.285 1864.620 562.515 ;
        RECT 1867.020 471.285 1931.320 562.515 ;
        RECT 1797.020 317.875 1931.320 471.285 ;
        RECT 1797.020 11.735 1861.320 317.875 ;
        RECT 1863.720 11.735 1864.620 317.875 ;
        RECT 1867.020 11.735 1931.320 317.875 ;
        RECT 1933.720 11.735 1934.620 562.515 ;
        RECT 1937.020 11.735 2001.320 562.515 ;
        RECT 2003.720 11.735 2004.620 2936.745 ;
        RECT 2007.020 2543.840 2071.320 2936.745 ;
        RECT 2007.020 2314.080 2016.820 2543.840 ;
        RECT 2019.220 2314.080 2020.500 2543.840 ;
        RECT 2022.900 2519.925 2071.320 2543.840 ;
        RECT 2073.720 2519.925 2074.620 2936.745 ;
        RECT 2077.020 2519.925 2141.320 2936.745 ;
        RECT 2143.720 2519.925 2144.620 2936.745 ;
        RECT 2147.020 2519.925 2211.320 2936.745 ;
        RECT 2213.720 2546.860 2214.620 2936.745 ;
        RECT 2217.020 2546.860 2281.320 2936.745 ;
        RECT 2213.720 2519.925 2281.320 2546.860 ;
        RECT 2022.900 2331.835 2281.320 2519.925 ;
        RECT 2022.900 2314.080 2071.320 2331.835 ;
        RECT 2007.020 2293.600 2071.320 2314.080 ;
        RECT 2007.020 2074.720 2024.180 2293.600 ;
        RECT 2026.580 2074.720 2027.860 2293.600 ;
        RECT 2030.260 2074.720 2071.320 2293.600 ;
        RECT 2007.020 2035.200 2071.320 2074.720 ;
        RECT 2007.020 1805.440 2016.820 2035.200 ;
        RECT 2019.220 1805.440 2020.500 2035.200 ;
        RECT 2022.900 2009.925 2071.320 2035.200 ;
        RECT 2073.720 2277.820 2074.620 2331.835 ;
        RECT 2077.020 2277.820 2141.320 2331.835 ;
        RECT 2073.720 2269.925 2141.320 2277.820 ;
        RECT 2143.720 2269.925 2144.620 2331.835 ;
        RECT 2147.020 2269.925 2211.320 2331.835 ;
        RECT 2213.720 2330.740 2281.320 2331.835 ;
        RECT 2213.720 2269.925 2214.620 2330.740 ;
        RECT 2073.720 2085.915 2214.620 2269.925 ;
        RECT 2073.720 2080.740 2141.320 2085.915 ;
        RECT 2073.720 2009.925 2074.620 2080.740 ;
        RECT 2077.020 2009.925 2141.320 2080.740 ;
        RECT 2143.720 2009.925 2144.620 2085.915 ;
        RECT 2147.020 2009.925 2211.320 2085.915 ;
        RECT 2213.720 2036.860 2214.620 2085.915 ;
        RECT 2217.020 2036.860 2281.320 2330.740 ;
        RECT 2213.720 2009.925 2281.320 2036.860 ;
        RECT 2022.900 1821.835 2281.320 2009.925 ;
        RECT 2022.900 1805.440 2071.320 1821.835 ;
        RECT 2007.020 1784.960 2071.320 1805.440 ;
        RECT 2007.020 1566.080 2024.180 1784.960 ;
        RECT 2026.580 1566.080 2027.860 1784.960 ;
        RECT 2030.260 1566.080 2071.320 1784.960 ;
        RECT 2007.020 1523.840 2071.320 1566.080 ;
        RECT 2007.020 1294.080 2016.820 1523.840 ;
        RECT 2019.220 1294.080 2020.500 1523.840 ;
        RECT 2022.900 1499.925 2071.320 1523.840 ;
        RECT 2073.720 1767.820 2074.620 1821.835 ;
        RECT 2077.020 1767.820 2141.320 1821.835 ;
        RECT 2073.720 1570.740 2141.320 1767.820 ;
        RECT 2073.720 1499.925 2074.620 1570.740 ;
        RECT 2077.020 1499.925 2141.320 1570.740 ;
        RECT 2143.720 1499.925 2144.620 1821.835 ;
        RECT 2147.020 1499.925 2211.320 1821.835 ;
        RECT 2213.720 1820.740 2281.320 1821.835 ;
        RECT 2213.720 1526.860 2214.620 1820.740 ;
        RECT 2217.020 1526.860 2281.320 1820.740 ;
        RECT 2213.720 1499.925 2281.320 1526.860 ;
        RECT 2022.900 1311.835 2281.320 1499.925 ;
        RECT 2022.900 1294.080 2071.320 1311.835 ;
        RECT 2007.020 1279.040 2071.320 1294.080 ;
        RECT 2007.020 1054.720 2024.180 1279.040 ;
        RECT 2026.580 1054.720 2027.860 1279.040 ;
        RECT 2030.260 1054.720 2071.320 1279.040 ;
        RECT 2007.020 1015.200 2071.320 1054.720 ;
        RECT 2007.020 785.440 2016.820 1015.200 ;
        RECT 2019.220 785.440 2020.500 1015.200 ;
        RECT 2022.900 989.925 2071.320 1015.200 ;
        RECT 2073.720 1260.820 2074.620 1311.835 ;
        RECT 2077.020 1260.820 2141.320 1311.835 ;
        RECT 2073.720 1063.740 2141.320 1260.820 ;
        RECT 2073.720 989.925 2074.620 1063.740 ;
        RECT 2077.020 989.925 2141.320 1063.740 ;
        RECT 2143.720 989.925 2144.620 1311.835 ;
        RECT 2147.020 989.925 2211.320 1311.835 ;
        RECT 2213.720 1310.740 2281.320 1311.835 ;
        RECT 2213.720 1016.860 2214.620 1310.740 ;
        RECT 2217.020 1016.860 2281.320 1310.740 ;
        RECT 2213.720 989.925 2281.320 1016.860 ;
        RECT 2022.900 801.835 2281.320 989.925 ;
        RECT 2022.900 785.440 2071.320 801.835 ;
        RECT 2007.020 764.960 2071.320 785.440 ;
        RECT 2007.020 546.080 2024.180 764.960 ;
        RECT 2026.580 546.080 2027.860 764.960 ;
        RECT 2030.260 546.080 2071.320 764.960 ;
        RECT 2007.020 495.680 2071.320 546.080 ;
        RECT 2007.020 265.920 2024.180 495.680 ;
        RECT 2026.580 265.920 2027.860 495.680 ;
        RECT 2030.260 265.920 2071.320 495.680 ;
        RECT 2007.020 11.735 2071.320 265.920 ;
        RECT 2073.720 747.820 2074.620 801.835 ;
        RECT 2077.020 747.820 2141.320 801.835 ;
        RECT 2073.720 550.740 2141.320 747.820 ;
        RECT 2073.720 477.820 2074.620 550.740 ;
        RECT 2077.020 477.820 2141.320 550.740 ;
        RECT 2073.720 386.965 2141.320 477.820 ;
        RECT 2143.720 386.965 2144.620 801.835 ;
        RECT 2147.020 386.965 2211.320 801.835 ;
        RECT 2213.720 800.740 2281.320 801.835 ;
        RECT 2213.720 386.965 2214.620 800.740 ;
        RECT 2217.020 386.965 2281.320 800.740 ;
        RECT 2073.720 282.515 2281.320 386.965 ;
        RECT 2073.720 280.740 2141.320 282.515 ;
        RECT 2073.720 11.735 2074.620 280.740 ;
        RECT 2077.020 11.735 2141.320 280.740 ;
        RECT 2143.720 11.735 2144.620 282.515 ;
        RECT 2147.020 11.735 2211.320 282.515 ;
        RECT 2213.720 11.735 2214.620 282.515 ;
        RECT 2217.020 11.735 2281.320 282.515 ;
        RECT 2283.720 11.735 2284.620 2936.745 ;
        RECT 2287.020 2393.125 2351.320 2936.745 ;
        RECT 2353.720 2393.125 2354.620 2936.745 ;
        RECT 2357.020 2393.125 2421.320 2936.745 ;
        RECT 2287.020 2308.395 2421.320 2393.125 ;
        RECT 2287.020 1883.125 2351.320 2308.395 ;
        RECT 2353.720 1883.125 2354.620 2308.395 ;
        RECT 2357.020 2171.445 2421.320 2308.395 ;
        RECT 2423.720 2188.860 2424.620 2936.745 ;
        RECT 2427.020 2188.860 2491.320 2936.745 ;
        RECT 2423.720 2171.445 2491.320 2188.860 ;
        RECT 2357.020 2047.955 2491.320 2171.445 ;
        RECT 2357.020 1883.125 2421.320 2047.955 ;
        RECT 2287.020 1798.395 2421.320 1883.125 ;
        RECT 2287.020 1724.005 2351.320 1798.395 ;
        RECT 2353.720 1724.005 2354.620 1798.395 ;
        RECT 2357.020 1724.005 2421.320 1798.395 ;
        RECT 2423.720 2040.740 2491.320 2047.955 ;
        RECT 2423.720 1724.005 2424.620 2040.740 ;
        RECT 2427.020 1724.005 2491.320 2040.740 ;
        RECT 2287.020 1532.515 2491.320 1724.005 ;
        RECT 2287.020 1373.125 2351.320 1532.515 ;
        RECT 2353.720 1373.125 2354.620 1532.515 ;
        RECT 2357.020 1373.125 2421.320 1532.515 ;
        RECT 2287.020 1288.395 2421.320 1373.125 ;
        RECT 2287.020 1214.005 2351.320 1288.395 ;
        RECT 2353.720 1214.005 2354.620 1288.395 ;
        RECT 2357.020 1214.005 2421.320 1288.395 ;
        RECT 2423.720 1214.005 2424.620 1532.515 ;
        RECT 2427.020 1214.005 2491.320 1532.515 ;
        RECT 2287.020 1022.515 2491.320 1214.005 ;
        RECT 2287.020 863.125 2351.320 1022.515 ;
        RECT 2353.720 863.125 2354.620 1022.515 ;
        RECT 2357.020 863.125 2421.320 1022.515 ;
        RECT 2287.020 778.395 2421.320 863.125 ;
        RECT 2287.020 704.005 2351.320 778.395 ;
        RECT 2353.720 704.005 2354.620 778.395 ;
        RECT 2357.020 704.005 2421.320 778.395 ;
        RECT 2423.720 704.005 2424.620 1022.515 ;
        RECT 2427.020 704.005 2491.320 1022.515 ;
        RECT 2287.020 512.515 2491.320 704.005 ;
        RECT 2287.020 472.645 2351.320 512.515 ;
        RECT 2353.720 472.645 2354.620 512.515 ;
        RECT 2357.020 472.645 2421.320 512.515 ;
        RECT 2287.020 289.995 2421.320 472.645 ;
        RECT 2287.020 11.735 2351.320 289.995 ;
        RECT 2353.720 11.735 2354.620 289.995 ;
        RECT 2357.020 11.735 2421.320 289.995 ;
        RECT 2423.720 11.735 2424.620 512.515 ;
        RECT 2427.020 11.735 2491.320 512.515 ;
        RECT 2493.720 2188.860 2494.620 2936.745 ;
        RECT 2497.020 2508.480 2561.320 2936.745 ;
        RECT 2497.020 2295.040 2532.020 2508.480 ;
        RECT 2534.420 2295.040 2535.700 2508.480 ;
        RECT 2538.100 2295.040 2561.320 2508.480 ;
        RECT 2497.020 2188.860 2561.320 2295.040 ;
        RECT 2493.720 2040.740 2561.320 2188.860 ;
        RECT 2493.720 11.735 2494.620 2040.740 ;
        RECT 2497.020 1999.840 2561.320 2040.740 ;
        RECT 2497.020 1786.400 2532.020 1999.840 ;
        RECT 2534.420 1786.400 2535.700 1999.840 ;
        RECT 2538.100 1786.400 2561.320 1999.840 ;
        RECT 2497.020 1488.480 2561.320 1786.400 ;
        RECT 2497.020 1275.040 2532.020 1488.480 ;
        RECT 2534.420 1275.040 2535.700 1488.480 ;
        RECT 2538.100 1275.040 2561.320 1488.480 ;
        RECT 2497.020 979.840 2561.320 1275.040 ;
        RECT 2497.020 766.400 2532.020 979.840 ;
        RECT 2534.420 766.400 2535.700 979.840 ;
        RECT 2538.100 766.400 2561.320 979.840 ;
        RECT 2497.020 11.735 2561.320 766.400 ;
        RECT 2563.720 11.735 2564.620 2936.745 ;
        RECT 2567.020 11.735 2631.320 2936.745 ;
        RECT 2633.720 11.735 2634.620 2936.745 ;
        RECT 2637.020 11.735 2701.320 2936.745 ;
        RECT 2703.720 11.735 2704.620 2936.745 ;
        RECT 2707.020 11.735 2767.065 2936.745 ;
      LAYER met5 ;
        RECT 35.540 2603.580 2583.700 2668.100 ;
        RECT 35.540 2528.580 2583.700 2595.480 ;
        RECT 35.540 2453.580 2583.700 2520.480 ;
        RECT 518.980 2445.480 631.660 2453.580 ;
        RECT 1028.980 2445.480 1141.660 2453.580 ;
        RECT 1538.980 2445.480 1651.660 2453.580 ;
        RECT 2048.980 2445.480 2161.660 2453.580 ;
        RECT 35.540 2378.580 2583.700 2445.480 ;
        RECT 35.540 2303.580 2583.700 2370.480 ;
        RECT 35.540 2228.580 2583.700 2295.480 ;
        RECT 35.540 2153.580 2583.700 2220.480 ;
        RECT 35.540 2078.580 2583.700 2145.480 ;
        RECT 35.540 2003.580 2583.700 2070.480 ;
        RECT 35.540 1928.580 2583.700 1995.480 ;
        RECT 518.980 1920.480 631.660 1928.580 ;
        RECT 1028.980 1920.480 1141.660 1928.580 ;
        RECT 1538.980 1920.480 1651.660 1928.580 ;
        RECT 2048.980 1920.480 2161.660 1928.580 ;
        RECT 35.540 1853.580 2583.700 1920.480 ;
        RECT 35.540 1778.580 2583.700 1845.480 ;
        RECT 35.540 1703.580 2583.700 1770.480 ;
        RECT 35.540 1628.580 2583.700 1695.480 ;
        RECT 35.540 1553.580 2583.700 1620.480 ;
        RECT 2358.980 1545.480 2485.460 1553.580 ;
        RECT 35.540 1478.580 2583.700 1545.480 ;
        RECT 518.980 1470.480 631.660 1478.580 ;
        RECT 1028.980 1470.480 1141.660 1478.580 ;
        RECT 1538.980 1470.480 1651.660 1478.580 ;
        RECT 2048.980 1470.480 2161.660 1478.580 ;
        RECT 35.540 1403.580 2583.700 1470.480 ;
        RECT 518.980 1395.480 631.660 1403.580 ;
        RECT 1028.980 1395.480 1141.660 1403.580 ;
        RECT 1538.980 1395.480 1651.660 1403.580 ;
        RECT 2048.980 1395.480 2161.660 1403.580 ;
        RECT 35.540 1328.580 2583.700 1395.480 ;
        RECT 35.540 1292.700 2583.700 1320.480 ;
        RECT 35.540 1284.500 250.120 1292.700 ;
        RECT 398.220 1284.500 2583.700 1292.700 ;
        RECT 35.540 1253.580 2583.700 1284.500 ;
        RECT 35.540 1178.580 2583.700 1245.480 ;
        RECT 35.540 1103.580 2583.700 1170.480 ;
        RECT 35.540 1028.580 2583.700 1095.480 ;
        RECT 2358.980 1025.280 2485.460 1028.580 ;
        RECT 35.540 953.580 2583.700 1020.480 ;
        RECT 518.980 945.480 631.660 953.580 ;
        RECT 1028.980 945.480 1141.660 953.580 ;
        RECT 1538.980 945.480 1651.660 953.580 ;
        RECT 2048.980 945.480 2161.660 953.580 ;
        RECT 35.540 878.580 2583.700 945.480 ;
        RECT 35.540 803.580 2583.700 870.480 ;
        RECT 35.540 728.580 2583.700 795.480 ;
        RECT 35.540 653.580 2583.700 720.480 ;
        RECT 35.540 578.580 2583.700 645.480 ;
        RECT 35.540 503.580 2583.700 570.480 ;
        RECT 35.540 428.580 2583.700 495.480 ;
        RECT 35.540 353.580 2583.700 420.480 ;
        RECT 35.540 278.580 2583.700 345.480 ;
        RECT 35.540 203.580 2583.700 270.480 ;
        RECT 35.540 128.580 2583.700 195.480 ;
        RECT 35.540 85.900 2583.700 120.480 ;
  END
END fpga_top
END LIBRARY

