VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__1_
  CLASS BLOCK ;
  FOREIGN cbx_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 190.000 BY 200.000 ;
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 156.440 4.000 157.040 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 129.240 189.000 129.840 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 176.840 189.000 177.440 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
  PIN bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 71.440 4.000 72.040 ;
    END
  END bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 156.440 189.000 157.040 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1.000 67.990 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 37.440 189.000 38.040 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1.000 42.230 4.000 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 139.440 189.000 140.040 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1.000 93.750 4.000 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.840 4.000 109.440 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 193.840 189.000 194.440 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 119.040 189.000 119.640 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1.000 180.690 4.000 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 196.000 26.130 199.000 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 199.000 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 196.000 106.630 199.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 10.240 189.000 10.840 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1.000 174.250 4.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 74.840 189.000 75.440 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1.000 164.590 4.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 196.000 122.730 199.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 196.000 10.030 199.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 196.000 80.870 199.000 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 119.040 4.000 119.640 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 149.640 189.000 150.240 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 6.840 4.000 7.440 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 146.240 4.000 146.840 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 196.000 142.050 199.000 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 17.040 4.000 17.640 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 196.000 174.250 199.000 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 85.040 189.000 85.640 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 196.000 96.970 199.000 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1.000 113.070 4.000 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.640 4.000 184.240 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 199.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 64.640 189.000 65.240 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 196.000 0.370 199.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1.000 148.490 4.000 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1.000 77.650 4.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 34.040 4.000 34.640 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 166.640 189.000 167.240 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 44.240 4.000 44.840 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1.000 16.470 4.000 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1.000 51.890 4.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1.000 154.930 4.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 54.440 189.000 55.040 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 27.240 189.000 27.840 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1.000 119.510 4.000 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.440 4.000 191.040 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 0.040 189.000 0.640 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 196.000 51.890 199.000 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 47.640 189.000 48.240 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 125.840 4.000 126.440 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1.000 138.830 4.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 91.840 4.000 92.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 196.000 35.790 199.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 196.000 71.210 199.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 163.240 4.000 163.840 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 98.640 4.000 99.240 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 196.000 61.550 199.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 196.000 113.070 199.000 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 196.000 167.810 199.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 136.040 4.000 136.640 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1.000 26.130 4.000 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1.000 6.810 4.000 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 196.000 183.910 199.000 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 27.240 4.000 27.840 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1.000 87.310 4.000 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 183.640 189.000 184.240 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 20.440 189.000 21.040 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 54.440 4.000 55.040 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 102.040 189.000 102.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1.000 32.570 4.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1.000 58.330 4.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 81.640 4.000 82.240 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 112.240 189.000 112.840 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1.000 103.410 4.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 196.000 158.150 199.000 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 196.000 148.490 199.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 196.000 19.690 199.000 ;
    END
  END chanx_right_out[9]
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 196.000 45.450 199.000 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1.000 129.170 4.000 ;
    END
  END prog_clk
  PIN top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 61.240 4.000 61.840 ;
    END
  END top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
  PIN top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 173.440 4.000 174.040 ;
    END
  END top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
  PIN top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 186.000 91.840 189.000 92.440 ;
    END
  END top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 184.460 187.765 ;
      LAYER met1 ;
        RECT 0.070 9.220 184.460 187.920 ;
      LAYER met2 ;
        RECT 0.650 195.720 9.470 196.000 ;
        RECT 10.310 195.720 19.130 196.000 ;
        RECT 19.970 195.720 25.570 196.000 ;
        RECT 26.410 195.720 35.230 196.000 ;
        RECT 36.070 195.720 44.890 196.000 ;
        RECT 45.730 195.720 51.330 196.000 ;
        RECT 52.170 195.720 60.990 196.000 ;
        RECT 61.830 195.720 70.650 196.000 ;
        RECT 71.490 195.720 80.310 196.000 ;
        RECT 81.150 195.720 86.750 196.000 ;
        RECT 87.590 195.720 96.410 196.000 ;
        RECT 97.250 195.720 106.070 196.000 ;
        RECT 106.910 195.720 112.510 196.000 ;
        RECT 113.350 195.720 122.170 196.000 ;
        RECT 123.010 195.720 131.830 196.000 ;
        RECT 132.670 195.720 141.490 196.000 ;
        RECT 142.330 195.720 147.930 196.000 ;
        RECT 148.770 195.720 157.590 196.000 ;
        RECT 158.430 195.720 167.250 196.000 ;
        RECT 168.090 195.720 173.690 196.000 ;
        RECT 174.530 195.720 183.350 196.000 ;
        RECT 0.100 4.280 183.900 195.720 ;
        RECT 0.650 0.720 6.250 4.280 ;
        RECT 7.090 0.720 15.910 4.280 ;
        RECT 16.750 0.720 25.570 4.280 ;
        RECT 26.410 0.720 32.010 4.280 ;
        RECT 32.850 0.720 41.670 4.280 ;
        RECT 42.510 0.720 51.330 4.280 ;
        RECT 52.170 0.720 57.770 4.280 ;
        RECT 58.610 0.720 67.430 4.280 ;
        RECT 68.270 0.720 77.090 4.280 ;
        RECT 77.930 0.720 86.750 4.280 ;
        RECT 87.590 0.720 93.190 4.280 ;
        RECT 94.030 0.720 102.850 4.280 ;
        RECT 103.690 0.720 112.510 4.280 ;
        RECT 113.350 0.720 118.950 4.280 ;
        RECT 119.790 0.720 128.610 4.280 ;
        RECT 129.450 0.720 138.270 4.280 ;
        RECT 139.110 0.720 147.930 4.280 ;
        RECT 148.770 0.720 154.370 4.280 ;
        RECT 155.210 0.720 164.030 4.280 ;
        RECT 164.870 0.720 173.690 4.280 ;
        RECT 174.530 0.720 180.130 4.280 ;
        RECT 180.970 0.720 183.900 4.280 ;
        RECT 0.100 0.155 183.900 0.720 ;
      LAYER met3 ;
        RECT 4.000 193.440 185.600 194.305 ;
        RECT 4.000 191.440 186.000 193.440 ;
        RECT 4.400 190.040 186.000 191.440 ;
        RECT 4.000 184.640 186.000 190.040 ;
        RECT 4.400 183.240 185.600 184.640 ;
        RECT 4.000 177.840 186.000 183.240 ;
        RECT 4.000 176.440 185.600 177.840 ;
        RECT 4.000 174.440 186.000 176.440 ;
        RECT 4.400 173.040 186.000 174.440 ;
        RECT 4.000 167.640 186.000 173.040 ;
        RECT 4.000 166.240 185.600 167.640 ;
        RECT 4.000 164.240 186.000 166.240 ;
        RECT 4.400 162.840 186.000 164.240 ;
        RECT 4.000 157.440 186.000 162.840 ;
        RECT 4.400 156.040 185.600 157.440 ;
        RECT 4.000 150.640 186.000 156.040 ;
        RECT 4.000 149.240 185.600 150.640 ;
        RECT 4.000 147.240 186.000 149.240 ;
        RECT 4.400 145.840 186.000 147.240 ;
        RECT 4.000 140.440 186.000 145.840 ;
        RECT 4.000 139.040 185.600 140.440 ;
        RECT 4.000 137.040 186.000 139.040 ;
        RECT 4.400 135.640 186.000 137.040 ;
        RECT 4.000 130.240 186.000 135.640 ;
        RECT 4.000 128.840 185.600 130.240 ;
        RECT 4.000 126.840 186.000 128.840 ;
        RECT 4.400 125.440 186.000 126.840 ;
        RECT 4.000 120.040 186.000 125.440 ;
        RECT 4.400 118.640 185.600 120.040 ;
        RECT 4.000 113.240 186.000 118.640 ;
        RECT 4.000 111.840 185.600 113.240 ;
        RECT 4.000 109.840 186.000 111.840 ;
        RECT 4.400 108.440 186.000 109.840 ;
        RECT 4.000 103.040 186.000 108.440 ;
        RECT 4.000 101.640 185.600 103.040 ;
        RECT 4.000 99.640 186.000 101.640 ;
        RECT 4.400 98.240 186.000 99.640 ;
        RECT 4.000 92.840 186.000 98.240 ;
        RECT 4.400 91.440 185.600 92.840 ;
        RECT 4.000 86.040 186.000 91.440 ;
        RECT 4.000 84.640 185.600 86.040 ;
        RECT 4.000 82.640 186.000 84.640 ;
        RECT 4.400 81.240 186.000 82.640 ;
        RECT 4.000 75.840 186.000 81.240 ;
        RECT 4.000 74.440 185.600 75.840 ;
        RECT 4.000 72.440 186.000 74.440 ;
        RECT 4.400 71.040 186.000 72.440 ;
        RECT 4.000 65.640 186.000 71.040 ;
        RECT 4.000 64.240 185.600 65.640 ;
        RECT 4.000 62.240 186.000 64.240 ;
        RECT 4.400 60.840 186.000 62.240 ;
        RECT 4.000 55.440 186.000 60.840 ;
        RECT 4.400 54.040 185.600 55.440 ;
        RECT 4.000 48.640 186.000 54.040 ;
        RECT 4.000 47.240 185.600 48.640 ;
        RECT 4.000 45.240 186.000 47.240 ;
        RECT 4.400 43.840 186.000 45.240 ;
        RECT 4.000 38.440 186.000 43.840 ;
        RECT 4.000 37.040 185.600 38.440 ;
        RECT 4.000 35.040 186.000 37.040 ;
        RECT 4.400 33.640 186.000 35.040 ;
        RECT 4.000 28.240 186.000 33.640 ;
        RECT 4.400 26.840 185.600 28.240 ;
        RECT 4.000 21.440 186.000 26.840 ;
        RECT 4.000 20.040 185.600 21.440 ;
        RECT 4.000 18.040 186.000 20.040 ;
        RECT 4.400 16.640 186.000 18.040 ;
        RECT 4.000 11.240 186.000 16.640 ;
        RECT 4.000 9.840 185.600 11.240 ;
        RECT 4.000 7.840 186.000 9.840 ;
        RECT 4.400 6.440 186.000 7.840 ;
        RECT 4.000 1.040 186.000 6.440 ;
        RECT 4.000 0.175 185.600 1.040 ;
      LAYER met4 ;
        RECT 123.575 15.815 123.905 55.585 ;
  END
END cbx_1__1_
END LIBRARY

