VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 142.840 4.000 143.440 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 196.000 29.350 199.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 1.000 64.770 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1.000 96.970 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 132.640 4.000 133.240 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 34.040 4.000 34.640 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.040 199.000 153.640 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
  PIN bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1.000 58.330 4.000 ;
    END
  END bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 196.000 125.950 199.000 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
  PIN bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.840 199.000 41.440 ;
    END
  END bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 3.440 4.000 4.040 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 199.000 177.440 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 95.240 4.000 95.840 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 196.000 132.390 199.000 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 115.640 4.000 116.240 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 196.000 61.550 199.000 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 199.000 55.040 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 1.000 142.050 4.000 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 196.000 22.910 199.000 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 196.000 180.690 199.000 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 196.000 187.130 199.000 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 27.240 4.000 27.840 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1.000 103.410 4.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 139.440 199.000 140.040 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 199.000 61.840 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 196.000 77.650 199.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1.000 196.790 4.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 196.000 164.590 199.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1.000 87.310 4.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 196.000 16.470 199.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1.000 55.110 4.000 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 78.240 4.000 78.840 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1.000 125.950 4.000 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 64.640 199.000 65.240 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.040 199.000 136.640 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1.000 174.250 4.000 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1.000 74.430 4.000 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 196.000 161.370 199.000 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 199.000 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1.000 167.810 4.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 199.000 82.240 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 196.000 39.010 199.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 199.000 119.640 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 196.000 84.090 199.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 199.000 163.840 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 20.440 4.000 21.040 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 199.000 89.040 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 156.440 4.000 157.040 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 176.840 4.000 177.440 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.840 199.000 160.440 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 199.000 7.440 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 196.000 106.630 199.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 196.000 93.750 199.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 196.000 154.930 199.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.040 199.000 187.640 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 196.000 116.290 199.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1.000 48.670 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 85.040 4.000 85.640 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 37.440 4.000 38.040 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 1.000 158.150 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 3.440 199.000 4.040 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 74.840 4.000 75.440 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 37.440 199.000 38.040 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 196.000 55.110 199.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 193.840 4.000 194.440 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.840 4.000 109.440 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1.000 80.870 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 125.840 4.000 126.440 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 196.000 171.030 199.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1.000 113.070 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1.000 148.490 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 122.440 199.000 123.040 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.840 199.000 24.440 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 196.000 138.830 199.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.840 199.000 194.440 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 199.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1.000 3.590 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1.000 26.130 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 196.000 67.990 199.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 196.000 45.450 199.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 105.440 199.000 106.040 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 199.000 72.040 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 199.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1.000 16.470 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 199.000 14.240 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 199.000 78.840 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 136.040 4.000 136.640 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 196.000 13.250 199.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1.000 183.910 4.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 102.040 4.000 102.640 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 196.000 0.370 199.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 196.000 193.570 199.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1.000 42.230 4.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 91.840 4.000 92.440 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1.000 119.510 4.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1.000 190.350 4.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 196.000 71.210 199.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1.000 151.710 4.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1.000 19.690 4.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 68.040 4.000 68.640 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 20.440 199.000 21.040 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 146.240 199.000 146.840 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.040 199.000 102.640 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1.000 164.590 4.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 119.040 4.000 119.640 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 47.640 199.000 48.240 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 159.840 4.000 160.440 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 199.000 112.840 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.040 199.000 170.640 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1.000 180.690 4.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.240 199.000 180.840 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 166.640 4.000 167.240 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 10.240 4.000 10.840 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 61.240 4.000 61.840 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1.000 129.170 4.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.440 4.000 191.040 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 196.000 48.670 199.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 196.000 122.730 199.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 149.640 4.000 150.240 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1.000 32.570 4.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1.000 10.030 4.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 44.240 4.000 44.840 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 196.000 109.850 199.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1.000 90.530 4.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 196.000 177.470 199.000 ;
    END
  END chany_top_out[9]
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 30.640 199.000 31.240 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 183.640 4.000 184.240 ;
    END
  END prog_clk
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 57.840 4.000 58.440 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1.000 35.790 4.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1.000 71.210 4.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 17.040 4.000 17.640 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.240 199.000 129.840 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1.000 109.850 4.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 196.000 148.490 199.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 196.000 142.050 199.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 196.000 6.810 199.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 196.000 32.570 199.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1.000 135.610 4.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
  PIN top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 51.040 4.000 51.640 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
  PIN top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 173.440 4.000 174.040 ;
    END
  END top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
  PIN top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 199.000 95.840 ;
    END
  END top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 0.070 10.240 196.810 188.320 ;
      LAYER met2 ;
        RECT 0.650 195.720 6.250 196.250 ;
        RECT 7.090 195.720 12.690 196.250 ;
        RECT 13.530 195.720 15.910 196.250 ;
        RECT 16.750 195.720 22.350 196.250 ;
        RECT 23.190 195.720 28.790 196.250 ;
        RECT 29.630 195.720 32.010 196.250 ;
        RECT 32.850 195.720 38.450 196.250 ;
        RECT 39.290 195.720 44.890 196.250 ;
        RECT 45.730 195.720 48.110 196.250 ;
        RECT 48.950 195.720 54.550 196.250 ;
        RECT 55.390 195.720 60.990 196.250 ;
        RECT 61.830 195.720 67.430 196.250 ;
        RECT 68.270 195.720 70.650 196.250 ;
        RECT 71.490 195.720 77.090 196.250 ;
        RECT 77.930 195.720 83.530 196.250 ;
        RECT 84.370 195.720 86.750 196.250 ;
        RECT 87.590 195.720 93.190 196.250 ;
        RECT 94.030 195.720 99.630 196.250 ;
        RECT 100.470 195.720 106.070 196.250 ;
        RECT 106.910 195.720 109.290 196.250 ;
        RECT 110.130 195.720 115.730 196.250 ;
        RECT 116.570 195.720 122.170 196.250 ;
        RECT 123.010 195.720 125.390 196.250 ;
        RECT 126.230 195.720 131.830 196.250 ;
        RECT 132.670 195.720 138.270 196.250 ;
        RECT 139.110 195.720 141.490 196.250 ;
        RECT 142.330 195.720 147.930 196.250 ;
        RECT 148.770 195.720 154.370 196.250 ;
        RECT 155.210 195.720 160.810 196.250 ;
        RECT 161.650 195.720 164.030 196.250 ;
        RECT 164.870 195.720 170.470 196.250 ;
        RECT 171.310 195.720 176.910 196.250 ;
        RECT 177.750 195.720 180.130 196.250 ;
        RECT 180.970 195.720 186.570 196.250 ;
        RECT 187.410 195.720 193.010 196.250 ;
        RECT 193.850 195.720 196.230 196.250 ;
        RECT 0.100 4.280 196.780 195.720 ;
        RECT 0.650 3.555 3.030 4.280 ;
        RECT 3.870 3.555 9.470 4.280 ;
        RECT 10.310 3.555 15.910 4.280 ;
        RECT 16.750 3.555 19.130 4.280 ;
        RECT 19.970 3.555 25.570 4.280 ;
        RECT 26.410 3.555 32.010 4.280 ;
        RECT 32.850 3.555 35.230 4.280 ;
        RECT 36.070 3.555 41.670 4.280 ;
        RECT 42.510 3.555 48.110 4.280 ;
        RECT 48.950 3.555 54.550 4.280 ;
        RECT 55.390 3.555 57.770 4.280 ;
        RECT 58.610 3.555 64.210 4.280 ;
        RECT 65.050 3.555 70.650 4.280 ;
        RECT 71.490 3.555 73.870 4.280 ;
        RECT 74.710 3.555 80.310 4.280 ;
        RECT 81.150 3.555 86.750 4.280 ;
        RECT 87.590 3.555 89.970 4.280 ;
        RECT 90.810 3.555 96.410 4.280 ;
        RECT 97.250 3.555 102.850 4.280 ;
        RECT 103.690 3.555 109.290 4.280 ;
        RECT 110.130 3.555 112.510 4.280 ;
        RECT 113.350 3.555 118.950 4.280 ;
        RECT 119.790 3.555 125.390 4.280 ;
        RECT 126.230 3.555 128.610 4.280 ;
        RECT 129.450 3.555 135.050 4.280 ;
        RECT 135.890 3.555 141.490 4.280 ;
        RECT 142.330 3.555 147.930 4.280 ;
        RECT 148.770 3.555 151.150 4.280 ;
        RECT 151.990 3.555 157.590 4.280 ;
        RECT 158.430 3.555 164.030 4.280 ;
        RECT 164.870 3.555 167.250 4.280 ;
        RECT 168.090 3.555 173.690 4.280 ;
        RECT 174.530 3.555 180.130 4.280 ;
        RECT 180.970 3.555 183.350 4.280 ;
        RECT 184.190 3.555 189.790 4.280 ;
        RECT 190.630 3.555 196.230 4.280 ;
      LAYER met3 ;
        RECT 4.400 193.440 195.600 194.305 ;
        RECT 4.000 191.440 196.000 193.440 ;
        RECT 4.400 190.040 196.000 191.440 ;
        RECT 4.000 188.040 196.000 190.040 ;
        RECT 4.000 186.640 195.600 188.040 ;
        RECT 4.000 184.640 196.000 186.640 ;
        RECT 4.400 183.240 196.000 184.640 ;
        RECT 4.000 181.240 196.000 183.240 ;
        RECT 4.000 179.840 195.600 181.240 ;
        RECT 4.000 177.840 196.000 179.840 ;
        RECT 4.400 176.440 195.600 177.840 ;
        RECT 4.000 174.440 196.000 176.440 ;
        RECT 4.400 173.040 196.000 174.440 ;
        RECT 4.000 171.040 196.000 173.040 ;
        RECT 4.000 169.640 195.600 171.040 ;
        RECT 4.000 167.640 196.000 169.640 ;
        RECT 4.400 166.240 196.000 167.640 ;
        RECT 4.000 164.240 196.000 166.240 ;
        RECT 4.000 162.840 195.600 164.240 ;
        RECT 4.000 160.840 196.000 162.840 ;
        RECT 4.400 159.440 195.600 160.840 ;
        RECT 4.000 157.440 196.000 159.440 ;
        RECT 4.400 156.040 196.000 157.440 ;
        RECT 4.000 154.040 196.000 156.040 ;
        RECT 4.000 152.640 195.600 154.040 ;
        RECT 4.000 150.640 196.000 152.640 ;
        RECT 4.400 149.240 196.000 150.640 ;
        RECT 4.000 147.240 196.000 149.240 ;
        RECT 4.000 145.840 195.600 147.240 ;
        RECT 4.000 143.840 196.000 145.840 ;
        RECT 4.400 142.440 196.000 143.840 ;
        RECT 4.000 140.440 196.000 142.440 ;
        RECT 4.000 139.040 195.600 140.440 ;
        RECT 4.000 137.040 196.000 139.040 ;
        RECT 4.400 135.640 195.600 137.040 ;
        RECT 4.000 133.640 196.000 135.640 ;
        RECT 4.400 132.240 196.000 133.640 ;
        RECT 4.000 130.240 196.000 132.240 ;
        RECT 4.000 128.840 195.600 130.240 ;
        RECT 4.000 126.840 196.000 128.840 ;
        RECT 4.400 125.440 196.000 126.840 ;
        RECT 4.000 123.440 196.000 125.440 ;
        RECT 4.000 122.040 195.600 123.440 ;
        RECT 4.000 120.040 196.000 122.040 ;
        RECT 4.400 118.640 195.600 120.040 ;
        RECT 4.000 116.640 196.000 118.640 ;
        RECT 4.400 115.240 196.000 116.640 ;
        RECT 4.000 113.240 196.000 115.240 ;
        RECT 4.000 111.840 195.600 113.240 ;
        RECT 4.000 109.840 196.000 111.840 ;
        RECT 4.400 108.440 196.000 109.840 ;
        RECT 4.000 106.440 196.000 108.440 ;
        RECT 4.000 105.040 195.600 106.440 ;
        RECT 4.000 103.040 196.000 105.040 ;
        RECT 4.400 101.640 195.600 103.040 ;
        RECT 4.000 96.240 196.000 101.640 ;
        RECT 4.400 94.840 195.600 96.240 ;
        RECT 4.000 92.840 196.000 94.840 ;
        RECT 4.400 91.440 196.000 92.840 ;
        RECT 4.000 89.440 196.000 91.440 ;
        RECT 4.000 88.040 195.600 89.440 ;
        RECT 4.000 86.040 196.000 88.040 ;
        RECT 4.400 84.640 196.000 86.040 ;
        RECT 4.000 82.640 196.000 84.640 ;
        RECT 4.000 81.240 195.600 82.640 ;
        RECT 4.000 79.240 196.000 81.240 ;
        RECT 4.400 77.840 195.600 79.240 ;
        RECT 4.000 75.840 196.000 77.840 ;
        RECT 4.400 74.440 196.000 75.840 ;
        RECT 4.000 72.440 196.000 74.440 ;
        RECT 4.000 71.040 195.600 72.440 ;
        RECT 4.000 69.040 196.000 71.040 ;
        RECT 4.400 67.640 196.000 69.040 ;
        RECT 4.000 65.640 196.000 67.640 ;
        RECT 4.000 64.240 195.600 65.640 ;
        RECT 4.000 62.240 196.000 64.240 ;
        RECT 4.400 60.840 195.600 62.240 ;
        RECT 4.000 58.840 196.000 60.840 ;
        RECT 4.400 57.440 196.000 58.840 ;
        RECT 4.000 55.440 196.000 57.440 ;
        RECT 4.000 54.040 195.600 55.440 ;
        RECT 4.000 52.040 196.000 54.040 ;
        RECT 4.400 50.640 196.000 52.040 ;
        RECT 4.000 48.640 196.000 50.640 ;
        RECT 4.000 47.240 195.600 48.640 ;
        RECT 4.000 45.240 196.000 47.240 ;
        RECT 4.400 43.840 196.000 45.240 ;
        RECT 4.000 41.840 196.000 43.840 ;
        RECT 4.000 40.440 195.600 41.840 ;
        RECT 4.000 38.440 196.000 40.440 ;
        RECT 4.400 37.040 195.600 38.440 ;
        RECT 4.000 35.040 196.000 37.040 ;
        RECT 4.400 33.640 196.000 35.040 ;
        RECT 4.000 31.640 196.000 33.640 ;
        RECT 4.000 30.240 195.600 31.640 ;
        RECT 4.000 28.240 196.000 30.240 ;
        RECT 4.400 26.840 196.000 28.240 ;
        RECT 4.000 24.840 196.000 26.840 ;
        RECT 4.000 23.440 195.600 24.840 ;
        RECT 4.000 21.440 196.000 23.440 ;
        RECT 4.400 20.040 195.600 21.440 ;
        RECT 4.000 18.040 196.000 20.040 ;
        RECT 4.400 16.640 196.000 18.040 ;
        RECT 4.000 14.640 196.000 16.640 ;
        RECT 4.000 13.240 195.600 14.640 ;
        RECT 4.000 11.240 196.000 13.240 ;
        RECT 4.400 9.840 196.000 11.240 ;
        RECT 4.000 7.840 196.000 9.840 ;
        RECT 4.000 6.440 195.600 7.840 ;
        RECT 4.000 4.440 196.000 6.440 ;
        RECT 4.400 3.575 195.600 4.440 ;
      LAYER met4 ;
        RECT 9.495 15.815 20.640 186.825 ;
        RECT 23.040 15.815 97.440 186.825 ;
        RECT 99.840 15.815 103.665 186.825 ;
  END
END sb_0__1_
END LIBRARY

