magic
tech sky130A
magscale 1 2
timestamp 1672422469
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 1640 39362 37584
<< metal2 >>
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 4526 39200 4582 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28354 39200 28410 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21914 200 21970 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
rect 39302 200 39358 800
<< obsm2 >>
rect 20 39144 1250 39545
rect 1418 39144 2538 39545
rect 2706 39144 4470 39545
rect 4638 39144 6402 39545
rect 6570 39144 7690 39545
rect 7858 39144 9622 39545
rect 9790 39144 11554 39545
rect 11722 39144 12842 39545
rect 13010 39144 14774 39545
rect 14942 39144 16706 39545
rect 16874 39144 17994 39545
rect 18162 39144 19926 39545
rect 20094 39144 21858 39545
rect 22026 39144 23146 39545
rect 23314 39144 25078 39545
rect 25246 39144 27010 39545
rect 27178 39144 28298 39545
rect 28466 39144 30230 39545
rect 30398 39144 32162 39545
rect 32330 39144 33450 39545
rect 33618 39144 35382 39545
rect 35550 39144 37314 39545
rect 37482 39144 38602 39545
rect 38770 39144 39356 39545
rect 20 856 39356 39144
rect 130 800 1250 856
rect 1418 800 3182 856
rect 3350 800 4470 856
rect 4638 800 6402 856
rect 6570 800 8334 856
rect 8502 800 9622 856
rect 9790 800 11554 856
rect 11722 800 13486 856
rect 13654 800 14774 856
rect 14942 800 16706 856
rect 16874 800 18638 856
rect 18806 800 19926 856
rect 20094 800 21858 856
rect 22026 800 23790 856
rect 23958 800 25078 856
rect 25246 800 27010 856
rect 27178 800 28942 856
rect 29110 800 30230 856
rect 30398 800 32162 856
rect 32330 800 34094 856
rect 34262 800 35382 856
rect 35550 800 37314 856
rect 37482 800 39246 856
<< metal3 >>
rect 200 39448 800 39568
rect 39200 38768 39800 38888
rect 200 37408 800 37528
rect 39200 37408 39800 37528
rect 200 36048 800 36168
rect 39200 35368 39800 35488
rect 200 34008 800 34128
rect 39200 33328 39800 33448
rect 200 31968 800 32088
rect 39200 31968 39800 32088
rect 200 30608 800 30728
rect 39200 29928 39800 30048
rect 200 28568 800 28688
rect 39200 27888 39800 28008
rect 200 26528 800 26648
rect 39200 26528 39800 26648
rect 200 25168 800 25288
rect 39200 24488 39800 24608
rect 200 23128 800 23248
rect 39200 22448 39800 22568
rect 200 21088 800 21208
rect 39200 21088 39800 21208
rect 200 19728 800 19848
rect 39200 19048 39800 19168
rect 200 17688 800 17808
rect 39200 17008 39800 17128
rect 200 15648 800 15768
rect 39200 15648 39800 15768
rect 200 14288 800 14408
rect 39200 13608 39800 13728
rect 200 12248 800 12368
rect 39200 11568 39800 11688
rect 200 10208 800 10328
rect 39200 10208 39800 10328
rect 200 8848 800 8968
rect 39200 8168 39800 8288
rect 200 6808 800 6928
rect 39200 6128 39800 6248
rect 200 4768 800 4888
rect 39200 4768 39800 4888
rect 200 3408 800 3528
rect 39200 2728 39800 2848
rect 200 1368 800 1488
rect 39200 688 39800 808
<< obsm3 >>
rect 880 39368 39314 39541
rect 800 38968 39314 39368
rect 800 38688 39120 38968
rect 800 37608 39314 38688
rect 880 37328 39120 37608
rect 800 36248 39314 37328
rect 880 35968 39314 36248
rect 800 35568 39314 35968
rect 800 35288 39120 35568
rect 800 34208 39314 35288
rect 880 33928 39314 34208
rect 800 33528 39314 33928
rect 800 33248 39120 33528
rect 800 32168 39314 33248
rect 880 31888 39120 32168
rect 800 30808 39314 31888
rect 880 30528 39314 30808
rect 800 30128 39314 30528
rect 800 29848 39120 30128
rect 800 28768 39314 29848
rect 880 28488 39314 28768
rect 800 28088 39314 28488
rect 800 27808 39120 28088
rect 800 26728 39314 27808
rect 880 26448 39120 26728
rect 800 25368 39314 26448
rect 880 25088 39314 25368
rect 800 24688 39314 25088
rect 800 24408 39120 24688
rect 800 23328 39314 24408
rect 880 23048 39314 23328
rect 800 22648 39314 23048
rect 800 22368 39120 22648
rect 800 21288 39314 22368
rect 880 21008 39120 21288
rect 800 19928 39314 21008
rect 880 19648 39314 19928
rect 800 19248 39314 19648
rect 800 18968 39120 19248
rect 800 17888 39314 18968
rect 880 17608 39314 17888
rect 800 17208 39314 17608
rect 800 16928 39120 17208
rect 800 15848 39314 16928
rect 880 15568 39120 15848
rect 800 14488 39314 15568
rect 880 14208 39314 14488
rect 800 13808 39314 14208
rect 800 13528 39120 13808
rect 800 12448 39314 13528
rect 880 12168 39314 12448
rect 800 11768 39314 12168
rect 800 11488 39120 11768
rect 800 10408 39314 11488
rect 880 10128 39120 10408
rect 800 9048 39314 10128
rect 880 8768 39314 9048
rect 800 8368 39314 8768
rect 800 8088 39120 8368
rect 800 7008 39314 8088
rect 880 6728 39314 7008
rect 800 6328 39314 6728
rect 800 6048 39120 6328
rect 800 4968 39314 6048
rect 880 4688 39120 4968
rect 800 3608 39314 4688
rect 880 3328 39314 3608
rect 800 2928 39314 3328
rect 800 2648 39120 2928
rect 800 1568 39314 2648
rect 880 1288 39314 1568
rect 800 888 39314 1288
rect 800 718 39120 888
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 16619 2483 19488 17645
rect 19968 2483 23309 17645
<< labels >>
rlabel metal3 s 200 3408 800 3528 6 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
port 1 nsew signal output
rlabel metal2 s 37370 39200 37426 39800 6 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
port 2 nsew signal output
rlabel metal3 s 200 17688 800 17808 6 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
port 3 nsew signal output
rlabel metal2 s 35438 200 35494 800 6 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
port 4 nsew signal output
rlabel metal2 s 14830 39200 14886 39800 6 bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
port 5 nsew signal output
rlabel metal2 s 16762 39200 16818 39800 6 bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
port 6 nsew signal output
rlabel metal2 s 18050 39200 18106 39800 6 bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_
port 7 nsew signal output
rlabel metal2 s 14830 200 14886 800 6 bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
port 8 nsew signal output
rlabel metal3 s 39200 8168 39800 8288 6 ccff_head
port 9 nsew signal input
rlabel metal2 s 35438 39200 35494 39800 6 ccff_tail
port 10 nsew signal output
rlabel metal2 s 21914 39200 21970 39800 6 chanx_left_in[0]
port 11 nsew signal input
rlabel metal2 s 13542 200 13598 800 6 chanx_left_in[10]
port 12 nsew signal input
rlabel metal3 s 39200 11568 39800 11688 6 chanx_left_in[11]
port 13 nsew signal input
rlabel metal3 s 39200 17008 39800 17128 6 chanx_left_in[12]
port 14 nsew signal input
rlabel metal3 s 39200 35368 39800 35488 6 chanx_left_in[13]
port 15 nsew signal input
rlabel metal3 s 39200 31968 39800 32088 6 chanx_left_in[14]
port 16 nsew signal input
rlabel metal3 s 39200 4768 39800 4888 6 chanx_left_in[15]
port 17 nsew signal input
rlabel metal3 s 200 28568 800 28688 6 chanx_left_in[16]
port 18 nsew signal input
rlabel metal2 s 8390 200 8446 800 6 chanx_left_in[17]
port 19 nsew signal input
rlabel metal3 s 39200 26528 39800 26648 6 chanx_left_in[18]
port 20 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 chanx_left_in[1]
port 21 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 chanx_left_in[2]
port 22 nsew signal input
rlabel metal3 s 39200 27888 39800 28008 6 chanx_left_in[3]
port 23 nsew signal input
rlabel metal2 s 37370 200 37426 800 6 chanx_left_in[4]
port 24 nsew signal input
rlabel metal2 s 25134 39200 25190 39800 6 chanx_left_in[5]
port 25 nsew signal input
rlabel metal2 s 1306 39200 1362 39800 6 chanx_left_in[6]
port 26 nsew signal input
rlabel metal3 s 39200 29928 39800 30048 6 chanx_left_in[7]
port 27 nsew signal input
rlabel metal3 s 200 19728 800 19848 6 chanx_left_in[8]
port 28 nsew signal input
rlabel metal3 s 200 23128 800 23248 6 chanx_left_in[9]
port 29 nsew signal input
rlabel metal3 s 200 1368 800 1488 6 chanx_left_out[0]
port 30 nsew signal output
rlabel metal2 s 30286 200 30342 800 6 chanx_left_out[10]
port 31 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 chanx_left_out[11]
port 32 nsew signal output
rlabel metal2 s 27066 39200 27122 39800 6 chanx_left_out[12]
port 33 nsew signal output
rlabel metal2 s 28354 39200 28410 39800 6 chanx_left_out[13]
port 34 nsew signal output
rlabel metal2 s 34150 200 34206 800 6 chanx_left_out[14]
port 35 nsew signal output
rlabel metal2 s 19982 39200 20038 39800 6 chanx_left_out[15]
port 36 nsew signal output
rlabel metal3 s 39200 33328 39800 33448 6 chanx_left_out[16]
port 37 nsew signal output
rlabel metal2 s 23846 200 23902 800 6 chanx_left_out[17]
port 38 nsew signal output
rlabel metal3 s 200 21088 800 21208 6 chanx_left_out[18]
port 39 nsew signal output
rlabel metal3 s 39200 688 39800 808 6 chanx_left_out[1]
port 40 nsew signal output
rlabel metal3 s 39200 15648 39800 15768 6 chanx_left_out[2]
port 41 nsew signal output
rlabel metal3 s 200 39448 800 39568 6 chanx_left_out[3]
port 42 nsew signal output
rlabel metal3 s 200 10208 800 10328 6 chanx_left_out[4]
port 43 nsew signal output
rlabel metal3 s 200 31968 800 32088 6 chanx_left_out[5]
port 44 nsew signal output
rlabel metal3 s 200 6808 800 6928 6 chanx_left_out[6]
port 45 nsew signal output
rlabel metal3 s 39200 37408 39800 37528 6 chanx_left_out[7]
port 46 nsew signal output
rlabel metal2 s 7746 39200 7802 39800 6 chanx_left_out[8]
port 47 nsew signal output
rlabel metal2 s 3238 200 3294 800 6 chanx_left_out[9]
port 48 nsew signal output
rlabel metal2 s 9678 200 9734 800 6 chanx_right_in[0]
port 49 nsew signal input
rlabel metal2 s 32218 200 32274 800 6 chanx_right_in[10]
port 50 nsew signal input
rlabel metal3 s 39200 13608 39800 13728 6 chanx_right_in[11]
port 51 nsew signal input
rlabel metal3 s 39200 6128 39800 6248 6 chanx_right_in[12]
port 52 nsew signal input
rlabel metal2 s 25134 200 25190 800 6 chanx_right_in[13]
port 53 nsew signal input
rlabel metal3 s 200 37408 800 37528 6 chanx_right_in[14]
port 54 nsew signal input
rlabel metal2 s 39302 200 39358 800 6 chanx_right_in[15]
port 55 nsew signal input
rlabel metal3 s 200 8848 800 8968 6 chanx_right_in[16]
port 56 nsew signal input
rlabel metal3 s 39200 10208 39800 10328 6 chanx_right_in[17]
port 57 nsew signal input
rlabel metal3 s 200 25168 800 25288 6 chanx_right_in[18]
port 58 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 chanx_right_in[1]
port 59 nsew signal input
rlabel metal3 s 39200 24488 39800 24608 6 chanx_right_in[2]
port 60 nsew signal input
rlabel metal2 s 11610 39200 11666 39800 6 chanx_right_in[3]
port 61 nsew signal input
rlabel metal2 s 6458 39200 6514 39800 6 chanx_right_in[4]
port 62 nsew signal input
rlabel metal2 s 18694 200 18750 800 6 chanx_right_in[5]
port 63 nsew signal input
rlabel metal2 s 18 200 74 800 6 chanx_right_in[6]
port 64 nsew signal input
rlabel metal2 s 21914 200 21970 800 6 chanx_right_in[7]
port 65 nsew signal input
rlabel metal2 s 12898 39200 12954 39800 6 chanx_right_in[8]
port 66 nsew signal input
rlabel metal2 s 23202 39200 23258 39800 6 chanx_right_in[9]
port 67 nsew signal input
rlabel metal2 s 33506 39200 33562 39800 6 chanx_right_out[0]
port 68 nsew signal output
rlabel metal3 s 200 26528 800 26648 6 chanx_right_out[10]
port 69 nsew signal output
rlabel metal2 s 4526 200 4582 800 6 chanx_right_out[11]
port 70 nsew signal output
rlabel metal2 s 1306 200 1362 800 6 chanx_right_out[12]
port 71 nsew signal output
rlabel metal2 s 38658 39200 38714 39800 6 chanx_right_out[13]
port 72 nsew signal output
rlabel metal2 s 30286 39200 30342 39800 6 chanx_right_out[14]
port 73 nsew signal output
rlabel metal2 s 16762 200 16818 800 6 chanx_right_out[15]
port 74 nsew signal output
rlabel metal3 s 39200 38768 39800 38888 6 chanx_right_out[16]
port 75 nsew signal output
rlabel metal3 s 39200 2728 39800 2848 6 chanx_right_out[17]
port 76 nsew signal output
rlabel metal2 s 4526 39200 4582 39800 6 chanx_right_out[18]
port 77 nsew signal output
rlabel metal3 s 39200 21088 39800 21208 6 chanx_right_out[1]
port 78 nsew signal output
rlabel metal2 s 6458 200 6514 800 6 chanx_right_out[2]
port 79 nsew signal output
rlabel metal2 s 11610 200 11666 800 6 chanx_right_out[3]
port 80 nsew signal output
rlabel metal3 s 200 15648 800 15768 6 chanx_right_out[4]
port 81 nsew signal output
rlabel metal3 s 39200 22448 39800 22568 6 chanx_right_out[5]
port 82 nsew signal output
rlabel metal2 s 19982 200 20038 800 6 chanx_right_out[6]
port 83 nsew signal output
rlabel metal3 s 200 4768 800 4888 6 chanx_right_out[7]
port 84 nsew signal output
rlabel metal2 s 32218 39200 32274 39800 6 chanx_right_out[8]
port 85 nsew signal output
rlabel metal2 s 2594 39200 2650 39800 6 chanx_right_out[9]
port 86 nsew signal output
rlabel metal2 s 9678 39200 9734 39800 6 pReset
port 87 nsew signal input
rlabel metal2 s 27066 200 27122 800 6 prog_clk
port 88 nsew signal input
rlabel metal3 s 200 12248 800 12368 6 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 89 nsew signal output
rlabel metal3 s 200 36048 800 36168 6 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 90 nsew signal output
rlabel metal3 s 39200 19048 39800 19168 6 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 91 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 93 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1898036
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/cbx_1__0_/runs/22_12_30_11_47/results/signoff/cbx_1__0_.magic.gds
string GDS_START 139574
<< end >>

