magic
tech sky130A
magscale 1 2
timestamp 1672416611
<< viali >>
rect 17693 37417 17727 37451
rect 18153 37349 18187 37383
rect 9321 37281 9355 37315
rect 12449 37281 12483 37315
rect 14473 37281 14507 37315
rect 14933 37281 14967 37315
rect 16313 37281 16347 37315
rect 17141 37281 17175 37315
rect 20821 37281 20855 37315
rect 21465 37281 21499 37315
rect 22017 37281 22051 37315
rect 35081 37281 35115 37315
rect 35541 37281 35575 37315
rect 38301 37281 38335 37315
rect 1869 37213 1903 37247
rect 2973 37213 3007 37247
rect 4905 37213 4939 37247
rect 6837 37213 6871 37247
rect 7389 37213 7423 37247
rect 7941 37213 7975 37247
rect 9873 37213 9907 37247
rect 11989 37213 12023 37247
rect 13277 37213 13311 37247
rect 15209 37213 15243 37247
rect 16957 37213 16991 37247
rect 18337 37213 18371 37247
rect 20361 37213 20395 37247
rect 22293 37213 22327 37247
rect 23305 37213 23339 37247
rect 25237 37213 25271 37247
rect 27169 37213 27203 37247
rect 27997 37213 28031 37247
rect 28457 37213 28491 37247
rect 30389 37213 30423 37247
rect 32597 37213 32631 37247
rect 33609 37213 33643 37247
rect 35817 37213 35851 37247
rect 38025 37213 38059 37247
rect 1685 37077 1719 37111
rect 2789 37077 2823 37111
rect 4721 37077 4755 37111
rect 5457 37077 5491 37111
rect 6653 37077 6687 37111
rect 8033 37077 8067 37111
rect 9965 37077 9999 37111
rect 11805 37077 11839 37111
rect 13093 37077 13127 37111
rect 20177 37077 20211 37111
rect 23489 37077 23523 37111
rect 25421 37077 25455 37111
rect 27353 37077 27387 37111
rect 28641 37077 28675 37111
rect 30573 37077 30607 37111
rect 32413 37077 32447 37111
rect 33793 37077 33827 37111
rect 22569 36873 22603 36907
rect 27905 36873 27939 36907
rect 37657 36873 37691 36907
rect 38301 36873 38335 36907
rect 2421 36805 2455 36839
rect 1685 36737 1719 36771
rect 3065 36737 3099 36771
rect 10701 36737 10735 36771
rect 22385 36737 22419 36771
rect 27721 36737 27755 36771
rect 37473 36737 37507 36771
rect 1869 36601 1903 36635
rect 2605 36601 2639 36635
rect 10517 36533 10551 36567
rect 13369 36533 13403 36567
rect 23121 36533 23155 36567
rect 36829 36533 36863 36567
rect 2421 36329 2455 36363
rect 37473 36329 37507 36363
rect 38209 36329 38243 36363
rect 1869 36125 1903 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 1685 35989 1719 36023
rect 36737 35989 36771 36023
rect 36921 35581 36955 35615
rect 37473 35581 37507 35615
rect 37749 35581 37783 35615
rect 21649 35241 21683 35275
rect 29929 35241 29963 35275
rect 38025 35241 38059 35275
rect 21465 35037 21499 35071
rect 22109 35037 22143 35071
rect 29745 35037 29779 35071
rect 30389 35037 30423 35071
rect 37841 35037 37875 35071
rect 2421 34697 2455 34731
rect 1869 34561 1903 34595
rect 2513 34561 2547 34595
rect 3065 34493 3099 34527
rect 1685 34357 1719 34391
rect 2053 33813 2087 33847
rect 38025 33473 38059 33507
rect 38209 33337 38243 33371
rect 37473 33269 37507 33303
rect 32597 32521 32631 32555
rect 1685 32385 1719 32419
rect 32689 32385 32723 32419
rect 33149 32385 33183 32419
rect 38025 32317 38059 32351
rect 38301 32317 38335 32351
rect 1777 32181 1811 32215
rect 1593 31977 1627 32011
rect 38301 31977 38335 32011
rect 1685 30617 1719 30651
rect 1869 30617 1903 30651
rect 1685 30345 1719 30379
rect 11897 30209 11931 30243
rect 38025 30209 38059 30243
rect 11805 30073 11839 30107
rect 12449 30005 12483 30039
rect 38209 30005 38243 30039
rect 22385 29801 22419 29835
rect 38025 29801 38059 29835
rect 37841 29597 37875 29631
rect 20085 29529 20119 29563
rect 20637 29529 20671 29563
rect 20821 29529 20855 29563
rect 1685 29121 1719 29155
rect 22201 29121 22235 29155
rect 22661 29121 22695 29155
rect 1869 28985 1903 29019
rect 22109 28985 22143 29019
rect 22753 28985 22787 29019
rect 21189 28713 21223 28747
rect 1593 28645 1627 28679
rect 21281 28441 21315 28475
rect 21925 28373 21959 28407
rect 15945 28033 15979 28067
rect 38025 28033 38059 28067
rect 38209 27897 38243 27931
rect 16037 27829 16071 27863
rect 37473 27829 37507 27863
rect 30757 27421 30791 27455
rect 30665 27285 30699 27319
rect 19625 27081 19659 27115
rect 38025 27013 38059 27047
rect 1869 26945 1903 26979
rect 19441 26945 19475 26979
rect 20085 26945 20119 26979
rect 37565 26945 37599 26979
rect 38209 26945 38243 26979
rect 1685 26741 1719 26775
rect 1777 25993 1811 26027
rect 1961 25857 1995 25891
rect 2421 25857 2455 25891
rect 21189 25449 21223 25483
rect 28365 25449 28399 25483
rect 1593 25245 1627 25279
rect 1869 25245 1903 25279
rect 20729 25245 20763 25279
rect 27813 25245 27847 25279
rect 32137 25245 32171 25279
rect 20637 25109 20671 25143
rect 27721 25109 27755 25143
rect 32045 25109 32079 25143
rect 1593 24905 1627 24939
rect 25789 24769 25823 24803
rect 38025 24769 38059 24803
rect 25973 24633 26007 24667
rect 26525 24565 26559 24599
rect 38209 24565 38243 24599
rect 1869 23681 1903 23715
rect 1685 23477 1719 23511
rect 20269 22729 20303 22763
rect 19625 22593 19659 22627
rect 38025 22593 38059 22627
rect 38209 22457 38243 22491
rect 19717 22389 19751 22423
rect 20729 21641 20763 21675
rect 1869 21505 1903 21539
rect 21189 21505 21223 21539
rect 38025 21505 38059 21539
rect 1685 21301 1719 21335
rect 21281 21301 21315 21335
rect 37473 21301 37507 21335
rect 38209 21301 38243 21335
rect 1777 21097 1811 21131
rect 7113 21097 7147 21131
rect 1961 20893 1995 20927
rect 7297 20893 7331 20927
rect 28641 20893 28675 20927
rect 7849 20757 7883 20791
rect 28089 20757 28123 20791
rect 28825 20757 28859 20791
rect 23581 20553 23615 20587
rect 22017 20417 22051 20451
rect 22937 20417 22971 20451
rect 25237 20417 25271 20451
rect 25881 20349 25915 20383
rect 23029 20281 23063 20315
rect 25329 20281 25363 20315
rect 19809 20213 19843 20247
rect 22109 20213 22143 20247
rect 24501 20213 24535 20247
rect 25789 20009 25823 20043
rect 22017 19873 22051 19907
rect 1869 19805 1903 19839
rect 21097 19805 21131 19839
rect 24961 19805 24995 19839
rect 25605 19805 25639 19839
rect 22109 19737 22143 19771
rect 22661 19737 22695 19771
rect 1685 19669 1719 19703
rect 19625 19669 19659 19703
rect 20269 19669 20303 19703
rect 21005 19669 21039 19703
rect 23213 19669 23247 19703
rect 24041 19669 24075 19703
rect 24869 19669 24903 19703
rect 20177 19465 20211 19499
rect 34069 19465 34103 19499
rect 18889 19397 18923 19431
rect 18981 19397 19015 19431
rect 20821 19397 20855 19431
rect 22385 19397 22419 19431
rect 22477 19397 22511 19431
rect 23949 19397 23983 19431
rect 24869 19397 24903 19431
rect 26065 19397 26099 19431
rect 26157 19397 26191 19431
rect 19993 19329 20027 19363
rect 33977 19329 34011 19363
rect 38025 19329 38059 19363
rect 20729 19261 20763 19295
rect 21005 19261 21039 19295
rect 23029 19261 23063 19295
rect 24961 19261 24995 19295
rect 25513 19261 25547 19295
rect 19441 19193 19475 19227
rect 38209 19125 38243 19159
rect 4721 18921 4755 18955
rect 19625 18921 19659 18955
rect 21465 18921 21499 18955
rect 26801 18853 26835 18887
rect 20269 18785 20303 18819
rect 22109 18785 22143 18819
rect 22385 18785 22419 18819
rect 23949 18785 23983 18819
rect 26249 18785 26283 18819
rect 4905 18717 4939 18751
rect 18245 18717 18279 18751
rect 18705 18717 18739 18751
rect 19533 18717 19567 18751
rect 21373 18717 21407 18751
rect 23397 18717 23431 18751
rect 23857 18717 23891 18751
rect 20361 18649 20395 18683
rect 20913 18649 20947 18683
rect 22201 18649 22235 18683
rect 24593 18649 24627 18683
rect 25513 18649 25547 18683
rect 25605 18649 25639 18683
rect 26341 18649 26375 18683
rect 5457 18581 5491 18615
rect 18797 18581 18831 18615
rect 23305 18581 23339 18615
rect 27353 18581 27387 18615
rect 15853 18377 15887 18411
rect 18981 18377 19015 18411
rect 20729 18377 20763 18411
rect 22109 18377 22143 18411
rect 37565 18377 37599 18411
rect 1869 18309 1903 18343
rect 19625 18309 19659 18343
rect 22845 18309 22879 18343
rect 23765 18309 23799 18343
rect 25605 18309 25639 18343
rect 25697 18309 25731 18343
rect 27169 18309 27203 18343
rect 27721 18309 27755 18343
rect 27813 18309 27847 18343
rect 1685 18241 1719 18275
rect 9689 18241 9723 18275
rect 15209 18241 15243 18275
rect 15761 18241 15795 18275
rect 20821 18241 20855 18275
rect 21281 18241 21315 18275
rect 22017 18241 22051 18275
rect 24409 18241 24443 18275
rect 26249 18241 26283 18275
rect 37473 18241 37507 18275
rect 19533 18173 19567 18207
rect 19809 18173 19843 18207
rect 22753 18173 22787 18207
rect 25053 18173 25087 18207
rect 9781 18105 9815 18139
rect 18429 18105 18463 18139
rect 28365 18105 28399 18139
rect 21373 18037 21407 18071
rect 24317 18037 24351 18071
rect 26341 18037 26375 18071
rect 26525 17833 26559 17867
rect 1593 17765 1627 17799
rect 20269 17765 20303 17799
rect 21833 17765 21867 17799
rect 22937 17765 22971 17799
rect 25329 17765 25363 17799
rect 25881 17697 25915 17731
rect 17969 17629 18003 17663
rect 18797 17629 18831 17663
rect 19533 17629 19567 17663
rect 20177 17629 20211 17663
rect 21097 17629 21131 17663
rect 23673 17629 23707 17663
rect 24593 17629 24627 17663
rect 26617 17629 26651 17663
rect 27261 17629 27295 17663
rect 27905 17629 27939 17663
rect 28365 17629 28399 17663
rect 18061 17561 18095 17595
rect 19625 17561 19659 17595
rect 22385 17561 22419 17595
rect 22477 17561 22511 17595
rect 25789 17561 25823 17595
rect 27169 17561 27203 17595
rect 18705 17493 18739 17527
rect 21189 17493 21223 17527
rect 23581 17493 23615 17527
rect 24685 17493 24719 17527
rect 27813 17493 27847 17527
rect 28457 17493 28491 17527
rect 26341 17289 26375 17323
rect 17417 17221 17451 17255
rect 17509 17221 17543 17255
rect 18521 17221 18555 17255
rect 19073 17221 19107 17255
rect 22201 17221 22235 17255
rect 23765 17221 23799 17255
rect 24961 17221 24995 17255
rect 25053 17221 25087 17255
rect 20269 17153 20303 17187
rect 21097 17153 21131 17187
rect 25605 17153 25639 17187
rect 26433 17153 26467 17187
rect 27353 17153 27387 17187
rect 27997 17153 28031 17187
rect 29009 17153 29043 17187
rect 37565 17153 37599 17187
rect 38209 17153 38243 17187
rect 17233 17085 17267 17119
rect 18429 17085 18463 17119
rect 22109 17085 22143 17119
rect 23213 17085 23247 17119
rect 23857 17085 23891 17119
rect 27261 17085 27295 17119
rect 22661 17017 22695 17051
rect 24501 17017 24535 17051
rect 27905 17017 27939 17051
rect 38025 17017 38059 17051
rect 19809 16949 19843 16983
rect 20361 16949 20395 16983
rect 21005 16949 21039 16983
rect 25697 16949 25731 16983
rect 28549 16949 28583 16983
rect 17509 16745 17543 16779
rect 18061 16745 18095 16779
rect 22937 16677 22971 16711
rect 26433 16677 26467 16711
rect 13645 16609 13679 16643
rect 15945 16609 15979 16643
rect 20545 16609 20579 16643
rect 21189 16609 21223 16643
rect 22385 16609 22419 16643
rect 24777 16609 24811 16643
rect 25237 16609 25271 16643
rect 28365 16609 28399 16643
rect 28825 16609 28859 16643
rect 3065 16541 3099 16575
rect 13001 16541 13035 16575
rect 15301 16541 15335 16575
rect 15393 16541 15427 16575
rect 18705 16541 18739 16575
rect 18797 16541 18831 16575
rect 19809 16541 19843 16575
rect 26985 16541 27019 16575
rect 27813 16541 27847 16575
rect 13093 16473 13127 16507
rect 20637 16473 20671 16507
rect 21741 16473 21775 16507
rect 21833 16473 21867 16507
rect 23397 16473 23431 16507
rect 23489 16473 23523 16507
rect 25145 16473 25179 16507
rect 25881 16473 25915 16507
rect 25973 16473 26007 16507
rect 2881 16405 2915 16439
rect 4077 16405 4111 16439
rect 17049 16405 17083 16439
rect 19901 16405 19935 16439
rect 27077 16405 27111 16439
rect 27721 16405 27755 16439
rect 19993 16201 20027 16235
rect 15761 16133 15795 16167
rect 17233 16133 17267 16167
rect 18613 16133 18647 16167
rect 21189 16133 21223 16167
rect 22194 16133 22228 16167
rect 23765 16133 23799 16167
rect 23857 16133 23891 16167
rect 24961 16133 24995 16167
rect 26433 16133 26467 16167
rect 26525 16133 26559 16167
rect 27353 16133 27387 16167
rect 1869 16065 1903 16099
rect 18521 16065 18555 16099
rect 19257 16065 19291 16099
rect 20085 16065 20119 16099
rect 28917 16065 28951 16099
rect 37565 16065 37599 16099
rect 38209 16065 38243 16099
rect 17141 15997 17175 16031
rect 19441 15997 19475 16031
rect 21281 15997 21315 16031
rect 22109 15997 22143 16031
rect 23213 15997 23247 16031
rect 24777 15997 24811 16031
rect 25053 15997 25087 16031
rect 27261 15997 27295 16031
rect 28089 15997 28123 16031
rect 17693 15929 17727 15963
rect 20729 15929 20763 15963
rect 22661 15929 22695 15963
rect 25973 15929 26007 15963
rect 1685 15861 1719 15895
rect 16313 15861 16347 15895
rect 28825 15861 28859 15895
rect 29469 15861 29503 15895
rect 38117 15861 38151 15895
rect 10517 15657 10551 15691
rect 17141 15657 17175 15691
rect 25881 15657 25915 15691
rect 29745 15657 29779 15691
rect 15393 15589 15427 15623
rect 29101 15589 29135 15623
rect 18153 15521 18187 15555
rect 19901 15521 19935 15555
rect 20085 15521 20119 15555
rect 21005 15521 21039 15555
rect 21189 15521 21223 15555
rect 25237 15521 25271 15555
rect 10425 15453 10459 15487
rect 11069 15453 11103 15487
rect 16405 15453 16439 15487
rect 17233 15453 17267 15487
rect 18061 15453 18095 15487
rect 18889 15453 18923 15487
rect 25973 15453 26007 15487
rect 28641 15453 28675 15487
rect 15945 15385 15979 15419
rect 21741 15385 21775 15419
rect 21833 15385 21867 15419
rect 22385 15385 22419 15419
rect 23397 15385 23431 15419
rect 23489 15385 23523 15419
rect 24041 15385 24075 15419
rect 24593 15385 24627 15419
rect 25152 15385 25186 15419
rect 26985 15385 27019 15419
rect 27077 15385 27111 15419
rect 27997 15385 28031 15419
rect 14841 15317 14875 15351
rect 16497 15317 16531 15351
rect 18797 15317 18831 15351
rect 19441 15317 19475 15351
rect 20545 15317 20579 15351
rect 28549 15317 28583 15351
rect 30389 15317 30423 15351
rect 15669 15113 15703 15147
rect 22109 15113 22143 15147
rect 31217 15113 31251 15147
rect 17049 15045 17083 15079
rect 18337 15045 18371 15079
rect 19533 15045 19567 15079
rect 21281 15045 21315 15079
rect 22753 15045 22787 15079
rect 24409 15045 24443 15079
rect 24501 15045 24535 15079
rect 26433 15045 26467 15079
rect 27261 15045 27295 15079
rect 27353 15045 27387 15079
rect 14657 14977 14691 15011
rect 16313 14977 16347 15011
rect 22201 14977 22235 15011
rect 22937 14977 22971 15011
rect 25053 14977 25087 15011
rect 25237 14977 25271 15011
rect 28917 14977 28951 15011
rect 29561 14977 29595 15011
rect 30205 14977 30239 15011
rect 16957 14909 16991 14943
rect 17325 14909 17359 14943
rect 18245 14909 18279 14943
rect 19441 14909 19475 14943
rect 25881 14909 25915 14943
rect 26525 14909 26559 14943
rect 28089 14909 28123 14943
rect 14749 14841 14783 14875
rect 18797 14841 18831 14875
rect 19993 14841 20027 14875
rect 23949 14841 23983 14875
rect 29469 14841 29503 14875
rect 30113 14841 30147 14875
rect 14105 14773 14139 14807
rect 16221 14773 16255 14807
rect 20637 14773 20671 14807
rect 21189 14773 21223 14807
rect 28825 14773 28859 14807
rect 30665 14773 30699 14807
rect 13185 14569 13219 14603
rect 13737 14569 13771 14603
rect 19533 14569 19567 14603
rect 27077 14569 27111 14603
rect 29837 14569 29871 14603
rect 9229 14501 9263 14535
rect 16681 14501 16715 14535
rect 29009 14501 29043 14535
rect 18061 14433 18095 14467
rect 21465 14433 21499 14467
rect 23029 14433 23063 14467
rect 26157 14433 26191 14467
rect 27629 14433 27663 14467
rect 30481 14433 30515 14467
rect 1869 14365 1903 14399
rect 8309 14365 8343 14399
rect 15485 14365 15519 14399
rect 15945 14365 15979 14399
rect 16589 14365 16623 14399
rect 17233 14365 17267 14399
rect 17877 14365 17911 14399
rect 19625 14365 19659 14399
rect 21557 14365 21591 14399
rect 22017 14365 22051 14399
rect 24041 14365 24075 14399
rect 24777 14365 24811 14399
rect 26985 14365 27019 14399
rect 28457 14365 28491 14399
rect 29101 14365 29135 14399
rect 29929 14365 29963 14399
rect 30389 14365 30423 14399
rect 17325 14297 17359 14331
rect 18521 14297 18555 14331
rect 20269 14297 20303 14331
rect 20361 14297 20395 14331
rect 20913 14297 20947 14331
rect 23213 14297 23247 14331
rect 23305 14297 23339 14331
rect 26341 14297 26375 14331
rect 26433 14297 26467 14331
rect 31585 14297 31619 14331
rect 1685 14229 1719 14263
rect 8125 14229 8159 14263
rect 14381 14229 14415 14263
rect 15393 14229 15427 14263
rect 16037 14229 16071 14263
rect 22109 14229 22143 14263
rect 23949 14229 23983 14263
rect 24685 14229 24719 14263
rect 25237 14229 25271 14263
rect 28365 14229 28399 14263
rect 31125 14229 31159 14263
rect 15577 14025 15611 14059
rect 16221 14025 16255 14059
rect 17509 14025 17543 14059
rect 19993 14025 20027 14059
rect 30297 14025 30331 14059
rect 31493 14025 31527 14059
rect 13645 13957 13679 13991
rect 14289 13957 14323 13991
rect 18153 13957 18187 13991
rect 19073 13957 19107 13991
rect 19165 13957 19199 13991
rect 20637 13957 20671 13991
rect 20729 13957 20763 13991
rect 23949 13957 23983 13991
rect 25789 13957 25823 13991
rect 26341 13957 26375 13991
rect 27169 13957 27203 13991
rect 27721 13957 27755 13991
rect 27813 13957 27847 13991
rect 28549 13957 28583 13991
rect 14197 13889 14231 13923
rect 15485 13889 15519 13923
rect 16129 13889 16163 13923
rect 16865 13889 16899 13923
rect 17049 13889 17083 13923
rect 19901 13889 19935 13923
rect 22201 13889 22235 13923
rect 24593 13889 24627 13923
rect 25237 13889 25271 13923
rect 29745 13889 29779 13923
rect 30205 13889 30239 13923
rect 30849 13889 30883 13923
rect 12633 13821 12667 13855
rect 15025 13821 15059 13855
rect 22017 13821 22051 13855
rect 23765 13821 23799 13855
rect 24041 13821 24075 13855
rect 26433 13821 26467 13855
rect 28457 13821 28491 13855
rect 28917 13821 28951 13855
rect 29653 13821 29687 13855
rect 30941 13821 30975 13855
rect 38025 13821 38059 13855
rect 38301 13821 38335 13855
rect 13185 13753 13219 13787
rect 21189 13753 21223 13787
rect 22385 13685 22419 13719
rect 24685 13685 24719 13719
rect 10609 13481 10643 13515
rect 16957 13481 16991 13515
rect 31125 13481 31159 13515
rect 38301 13481 38335 13515
rect 13645 13413 13679 13447
rect 21741 13413 21775 13447
rect 14381 13345 14415 13379
rect 15669 13345 15703 13379
rect 19901 13345 19935 13379
rect 25329 13345 25363 13379
rect 25973 13345 26007 13379
rect 26617 13345 26651 13379
rect 27353 13345 27387 13379
rect 29837 13345 29871 13379
rect 31769 13345 31803 13379
rect 10701 13277 10735 13311
rect 15025 13277 15059 13311
rect 16313 13277 16347 13311
rect 16865 13277 16899 13311
rect 18705 13277 18739 13311
rect 27997 13277 28031 13311
rect 29193 13277 29227 13311
rect 29929 13277 29963 13311
rect 30573 13277 30607 13311
rect 31033 13277 31067 13311
rect 12081 13209 12115 13243
rect 13185 13209 13219 13243
rect 14473 13209 14507 13243
rect 15761 13209 15795 13243
rect 17601 13209 17635 13243
rect 17693 13209 17727 13243
rect 18245 13209 18279 13243
rect 20821 13209 20855 13243
rect 20913 13209 20947 13243
rect 22201 13209 22235 13243
rect 22293 13209 22327 13243
rect 22845 13209 22879 13243
rect 23397 13209 23431 13243
rect 23489 13209 23523 13243
rect 24685 13209 24719 13243
rect 24777 13209 24811 13243
rect 26525 13209 26559 13243
rect 27445 13209 27479 13243
rect 28549 13209 28583 13243
rect 28641 13209 28675 13243
rect 12633 13141 12667 13175
rect 18797 13141 18831 13175
rect 30481 13141 30515 13175
rect 32321 13141 32355 13175
rect 12449 12937 12483 12971
rect 15577 12937 15611 12971
rect 29653 12937 29687 12971
rect 30941 12937 30975 12971
rect 11897 12869 11931 12903
rect 14933 12869 14967 12903
rect 17693 12869 17727 12903
rect 18797 12869 18831 12903
rect 18889 12869 18923 12903
rect 21097 12869 21131 12903
rect 22201 12869 22235 12903
rect 23765 12869 23799 12903
rect 24593 12869 24627 12903
rect 25605 12869 25639 12903
rect 26157 12869 26191 12903
rect 27728 12869 27762 12903
rect 28457 12869 28491 12903
rect 28549 12869 28583 12903
rect 1869 12801 1903 12835
rect 12909 12801 12943 12835
rect 13553 12801 13587 12835
rect 14197 12801 14231 12835
rect 14841 12801 14875 12835
rect 15485 12801 15519 12835
rect 16129 12801 16163 12835
rect 17049 12801 17083 12835
rect 20085 12801 20119 12835
rect 20545 12801 20579 12835
rect 21005 12801 21039 12835
rect 29745 12801 29779 12835
rect 30389 12801 30423 12835
rect 31033 12801 31067 12835
rect 33241 12801 33275 12835
rect 17601 12733 17635 12767
rect 18245 12733 18279 12767
rect 19901 12733 19935 12767
rect 22109 12733 22143 12767
rect 22753 12733 22787 12767
rect 23857 12733 23891 12767
rect 24501 12733 24535 12767
rect 24777 12733 24811 12767
rect 26249 12733 26283 12767
rect 27813 12733 27847 12767
rect 28825 12733 28859 12767
rect 31493 12733 31527 12767
rect 13001 12665 13035 12699
rect 14289 12665 14323 12699
rect 19349 12665 19383 12699
rect 23305 12665 23339 12699
rect 27261 12665 27295 12699
rect 30297 12665 30331 12699
rect 1685 12597 1719 12631
rect 13645 12597 13679 12631
rect 16221 12597 16255 12631
rect 16957 12597 16991 12631
rect 33333 12597 33367 12631
rect 13093 12393 13127 12427
rect 13645 12325 13679 12359
rect 20453 12325 20487 12359
rect 22845 12325 22879 12359
rect 27077 12325 27111 12359
rect 28825 12325 28859 12359
rect 16589 12257 16623 12291
rect 18245 12257 18279 12291
rect 19901 12257 19935 12291
rect 22293 12257 22327 12291
rect 23397 12257 23431 12291
rect 25237 12257 25271 12291
rect 26433 12257 26467 12291
rect 27629 12257 27663 12291
rect 30481 12257 30515 12291
rect 12541 12189 12575 12223
rect 13553 12189 13587 12223
rect 14657 12189 14691 12223
rect 24593 12189 24627 12223
rect 29929 12189 29963 12223
rect 30389 12189 30423 12223
rect 31033 12189 31067 12223
rect 31125 12189 31159 12223
rect 15393 12121 15427 12155
rect 15485 12121 15519 12155
rect 16037 12121 16071 12155
rect 16681 12121 16715 12155
rect 17233 12121 17267 12155
rect 18337 12121 18371 12155
rect 18889 12121 18923 12155
rect 19993 12121 20027 12155
rect 21097 12121 21131 12155
rect 21189 12121 21223 12155
rect 21741 12121 21775 12155
rect 22385 12121 22419 12155
rect 25145 12121 25179 12155
rect 25789 12121 25823 12155
rect 26341 12121 26375 12155
rect 27537 12121 27571 12155
rect 28273 12121 28307 12155
rect 28365 12121 28399 12155
rect 32229 12121 32263 12155
rect 14749 12053 14783 12087
rect 29837 12053 29871 12087
rect 31677 12053 31711 12087
rect 13737 11849 13771 11883
rect 15025 11849 15059 11883
rect 24317 11849 24351 11883
rect 31585 11849 31619 11883
rect 11989 11781 12023 11815
rect 14381 11781 14415 11815
rect 15761 11781 15795 11815
rect 16313 11781 16347 11815
rect 17785 11781 17819 11815
rect 18981 11781 19015 11815
rect 21281 11781 21315 11815
rect 23489 11781 23523 11815
rect 27169 11781 27203 11815
rect 27721 11781 27755 11815
rect 28457 11781 28491 11815
rect 28549 11781 28583 11815
rect 29101 11781 29135 11815
rect 29653 11781 29687 11815
rect 13185 11713 13219 11747
rect 13645 11713 13679 11747
rect 14473 11713 14507 11747
rect 14933 11713 14967 11747
rect 17141 11713 17175 11747
rect 24409 11713 24443 11747
rect 26617 11713 26651 11747
rect 29561 11713 29595 11747
rect 30389 11713 30423 11747
rect 30941 11713 30975 11747
rect 31033 11713 31067 11747
rect 31677 11713 31711 11747
rect 37565 11713 37599 11747
rect 38209 11713 38243 11747
rect 15669 11645 15703 11679
rect 17693 11645 17727 11679
rect 18889 11645 18923 11679
rect 19441 11645 19475 11679
rect 21097 11645 21131 11679
rect 21373 11645 21407 11679
rect 23765 11645 23799 11679
rect 24869 11645 24903 11679
rect 27813 11645 27847 11679
rect 12541 11577 12575 11611
rect 18245 11577 18279 11611
rect 30297 11577 30331 11611
rect 38025 11577 38059 11611
rect 13093 11509 13127 11543
rect 17049 11509 17083 11543
rect 22017 11509 22051 11543
rect 26359 11509 26393 11543
rect 32321 11509 32355 11543
rect 12173 11305 12207 11339
rect 14381 11305 14415 11339
rect 18153 11305 18187 11339
rect 27721 11305 27755 11339
rect 29837 11305 29871 11339
rect 17325 11237 17359 11271
rect 20269 11237 20303 11271
rect 22109 11237 22143 11271
rect 24685 11237 24719 11271
rect 28365 11237 28399 11271
rect 33241 11237 33275 11271
rect 15577 11169 15611 11203
rect 15761 11169 15795 11203
rect 16773 11169 16807 11203
rect 19717 11169 19751 11203
rect 25973 11169 26007 11203
rect 12909 11101 12943 11135
rect 13553 11101 13587 11135
rect 14289 11101 14323 11135
rect 14933 11101 14967 11135
rect 18245 11101 18279 11135
rect 18889 11101 18923 11135
rect 20821 11101 20855 11135
rect 23857 11101 23891 11135
rect 29929 11101 29963 11135
rect 30389 11101 30423 11135
rect 33425 11101 33459 11135
rect 13645 11033 13679 11067
rect 15025 11033 15059 11067
rect 16865 11033 16899 11067
rect 18797 11033 18831 11067
rect 19809 11033 19843 11067
rect 21373 11033 21407 11067
rect 21465 11033 21499 11067
rect 23581 11033 23615 11067
rect 25145 11033 25179 11067
rect 25237 11033 25271 11067
rect 26249 11033 26283 11067
rect 28825 11033 28859 11067
rect 28917 11033 28951 11067
rect 31033 11033 31067 11067
rect 31585 11033 31619 11067
rect 32137 11033 32171 11067
rect 12725 10965 12759 10999
rect 16221 10965 16255 10999
rect 30481 10965 30515 10999
rect 12357 10761 12391 10795
rect 13461 10761 13495 10795
rect 16957 10761 16991 10795
rect 26525 10761 26559 10795
rect 31125 10761 31159 10795
rect 31677 10761 31711 10795
rect 32873 10761 32907 10795
rect 38117 10761 38151 10795
rect 12817 10693 12851 10727
rect 18889 10693 18923 10727
rect 20453 10693 20487 10727
rect 21281 10693 21315 10727
rect 23581 10693 23615 10727
rect 25053 10693 25087 10727
rect 32413 10693 32447 10727
rect 1685 10625 1719 10659
rect 9229 10625 9263 10659
rect 9873 10625 9907 10659
rect 14749 10625 14783 10659
rect 15853 10625 15887 10659
rect 17417 10625 17451 10659
rect 21189 10625 21223 10659
rect 23857 10625 23891 10659
rect 24777 10625 24811 10659
rect 27353 10625 27387 10659
rect 30665 10625 30699 10659
rect 37657 10625 37691 10659
rect 38301 10625 38335 10659
rect 14105 10557 14139 10591
rect 14565 10557 14599 10591
rect 15669 10557 15703 10591
rect 18245 10557 18279 10591
rect 18797 10557 18831 10591
rect 20269 10557 20303 10591
rect 20545 10557 20579 10591
rect 27997 10557 28031 10591
rect 29745 10557 29779 10591
rect 30021 10557 30055 10591
rect 9321 10489 9355 10523
rect 19349 10489 19383 10523
rect 1777 10421 1811 10455
rect 15209 10421 15243 10455
rect 16037 10421 16071 10455
rect 17509 10421 17543 10455
rect 22109 10421 22143 10455
rect 27261 10421 27295 10455
rect 30573 10421 30607 10455
rect 33425 10421 33459 10455
rect 1593 10217 1627 10251
rect 10977 10217 11011 10251
rect 20821 10217 20855 10251
rect 25421 10217 25455 10251
rect 26911 10217 26945 10251
rect 28917 10217 28951 10251
rect 31321 10217 31355 10251
rect 32045 10217 32079 10251
rect 17233 10149 17267 10183
rect 19533 10149 19567 10183
rect 33701 10149 33735 10183
rect 13185 10081 13219 10115
rect 15393 10081 15427 10115
rect 18521 10081 18555 10115
rect 23397 10081 23431 10115
rect 24041 10081 24075 10115
rect 27169 10081 27203 10115
rect 27997 10081 28031 10115
rect 28273 10081 28307 10115
rect 31585 10081 31619 10115
rect 11069 10013 11103 10047
rect 14657 10013 14691 10047
rect 15301 10013 15335 10047
rect 16129 10013 16163 10047
rect 20913 10013 20947 10047
rect 24777 10013 24811 10047
rect 29009 10013 29043 10047
rect 35357 10013 35391 10047
rect 35817 10013 35851 10047
rect 13737 9945 13771 9979
rect 16681 9945 16715 9979
rect 16773 9945 16807 9979
rect 17877 9945 17911 9979
rect 17969 9945 18003 9979
rect 19993 9945 20027 9979
rect 20085 9945 20119 9979
rect 21373 9945 21407 9979
rect 23121 9945 23155 9979
rect 28181 9945 28215 9979
rect 32689 9945 32723 9979
rect 33149 9945 33183 9979
rect 35265 9945 35299 9979
rect 14749 9877 14783 9911
rect 16037 9877 16071 9911
rect 24685 9877 24719 9911
rect 29837 9877 29871 9911
rect 15025 9673 15059 9707
rect 9413 9605 9447 9639
rect 13185 9605 13219 9639
rect 14381 9605 14415 9639
rect 15761 9605 15795 9639
rect 17141 9605 17175 9639
rect 17693 9605 17727 9639
rect 18337 9605 18371 9639
rect 22109 9605 22143 9639
rect 22661 9605 22695 9639
rect 23213 9605 23247 9639
rect 26433 9605 26467 9639
rect 27261 9605 27295 9639
rect 29653 9605 29687 9639
rect 30481 9605 30515 9639
rect 8861 9537 8895 9571
rect 12633 9537 12667 9571
rect 13645 9537 13679 9571
rect 14289 9537 14323 9571
rect 14933 9537 14967 9571
rect 22017 9537 22051 9571
rect 25881 9537 25915 9571
rect 26525 9537 26559 9571
rect 27169 9537 27203 9571
rect 32413 9537 32447 9571
rect 32505 9537 32539 9571
rect 33149 9537 33183 9571
rect 15669 9469 15703 9503
rect 15945 9469 15979 9503
rect 17049 9469 17083 9503
rect 18245 9469 18279 9503
rect 19717 9469 19751 9503
rect 19993 9469 20027 9503
rect 21465 9469 21499 9503
rect 23305 9469 23339 9503
rect 23857 9469 23891 9503
rect 25605 9469 25639 9503
rect 27905 9469 27939 9503
rect 29929 9469 29963 9503
rect 18797 9401 18831 9435
rect 34161 9401 34195 9435
rect 8677 9333 8711 9367
rect 13737 9333 13771 9367
rect 30941 9333 30975 9367
rect 31493 9333 31527 9367
rect 33057 9333 33091 9367
rect 33609 9333 33643 9367
rect 37565 9333 37599 9367
rect 38301 9333 38335 9367
rect 23673 9129 23707 9163
rect 26985 9129 27019 9163
rect 29837 9129 29871 9163
rect 32045 9129 32079 9163
rect 14841 9061 14875 9095
rect 20729 9061 20763 9095
rect 33149 9061 33183 9095
rect 1869 8993 1903 9027
rect 15485 8993 15519 9027
rect 16129 8993 16163 9027
rect 17141 8993 17175 9027
rect 18705 8993 18739 9027
rect 19809 8993 19843 9027
rect 23121 8993 23155 9027
rect 26157 8993 26191 9027
rect 28733 8993 28767 9027
rect 31585 8993 31619 9027
rect 1593 8925 1627 8959
rect 12725 8925 12759 8959
rect 14749 8925 14783 8959
rect 20821 8925 20855 8959
rect 23765 8925 23799 8959
rect 26433 8925 26467 8959
rect 36093 8925 36127 8959
rect 36553 8925 36587 8959
rect 37565 8925 37599 8959
rect 38025 8925 38059 8959
rect 12817 8857 12851 8891
rect 13737 8857 13771 8891
rect 15577 8857 15611 8891
rect 16682 8857 16716 8891
rect 16773 8857 16807 8891
rect 18245 8857 18279 8891
rect 18337 8857 18371 8891
rect 19533 8857 19567 8891
rect 19625 8857 19659 8891
rect 22845 8857 22879 8891
rect 28457 8857 28491 8891
rect 31309 8857 31343 8891
rect 32597 8857 32631 8891
rect 33793 8857 33827 8891
rect 36001 8857 36035 8891
rect 21373 8789 21407 8823
rect 24685 8789 24719 8823
rect 37473 8789 37507 8823
rect 1593 8585 1627 8619
rect 13369 8585 13403 8619
rect 15577 8585 15611 8619
rect 16221 8585 16255 8619
rect 20361 8585 20395 8619
rect 21373 8585 21407 8619
rect 22109 8585 22143 8619
rect 27261 8585 27295 8619
rect 13921 8517 13955 8551
rect 14473 8517 14507 8551
rect 17969 8517 18003 8551
rect 19625 8517 19659 8551
rect 23581 8517 23615 8551
rect 30389 8517 30423 8551
rect 15485 8449 15519 8483
rect 16129 8449 16163 8483
rect 17141 8449 17175 8483
rect 20269 8449 20303 8483
rect 23857 8449 23891 8483
rect 24317 8449 24351 8483
rect 27353 8449 27387 8483
rect 30297 8449 30331 8483
rect 37749 8449 37783 8483
rect 17877 8381 17911 8415
rect 19717 8381 19751 8415
rect 24593 8381 24627 8415
rect 26065 8381 26099 8415
rect 27813 8381 27847 8415
rect 28089 8381 28123 8415
rect 29837 8381 29871 8415
rect 31493 8381 31527 8415
rect 36921 8381 36955 8415
rect 37473 8381 37507 8415
rect 14933 8313 14967 8347
rect 17233 8313 17267 8347
rect 18429 8313 18463 8347
rect 19165 8313 19199 8347
rect 30941 8313 30975 8347
rect 32321 8313 32355 8347
rect 32873 8313 32907 8347
rect 33425 8313 33459 8347
rect 34069 8313 34103 8347
rect 36369 8313 36403 8347
rect 12725 8041 12759 8075
rect 18797 8041 18831 8075
rect 20729 8041 20763 8075
rect 21649 8041 21683 8075
rect 23949 8041 23983 8075
rect 28929 8041 28963 8075
rect 36001 8041 36035 8075
rect 13369 7973 13403 8007
rect 27445 7973 27479 8007
rect 31493 7973 31527 8007
rect 33057 7973 33091 8007
rect 37933 7973 37967 8007
rect 14381 7905 14415 7939
rect 15669 7905 15703 7939
rect 16865 7905 16899 7939
rect 17785 7905 17819 7939
rect 18153 7905 18187 7939
rect 20085 7905 20119 7939
rect 23397 7905 23431 7939
rect 26433 7905 26467 7939
rect 30021 7905 30055 7939
rect 36645 7905 36679 7939
rect 12633 7837 12667 7871
rect 13277 7837 13311 7871
rect 15025 7837 15059 7871
rect 15577 7837 15611 7871
rect 18889 7837 18923 7871
rect 20821 7837 20855 7871
rect 24041 7837 24075 7871
rect 26709 7837 26743 7871
rect 29193 7837 29227 7871
rect 29745 7837 29779 7871
rect 35449 7837 35483 7871
rect 37197 7837 37231 7871
rect 37841 7837 37875 7871
rect 14473 7769 14507 7803
rect 16221 7769 16255 7803
rect 16773 7769 16807 7803
rect 18061 7769 18095 7803
rect 19441 7769 19475 7803
rect 19993 7769 20027 7803
rect 23121 7769 23155 7803
rect 24685 7769 24719 7803
rect 35357 7769 35391 7803
rect 31953 7701 31987 7735
rect 32597 7701 32631 7735
rect 33609 7701 33643 7735
rect 37381 7701 37415 7735
rect 13645 7497 13679 7531
rect 14933 7497 14967 7531
rect 29745 7497 29779 7531
rect 35081 7497 35115 7531
rect 36277 7497 36311 7531
rect 1869 7429 1903 7463
rect 16221 7429 16255 7463
rect 16957 7429 16991 7463
rect 17049 7429 17083 7463
rect 19533 7429 19567 7463
rect 24501 7429 24535 7463
rect 28273 7429 28307 7463
rect 30205 7429 30239 7463
rect 36829 7429 36863 7463
rect 1685 7361 1719 7395
rect 12633 7361 12667 7395
rect 13553 7361 13587 7395
rect 14197 7361 14231 7395
rect 15025 7361 15059 7395
rect 15485 7361 15519 7395
rect 15577 7361 15611 7395
rect 16313 7361 16347 7395
rect 18337 7361 18371 7395
rect 24041 7361 24075 7395
rect 27169 7361 27203 7395
rect 37657 7361 37691 7395
rect 38117 7361 38151 7395
rect 12173 7293 12207 7327
rect 14289 7293 14323 7327
rect 19625 7293 19659 7327
rect 22017 7293 22051 7327
rect 23765 7293 23799 7327
rect 26249 7293 26283 7327
rect 26525 7293 26559 7327
rect 27997 7293 28031 7327
rect 31401 7293 31435 7327
rect 37565 7293 37599 7327
rect 17509 7225 17543 7259
rect 19073 7225 19107 7259
rect 27261 7225 27295 7259
rect 32413 7225 32447 7259
rect 32965 7225 32999 7259
rect 33425 7225 33459 7259
rect 34529 7225 34563 7259
rect 38209 7225 38243 7259
rect 12725 7157 12759 7191
rect 18429 7157 18463 7191
rect 20361 7157 20395 7191
rect 20913 7157 20947 7191
rect 21373 7157 21407 7191
rect 30849 7157 30883 7191
rect 33977 7157 34011 7191
rect 35725 7157 35759 7191
rect 1593 6953 1627 6987
rect 13001 6953 13035 6987
rect 30002 6953 30036 6987
rect 31493 6953 31527 6987
rect 32045 6953 32079 6987
rect 37105 6953 37139 6987
rect 37657 6953 37691 6987
rect 38209 6953 38243 6987
rect 21189 6885 21223 6919
rect 23397 6885 23431 6919
rect 12357 6817 12391 6851
rect 15853 6817 15887 6851
rect 16497 6817 16531 6851
rect 17785 6817 17819 6851
rect 19441 6817 19475 6851
rect 21649 6817 21683 6851
rect 25513 6817 25547 6851
rect 26249 6817 26283 6851
rect 32505 6817 32539 6851
rect 35449 6817 35483 6851
rect 12265 6749 12299 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 14473 6749 14507 6783
rect 15117 6749 15151 6783
rect 15209 6749 15243 6783
rect 15761 6749 15795 6783
rect 16589 6749 16623 6783
rect 17233 6749 17267 6783
rect 17877 6749 17911 6783
rect 18337 6749 18371 6783
rect 24041 6749 24075 6783
rect 24777 6749 24811 6783
rect 25421 6749 25455 6783
rect 28733 6749 28767 6783
rect 29745 6749 29779 6783
rect 13645 6681 13679 6715
rect 14565 6681 14599 6715
rect 17141 6681 17175 6715
rect 19717 6681 19751 6715
rect 21925 6681 21959 6715
rect 23949 6681 23983 6715
rect 26525 6681 26559 6715
rect 28641 6681 28675 6715
rect 34161 6681 34195 6715
rect 18521 6613 18555 6647
rect 24685 6613 24719 6647
rect 27997 6613 28031 6647
rect 33149 6613 33183 6647
rect 33609 6613 33643 6647
rect 34897 6613 34931 6647
rect 36001 6613 36035 6647
rect 36645 6613 36679 6647
rect 12449 6409 12483 6443
rect 13093 6409 13127 6443
rect 13737 6409 13771 6443
rect 15025 6409 15059 6443
rect 20269 6409 20303 6443
rect 27261 6409 27295 6443
rect 27997 6409 28031 6443
rect 33977 6409 34011 6443
rect 15761 6341 15795 6375
rect 18337 6341 18371 6375
rect 19533 6341 19567 6375
rect 19625 6341 19659 6375
rect 29469 6341 29503 6375
rect 36001 6341 36035 6375
rect 38025 6341 38059 6375
rect 12541 6273 12575 6307
rect 13185 6273 13219 6307
rect 13645 6273 13679 6307
rect 14289 6273 14323 6307
rect 14933 6273 14967 6307
rect 16313 6273 16347 6307
rect 20361 6273 20395 6307
rect 23857 6273 23891 6307
rect 27169 6273 27203 6307
rect 30389 6273 30423 6307
rect 35449 6273 35483 6307
rect 36093 6273 36127 6307
rect 36553 6273 36587 6307
rect 37565 6273 37599 6307
rect 38209 6273 38243 6307
rect 15669 6205 15703 6239
rect 17325 6205 17359 6239
rect 18429 6205 18463 6239
rect 22109 6205 22143 6239
rect 23581 6205 23615 6239
rect 24593 6205 24627 6239
rect 26341 6205 26375 6239
rect 26617 6205 26651 6239
rect 29745 6205 29779 6239
rect 30941 6205 30975 6239
rect 32413 6205 32447 6239
rect 32965 6205 32999 6239
rect 14381 6137 14415 6171
rect 17877 6137 17911 6171
rect 19073 6137 19107 6171
rect 33425 6137 33459 6171
rect 20913 6069 20947 6103
rect 21373 6069 21407 6103
rect 30297 6069 30331 6103
rect 31401 6069 31435 6103
rect 34529 6069 34563 6103
rect 35357 6069 35391 6103
rect 12265 5865 12299 5899
rect 13645 5865 13679 5899
rect 14381 5865 14415 5899
rect 15577 5865 15611 5899
rect 17049 5865 17083 5899
rect 33701 5865 33735 5899
rect 37105 5865 37139 5899
rect 38209 5865 38243 5899
rect 17601 5797 17635 5831
rect 20821 5797 20855 5831
rect 26341 5797 26375 5831
rect 28917 5797 28951 5831
rect 31493 5797 31527 5831
rect 36001 5797 36035 5831
rect 37657 5797 37691 5831
rect 18245 5729 18279 5763
rect 24593 5729 24627 5763
rect 24869 5729 24903 5763
rect 27445 5729 27479 5763
rect 29745 5729 29779 5763
rect 30021 5729 30055 5763
rect 31953 5729 31987 5763
rect 35449 5729 35483 5763
rect 11713 5661 11747 5695
rect 13553 5661 13587 5695
rect 14841 5661 14875 5695
rect 15669 5661 15703 5695
rect 16129 5661 16163 5695
rect 16949 5663 16983 5697
rect 18889 5661 18923 5695
rect 21373 5661 21407 5695
rect 24041 5661 24075 5695
rect 27169 5661 27203 5695
rect 16221 5593 16255 5627
rect 18330 5593 18364 5627
rect 19809 5593 19843 5627
rect 20269 5593 20303 5627
rect 21649 5593 21683 5627
rect 23397 5593 23431 5627
rect 32229 5593 32263 5627
rect 11529 5525 11563 5559
rect 14933 5525 14967 5559
rect 23949 5525 23983 5559
rect 34253 5525 34287 5559
rect 34897 5525 34931 5559
rect 36553 5525 36587 5559
rect 14013 5321 14047 5355
rect 15209 5321 15243 5355
rect 16957 5321 16991 5355
rect 23765 5321 23799 5355
rect 30021 5321 30055 5355
rect 34529 5321 34563 5355
rect 36093 5321 36127 5355
rect 37473 5321 37507 5355
rect 13461 5253 13495 5287
rect 16129 5253 16163 5287
rect 18429 5253 18463 5287
rect 18521 5253 18555 5287
rect 19073 5253 19107 5287
rect 20729 5253 20763 5287
rect 25789 5253 25823 5287
rect 26617 5253 26651 5287
rect 33885 5253 33919 5287
rect 38025 5253 38059 5287
rect 1869 5185 1903 5219
rect 12265 5185 12299 5219
rect 14473 5185 14507 5219
rect 15301 5185 15335 5219
rect 16037 5185 16071 5219
rect 17049 5185 17083 5219
rect 20637 5185 20671 5219
rect 21281 5185 21315 5219
rect 26065 5185 26099 5219
rect 27353 5185 27387 5219
rect 30757 5185 30791 5219
rect 32505 5185 32539 5219
rect 33425 5185 33459 5219
rect 38209 5185 38243 5219
rect 12357 5117 12391 5151
rect 22017 5117 22051 5151
rect 22293 5117 22327 5151
rect 28273 5117 28307 5151
rect 28549 5117 28583 5151
rect 30481 5117 30515 5151
rect 17969 5049 18003 5083
rect 36645 5049 36679 5083
rect 1685 4981 1719 5015
rect 14565 4981 14599 5015
rect 20177 4981 20211 5015
rect 21373 4981 21407 5015
rect 24317 4981 24351 5015
rect 27261 4981 27295 5015
rect 32597 4981 32631 5015
rect 33333 4981 33367 5015
rect 34989 4981 35023 5015
rect 35541 4981 35575 5015
rect 10333 4777 10367 4811
rect 14565 4777 14599 4811
rect 18245 4777 18279 4811
rect 31493 4777 31527 4811
rect 32505 4777 32539 4811
rect 13737 4709 13771 4743
rect 20177 4709 20211 4743
rect 20729 4709 20763 4743
rect 21189 4709 21223 4743
rect 36185 4709 36219 4743
rect 15761 4641 15795 4675
rect 16405 4641 16439 4675
rect 17049 4641 17083 4675
rect 22937 4641 22971 4675
rect 26065 4641 26099 4675
rect 28549 4641 28583 4675
rect 35541 4641 35575 4675
rect 10425 4573 10459 4607
rect 14473 4573 14507 4607
rect 15677 4567 15711 4601
rect 18337 4573 18371 4607
rect 18889 4573 18923 4607
rect 24041 4573 24075 4607
rect 26341 4573 26375 4607
rect 28825 4573 28859 4607
rect 29745 4573 29779 4607
rect 32321 4573 32355 4607
rect 34253 4573 34287 4607
rect 35633 4573 35667 4607
rect 36277 4573 36311 4607
rect 37841 4573 37875 4607
rect 17118 4505 17152 4539
rect 17693 4505 17727 4539
rect 22661 4505 22695 4539
rect 30021 4505 30055 4539
rect 33057 4505 33091 4539
rect 33609 4505 33643 4539
rect 36737 4505 36771 4539
rect 15209 4437 15243 4471
rect 19533 4437 19567 4471
rect 23949 4437 23983 4471
rect 24593 4437 24627 4471
rect 27077 4437 27111 4471
rect 34161 4437 34195 4471
rect 34897 4437 34931 4471
rect 37749 4437 37783 4471
rect 22201 4233 22235 4267
rect 33425 4233 33459 4267
rect 14657 4165 14691 4199
rect 17601 4165 17635 4199
rect 24409 4165 24443 4199
rect 26617 4165 26651 4199
rect 13461 4097 13495 4131
rect 14013 4097 14047 4131
rect 14933 4097 14967 4131
rect 15485 4097 15519 4131
rect 16313 4097 16347 4131
rect 17233 4097 17267 4131
rect 18245 4097 18279 4131
rect 18337 4097 18371 4131
rect 18981 4097 19015 4131
rect 22017 4097 22051 4131
rect 25789 4097 25823 4131
rect 28917 4097 28951 4131
rect 31585 4097 31619 4131
rect 32689 4097 32723 4131
rect 36921 4097 36955 4131
rect 37749 4097 37783 4131
rect 15577 4029 15611 4063
rect 24685 4029 24719 4063
rect 26065 4029 26099 4063
rect 27169 4029 27203 4063
rect 29377 4029 29411 4063
rect 31125 4029 31159 4063
rect 36829 4029 36863 4063
rect 19717 3961 19751 3995
rect 20269 3961 20303 3995
rect 22937 3961 22971 3995
rect 32873 3961 32907 3995
rect 37657 3961 37691 3995
rect 16221 3893 16255 3927
rect 18889 3893 18923 3927
rect 20821 3893 20855 3927
rect 21465 3893 21499 3927
rect 28653 3893 28687 3927
rect 30867 3893 30901 3927
rect 31769 3893 31803 3927
rect 33885 3893 33919 3927
rect 34529 3893 34563 3927
rect 35081 3893 35115 3927
rect 35633 3893 35667 3927
rect 36093 3893 36127 3927
rect 38209 3893 38243 3927
rect 12081 3689 12115 3723
rect 13185 3689 13219 3723
rect 16129 3689 16163 3723
rect 19625 3689 19659 3723
rect 21538 3689 21572 3723
rect 28285 3689 28319 3723
rect 23029 3621 23063 3655
rect 33701 3621 33735 3655
rect 37473 3621 37507 3655
rect 17693 3553 17727 3587
rect 21281 3553 21315 3587
rect 26065 3553 26099 3587
rect 26341 3553 26375 3587
rect 28549 3553 28583 3587
rect 29101 3553 29135 3587
rect 29745 3553 29779 3587
rect 31942 3553 31976 3587
rect 38025 3553 38059 3587
rect 1593 3485 1627 3519
rect 2237 3485 2271 3519
rect 12173 3485 12207 3519
rect 14473 3485 14507 3519
rect 16221 3485 16255 3519
rect 16865 3485 16899 3519
rect 17969 3485 18003 3519
rect 18429 3485 18463 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 24041 3485 24075 3519
rect 37565 3485 37599 3519
rect 38209 3485 38243 3519
rect 15301 3417 15335 3451
rect 18705 3417 18739 3451
rect 30021 3417 30055 3451
rect 32229 3417 32263 3451
rect 34253 3417 34287 3451
rect 34989 3417 35023 3451
rect 35541 3417 35575 3451
rect 36093 3417 36127 3451
rect 1777 3349 1811 3383
rect 13737 3349 13771 3383
rect 16865 3349 16899 3383
rect 20269 3349 20303 3383
rect 23857 3349 23891 3383
rect 24593 3349 24627 3383
rect 26801 3349 26835 3383
rect 31493 3349 31527 3383
rect 36645 3349 36679 3383
rect 4721 3145 4755 3179
rect 13369 3145 13403 3179
rect 34069 3145 34103 3179
rect 35909 3145 35943 3179
rect 36921 3145 36955 3179
rect 17141 3077 17175 3111
rect 17233 3077 17267 3111
rect 18429 3077 18463 3111
rect 24041 3077 24075 3111
rect 24593 3077 24627 3111
rect 27445 3077 27479 3111
rect 29653 3077 29687 3111
rect 32597 3077 32631 3111
rect 1869 3009 1903 3043
rect 4905 3009 4939 3043
rect 8401 3009 8435 3043
rect 14841 3009 14875 3043
rect 15761 3009 15795 3043
rect 18521 3009 18555 3043
rect 19165 3009 19199 3043
rect 21465 3009 21499 3043
rect 22017 3009 22051 3043
rect 26617 3009 26651 3043
rect 27169 3009 27203 3043
rect 34805 3009 34839 3043
rect 36737 3009 36771 3043
rect 38025 3009 38059 3043
rect 2421 2941 2455 2975
rect 12265 2941 12299 2975
rect 14565 2941 14599 2975
rect 15577 2941 15611 2975
rect 21189 2941 21223 2975
rect 26341 2941 26375 2975
rect 29193 2941 29227 2975
rect 31401 2941 31435 2975
rect 31677 2941 31711 2975
rect 32321 2941 32355 2975
rect 12817 2873 12851 2907
rect 17693 2873 17727 2907
rect 19073 2873 19107 2907
rect 35265 2873 35299 2907
rect 1685 2805 1719 2839
rect 8309 2805 8343 2839
rect 11161 2805 11195 2839
rect 13921 2805 13955 2839
rect 16221 2805 16255 2839
rect 19717 2805 19751 2839
rect 22280 2805 22314 2839
rect 34621 2805 34655 2839
rect 37565 2805 37599 2839
rect 38209 2805 38243 2839
rect 10057 2601 10091 2635
rect 12541 2601 12575 2635
rect 18061 2601 18095 2635
rect 28917 2601 28951 2635
rect 38209 2601 38243 2635
rect 2421 2533 2455 2567
rect 9413 2533 9447 2567
rect 14289 2533 14323 2567
rect 4261 2465 4295 2499
rect 21465 2465 21499 2499
rect 22017 2465 22051 2499
rect 24685 2465 24719 2499
rect 27445 2465 27479 2499
rect 29745 2465 29779 2499
rect 31493 2465 31527 2499
rect 34069 2465 34103 2499
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 5549 2397 5583 2431
rect 6837 2397 6871 2431
rect 9873 2397 9907 2431
rect 10517 2397 10551 2431
rect 11989 2397 12023 2431
rect 13553 2397 13587 2431
rect 15209 2397 15243 2431
rect 16129 2397 16163 2431
rect 16865 2397 16899 2431
rect 17969 2397 18003 2431
rect 18613 2397 18647 2431
rect 27169 2397 27203 2431
rect 34897 2397 34931 2431
rect 35817 2397 35851 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 9229 2329 9263 2363
rect 11161 2329 11195 2363
rect 14473 2329 14507 2363
rect 21189 2329 21223 2363
rect 22293 2329 22327 2363
rect 24961 2329 24995 2363
rect 31217 2329 31251 2363
rect 33793 2329 33827 2363
rect 1685 2261 1719 2295
rect 3341 2261 3375 2295
rect 5365 2261 5399 2295
rect 6653 2261 6687 2295
rect 8493 2261 8527 2295
rect 11805 2261 11839 2295
rect 13093 2261 13127 2295
rect 13737 2261 13771 2295
rect 15301 2261 15335 2295
rect 16313 2261 16347 2295
rect 17049 2261 17083 2295
rect 18797 2261 18831 2295
rect 19717 2261 19751 2295
rect 23765 2261 23799 2295
rect 26433 2261 26467 2295
rect 32321 2261 32355 2295
rect 35081 2261 35115 2295
rect 35725 2261 35759 2295
rect 36829 2261 36863 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 17681 37451 17739 37457
rect 17681 37417 17693 37451
rect 17727 37448 17739 37451
rect 18046 37448 18052 37460
rect 17727 37420 18052 37448
rect 17727 37417 17739 37420
rect 17681 37411 17739 37417
rect 18046 37408 18052 37420
rect 18104 37408 18110 37460
rect 14550 37340 14556 37392
rect 14608 37380 14614 37392
rect 18141 37383 18199 37389
rect 18141 37380 18153 37383
rect 14608 37352 18153 37380
rect 14608 37340 14614 37352
rect 18141 37349 18153 37352
rect 18187 37349 18199 37383
rect 18141 37343 18199 37349
rect 9309 37315 9367 37321
rect 9309 37281 9321 37315
rect 9355 37312 9367 37315
rect 12437 37315 12495 37321
rect 9355 37284 9720 37312
rect 9355 37281 9367 37284
rect 9309 37275 9367 37281
rect 9692 37256 9720 37284
rect 12437 37281 12449 37315
rect 12483 37281 12495 37315
rect 12437 37275 12495 37281
rect 14461 37315 14519 37321
rect 14461 37281 14473 37315
rect 14507 37312 14519 37315
rect 14826 37312 14832 37324
rect 14507 37284 14832 37312
rect 14507 37281 14519 37284
rect 14461 37275 14519 37281
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 1857 37247 1915 37253
rect 1857 37244 1869 37247
rect 1820 37216 1869 37244
rect 1820 37204 1826 37216
rect 1857 37213 1869 37216
rect 1903 37213 1915 37247
rect 1857 37207 1915 37213
rect 2961 37247 3019 37253
rect 2961 37213 2973 37247
rect 3007 37244 3019 37247
rect 4062 37244 4068 37256
rect 3007 37216 4068 37244
rect 3007 37213 3019 37216
rect 2961 37207 3019 37213
rect 4062 37204 4068 37216
rect 4120 37204 4126 37256
rect 4893 37247 4951 37253
rect 4893 37213 4905 37247
rect 4939 37244 4951 37247
rect 6825 37247 6883 37253
rect 4939 37216 5488 37244
rect 4939 37213 4951 37216
rect 4893 37207 4951 37213
rect 5460 37120 5488 37216
rect 6825 37213 6837 37247
rect 6871 37244 6883 37247
rect 7282 37244 7288 37256
rect 6871 37216 7288 37244
rect 6871 37213 6883 37216
rect 6825 37207 6883 37213
rect 7282 37204 7288 37216
rect 7340 37204 7346 37256
rect 7377 37247 7435 37253
rect 7377 37213 7389 37247
rect 7423 37244 7435 37247
rect 7742 37244 7748 37256
rect 7423 37216 7748 37244
rect 7423 37213 7435 37216
rect 7377 37207 7435 37213
rect 7742 37204 7748 37216
rect 7800 37244 7806 37256
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 7800 37216 7941 37244
rect 7800 37204 7806 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 7929 37207 7987 37213
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9732 37216 9873 37244
rect 9732 37204 9738 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 11974 37244 11980 37256
rect 11935 37216 11980 37244
rect 9861 37207 9919 37213
rect 11974 37204 11980 37216
rect 12032 37244 12038 37256
rect 12452 37244 12480 37275
rect 14826 37272 14832 37284
rect 14884 37312 14890 37324
rect 14921 37315 14979 37321
rect 14921 37312 14933 37315
rect 14884 37284 14933 37312
rect 14884 37272 14890 37284
rect 14921 37281 14933 37284
rect 14967 37281 14979 37315
rect 14921 37275 14979 37281
rect 16301 37315 16359 37321
rect 16301 37281 16313 37315
rect 16347 37312 16359 37315
rect 16666 37312 16672 37324
rect 16347 37284 16672 37312
rect 16347 37281 16359 37284
rect 16301 37275 16359 37281
rect 16666 37272 16672 37284
rect 16724 37272 16730 37324
rect 16758 37272 16764 37324
rect 16816 37312 16822 37324
rect 17129 37315 17187 37321
rect 17129 37312 17141 37315
rect 16816 37284 17141 37312
rect 16816 37272 16822 37284
rect 17129 37281 17141 37284
rect 17175 37281 17187 37315
rect 17129 37275 17187 37281
rect 20809 37315 20867 37321
rect 20809 37281 20821 37315
rect 20855 37281 20867 37315
rect 20809 37275 20867 37281
rect 21453 37315 21511 37321
rect 21453 37281 21465 37315
rect 21499 37312 21511 37315
rect 21910 37312 21916 37324
rect 21499 37284 21916 37312
rect 21499 37281 21511 37284
rect 21453 37275 21511 37281
rect 13262 37244 13268 37256
rect 12032 37216 12480 37244
rect 13223 37216 13268 37244
rect 12032 37204 12038 37216
rect 13262 37204 13268 37216
rect 13320 37204 13326 37256
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 16684 37244 16712 37272
rect 16945 37247 17003 37253
rect 16945 37244 16957 37247
rect 16684 37216 16957 37244
rect 16945 37213 16957 37216
rect 16991 37213 17003 37247
rect 16945 37207 17003 37213
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 20346 37244 20352 37256
rect 20307 37216 20352 37244
rect 18325 37207 18383 37213
rect 20346 37204 20352 37216
rect 20404 37244 20410 37256
rect 20824 37244 20852 37275
rect 21910 37272 21916 37284
rect 21968 37312 21974 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21968 37284 22017 37312
rect 21968 37272 21974 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 35069 37315 35127 37321
rect 35069 37281 35081 37315
rect 35115 37312 35127 37315
rect 35434 37312 35440 37324
rect 35115 37284 35440 37312
rect 35115 37281 35127 37284
rect 35069 37275 35127 37281
rect 35434 37272 35440 37284
rect 35492 37312 35498 37324
rect 35529 37315 35587 37321
rect 35529 37312 35541 37315
rect 35492 37284 35541 37312
rect 35492 37272 35498 37284
rect 35529 37281 35541 37284
rect 35575 37281 35587 37315
rect 38286 37312 38292 37324
rect 38247 37284 38292 37312
rect 35529 37275 35587 37281
rect 38286 37272 38292 37284
rect 38344 37272 38350 37324
rect 22278 37244 22284 37256
rect 20404 37216 20852 37244
rect 22239 37216 22284 37244
rect 20404 37204 20410 37216
rect 22278 37204 22284 37216
rect 22336 37204 22342 37256
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 23293 37247 23351 37253
rect 23293 37244 23305 37247
rect 22612 37216 23305 37244
rect 22612 37204 22618 37216
rect 23293 37213 23305 37216
rect 23339 37213 23351 37247
rect 23293 37207 23351 37213
rect 23382 37204 23388 37256
rect 23440 37244 23446 37256
rect 25225 37247 25283 37253
rect 25225 37244 25237 37247
rect 23440 37216 25237 37244
rect 23440 37204 23446 37216
rect 25225 37213 25237 37216
rect 25271 37213 25283 37247
rect 27154 37244 27160 37256
rect 27115 37216 27160 37244
rect 25225 37207 25283 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 27985 37247 28043 37253
rect 27985 37213 27997 37247
rect 28031 37244 28043 37247
rect 28442 37244 28448 37256
rect 28031 37216 28448 37244
rect 28031 37213 28043 37216
rect 27985 37207 28043 37213
rect 28442 37204 28448 37216
rect 28500 37204 28506 37256
rect 30377 37247 30435 37253
rect 30377 37213 30389 37247
rect 30423 37244 30435 37247
rect 30466 37244 30472 37256
rect 30423 37216 30472 37244
rect 30423 37213 30435 37216
rect 30377 37207 30435 37213
rect 30466 37204 30472 37216
rect 30524 37204 30530 37256
rect 32582 37244 32588 37256
rect 32543 37216 32588 37244
rect 32582 37204 32588 37216
rect 32640 37204 32646 37256
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 35802 37244 35808 37256
rect 35763 37216 35808 37244
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 37826 37204 37832 37256
rect 37884 37244 37890 37256
rect 38013 37247 38071 37253
rect 38013 37244 38025 37247
rect 37884 37216 38025 37244
rect 37884 37204 37890 37216
rect 38013 37213 38025 37216
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 1673 37111 1731 37117
rect 1673 37108 1685 37111
rect 1360 37080 1685 37108
rect 1360 37068 1366 37080
rect 1673 37077 1685 37080
rect 1719 37077 1731 37111
rect 2774 37108 2780 37120
rect 2735 37080 2780 37108
rect 1673 37071 1731 37077
rect 2774 37068 2780 37080
rect 2832 37068 2838 37120
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4709 37111 4767 37117
rect 4709 37108 4721 37111
rect 4672 37080 4721 37108
rect 4672 37068 4678 37080
rect 4709 37077 4721 37080
rect 4755 37077 4767 37111
rect 5442 37108 5448 37120
rect 5403 37080 5448 37108
rect 4709 37071 4767 37077
rect 5442 37068 5448 37080
rect 5500 37068 5506 37120
rect 6454 37068 6460 37120
rect 6512 37108 6518 37120
rect 6641 37111 6699 37117
rect 6641 37108 6653 37111
rect 6512 37080 6653 37108
rect 6512 37068 6518 37080
rect 6641 37077 6653 37080
rect 6687 37077 6699 37111
rect 8018 37108 8024 37120
rect 7979 37080 8024 37108
rect 6641 37071 6699 37077
rect 8018 37068 8024 37080
rect 8076 37068 8082 37120
rect 9950 37108 9956 37120
rect 9911 37080 9956 37108
rect 9950 37068 9956 37080
rect 10008 37068 10014 37120
rect 11606 37068 11612 37120
rect 11664 37108 11670 37120
rect 11793 37111 11851 37117
rect 11793 37108 11805 37111
rect 11664 37080 11805 37108
rect 11664 37068 11670 37080
rect 11793 37077 11805 37080
rect 11839 37077 11851 37111
rect 11793 37071 11851 37077
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 13081 37111 13139 37117
rect 13081 37108 13093 37111
rect 12952 37080 13093 37108
rect 12952 37068 12958 37080
rect 13081 37077 13093 37080
rect 13127 37077 13139 37111
rect 13081 37071 13139 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20165 37111 20223 37117
rect 20165 37108 20177 37111
rect 20036 37080 20177 37108
rect 20036 37068 20042 37080
rect 20165 37077 20177 37080
rect 20211 37077 20223 37111
rect 20165 37071 20223 37077
rect 23198 37068 23204 37120
rect 23256 37108 23262 37120
rect 23477 37111 23535 37117
rect 23477 37108 23489 37111
rect 23256 37080 23489 37108
rect 23256 37068 23262 37080
rect 23477 37077 23489 37080
rect 23523 37077 23535 37111
rect 23477 37071 23535 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25409 37111 25467 37117
rect 25409 37108 25421 37111
rect 25188 37080 25421 37108
rect 25188 37068 25194 37080
rect 25409 37077 25421 37080
rect 25455 37077 25467 37111
rect 25409 37071 25467 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28350 37068 28356 37120
rect 28408 37108 28414 37120
rect 28629 37111 28687 37117
rect 28629 37108 28641 37111
rect 28408 37080 28641 37108
rect 28408 37068 28414 37080
rect 28629 37077 28641 37080
rect 28675 37077 28687 37111
rect 28629 37071 28687 37077
rect 30374 37068 30380 37120
rect 30432 37108 30438 37120
rect 30561 37111 30619 37117
rect 30561 37108 30573 37111
rect 30432 37080 30573 37108
rect 30432 37068 30438 37080
rect 30561 37077 30573 37080
rect 30607 37077 30619 37111
rect 30561 37071 30619 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32401 37111 32459 37117
rect 32401 37108 32413 37111
rect 32272 37080 32413 37108
rect 32272 37068 32278 37080
rect 32401 37077 32413 37080
rect 32447 37077 32459 37111
rect 32401 37071 32459 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 5442 36864 5448 36916
rect 5500 36904 5506 36916
rect 21174 36904 21180 36916
rect 5500 36876 21180 36904
rect 5500 36864 5506 36876
rect 21174 36864 21180 36876
rect 21232 36864 21238 36916
rect 22554 36904 22560 36916
rect 22515 36876 22560 36904
rect 22554 36864 22560 36876
rect 22612 36864 22618 36916
rect 27893 36907 27951 36913
rect 27893 36873 27905 36907
rect 27939 36904 27951 36907
rect 33594 36904 33600 36916
rect 27939 36876 33600 36904
rect 27939 36873 27951 36876
rect 27893 36867 27951 36873
rect 33594 36864 33600 36876
rect 33652 36864 33658 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37645 36907 37703 36913
rect 37645 36904 37657 36907
rect 37424 36876 37657 36904
rect 37424 36864 37430 36876
rect 37645 36873 37657 36876
rect 37691 36873 37703 36907
rect 38286 36904 38292 36916
rect 38247 36876 38292 36904
rect 37645 36867 37703 36873
rect 38286 36864 38292 36876
rect 38344 36864 38350 36916
rect 2409 36839 2467 36845
rect 2409 36805 2421 36839
rect 2455 36836 2467 36839
rect 2866 36836 2872 36848
rect 2455 36808 2872 36836
rect 2455 36805 2467 36808
rect 2409 36799 2467 36805
rect 2866 36796 2872 36808
rect 2924 36796 2930 36848
rect 22278 36796 22284 36848
rect 22336 36836 22342 36848
rect 22336 36808 26234 36836
rect 22336 36796 22342 36808
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 2958 36768 2964 36780
rect 1719 36740 2964 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 2958 36728 2964 36740
rect 3016 36768 3022 36780
rect 3053 36771 3111 36777
rect 3053 36768 3065 36771
rect 3016 36740 3065 36768
rect 3016 36728 3022 36740
rect 3053 36737 3065 36740
rect 3099 36737 3111 36771
rect 3053 36731 3111 36737
rect 10689 36771 10747 36777
rect 10689 36737 10701 36771
rect 10735 36768 10747 36771
rect 15194 36768 15200 36780
rect 10735 36740 15200 36768
rect 10735 36737 10747 36740
rect 10689 36731 10747 36737
rect 15194 36728 15200 36740
rect 15252 36768 15258 36780
rect 15930 36768 15936 36780
rect 15252 36740 15936 36768
rect 15252 36728 15258 36740
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 22373 36771 22431 36777
rect 22373 36737 22385 36771
rect 22419 36768 22431 36771
rect 23106 36768 23112 36780
rect 22419 36740 23112 36768
rect 22419 36737 22431 36740
rect 22373 36731 22431 36737
rect 23106 36728 23112 36740
rect 23164 36728 23170 36780
rect 26206 36768 26234 36808
rect 27709 36771 27767 36777
rect 27709 36768 27721 36771
rect 26206 36740 27721 36768
rect 27709 36737 27721 36740
rect 27755 36737 27767 36771
rect 27709 36731 27767 36737
rect 36814 36728 36820 36780
rect 36872 36768 36878 36780
rect 37461 36771 37519 36777
rect 37461 36768 37473 36771
rect 36872 36740 37473 36768
rect 36872 36728 36878 36740
rect 37461 36737 37473 36740
rect 37507 36737 37519 36771
rect 37461 36731 37519 36737
rect 1857 36635 1915 36641
rect 1857 36601 1869 36635
rect 1903 36632 1915 36635
rect 2038 36632 2044 36644
rect 1903 36604 2044 36632
rect 1903 36601 1915 36604
rect 1857 36595 1915 36601
rect 2038 36592 2044 36604
rect 2096 36592 2102 36644
rect 2593 36635 2651 36641
rect 2593 36601 2605 36635
rect 2639 36632 2651 36635
rect 17494 36632 17500 36644
rect 2639 36604 17500 36632
rect 2639 36601 2651 36604
rect 2593 36595 2651 36601
rect 17494 36592 17500 36604
rect 17552 36592 17558 36644
rect 7282 36524 7288 36576
rect 7340 36564 7346 36576
rect 10505 36567 10563 36573
rect 10505 36564 10517 36567
rect 7340 36536 10517 36564
rect 7340 36524 7346 36536
rect 10505 36533 10517 36536
rect 10551 36533 10563 36567
rect 10505 36527 10563 36533
rect 13262 36524 13268 36576
rect 13320 36564 13326 36576
rect 13357 36567 13415 36573
rect 13357 36564 13369 36567
rect 13320 36536 13369 36564
rect 13320 36524 13326 36536
rect 13357 36533 13369 36536
rect 13403 36533 13415 36567
rect 23106 36564 23112 36576
rect 23067 36536 23112 36564
rect 13357 36527 13415 36533
rect 23106 36524 23112 36536
rect 23164 36524 23170 36576
rect 36814 36564 36820 36576
rect 36775 36536 36820 36564
rect 36814 36524 36820 36536
rect 36872 36524 36878 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 2409 36363 2467 36369
rect 2409 36329 2421 36363
rect 2455 36360 2467 36363
rect 2866 36360 2872 36372
rect 2455 36332 2872 36360
rect 2455 36329 2467 36332
rect 2409 36323 2467 36329
rect 2866 36320 2872 36332
rect 2924 36320 2930 36372
rect 23106 36320 23112 36372
rect 23164 36360 23170 36372
rect 35802 36360 35808 36372
rect 23164 36332 35808 36360
rect 23164 36320 23170 36332
rect 35802 36320 35808 36332
rect 35860 36320 35866 36372
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37240 36332 37473 36360
rect 37240 36320 37246 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 38197 36363 38255 36369
rect 38197 36329 38209 36363
rect 38243 36360 38255 36363
rect 38654 36360 38660 36372
rect 38243 36332 38660 36360
rect 38243 36329 38255 36332
rect 38197 36323 38255 36329
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 1854 36156 1860 36168
rect 1815 36128 1860 36156
rect 1854 36116 1860 36128
rect 1912 36116 1918 36168
rect 37277 36159 37335 36165
rect 37277 36156 37289 36159
rect 36740 36128 37289 36156
rect 36740 36032 36768 36128
rect 37277 36125 37289 36128
rect 37323 36125 37335 36159
rect 38010 36156 38016 36168
rect 37971 36128 38016 36156
rect 37277 36119 37335 36125
rect 38010 36116 38016 36128
rect 38068 36116 38074 36168
rect 1670 36020 1676 36032
rect 1631 35992 1676 36020
rect 1670 35980 1676 35992
rect 1728 35980 1734 36032
rect 36722 36020 36728 36032
rect 36683 35992 36728 36020
rect 36722 35980 36728 35992
rect 36780 35980 36786 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 36909 35615 36967 35621
rect 36909 35581 36921 35615
rect 36955 35612 36967 35615
rect 37458 35612 37464 35624
rect 36955 35584 37464 35612
rect 36955 35581 36967 35584
rect 36909 35575 36967 35581
rect 37458 35572 37464 35584
rect 37516 35572 37522 35624
rect 37734 35612 37740 35624
rect 37695 35584 37740 35612
rect 37734 35572 37740 35584
rect 37792 35572 37798 35624
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 21637 35275 21695 35281
rect 21637 35241 21649 35275
rect 21683 35272 21695 35275
rect 23382 35272 23388 35284
rect 21683 35244 23388 35272
rect 21683 35241 21695 35244
rect 21637 35235 21695 35241
rect 23382 35232 23388 35244
rect 23440 35232 23446 35284
rect 29917 35275 29975 35281
rect 29917 35241 29929 35275
rect 29963 35272 29975 35275
rect 30466 35272 30472 35284
rect 29963 35244 30472 35272
rect 29963 35241 29975 35244
rect 29917 35235 29975 35241
rect 30466 35232 30472 35244
rect 30524 35232 30530 35284
rect 38010 35272 38016 35284
rect 37971 35244 38016 35272
rect 38010 35232 38016 35244
rect 38068 35232 38074 35284
rect 21082 35028 21088 35080
rect 21140 35068 21146 35080
rect 21453 35071 21511 35077
rect 21453 35068 21465 35071
rect 21140 35040 21465 35068
rect 21140 35028 21146 35040
rect 21453 35037 21465 35040
rect 21499 35068 21511 35071
rect 22097 35071 22155 35077
rect 22097 35068 22109 35071
rect 21499 35040 22109 35068
rect 21499 35037 21511 35040
rect 21453 35031 21511 35037
rect 22097 35037 22109 35040
rect 22143 35037 22155 35071
rect 22097 35031 22155 35037
rect 29638 35028 29644 35080
rect 29696 35068 29702 35080
rect 29733 35071 29791 35077
rect 29733 35068 29745 35071
rect 29696 35040 29745 35068
rect 29696 35028 29702 35040
rect 29733 35037 29745 35040
rect 29779 35068 29791 35071
rect 30377 35071 30435 35077
rect 30377 35068 30389 35071
rect 29779 35040 30389 35068
rect 29779 35037 29791 35040
rect 29733 35031 29791 35037
rect 30377 35037 30389 35040
rect 30423 35037 30435 35071
rect 30377 35031 30435 35037
rect 30742 35028 30748 35080
rect 30800 35068 30806 35080
rect 37734 35068 37740 35080
rect 30800 35040 37740 35068
rect 30800 35028 30806 35040
rect 37734 35028 37740 35040
rect 37792 35068 37798 35080
rect 37829 35071 37887 35077
rect 37829 35068 37841 35071
rect 37792 35040 37841 35068
rect 37792 35028 37798 35040
rect 37829 35037 37841 35040
rect 37875 35037 37887 35071
rect 37829 35031 37887 35037
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1854 34688 1860 34740
rect 1912 34728 1918 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 1912 34700 2421 34728
rect 1912 34688 1918 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 2409 34691 2467 34697
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 2130 34592 2136 34604
rect 1903 34564 2136 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 2130 34552 2136 34564
rect 2188 34552 2194 34604
rect 2501 34595 2559 34601
rect 2501 34561 2513 34595
rect 2547 34592 2559 34595
rect 2547 34564 3096 34592
rect 2547 34561 2559 34564
rect 2501 34555 2559 34561
rect 3068 34533 3096 34564
rect 3053 34527 3111 34533
rect 3053 34493 3065 34527
rect 3099 34524 3111 34527
rect 18138 34524 18144 34536
rect 3099 34496 18144 34524
rect 3099 34493 3111 34496
rect 3053 34487 3111 34493
rect 18138 34484 18144 34496
rect 18196 34484 18202 34536
rect 1670 34388 1676 34400
rect 1631 34360 1676 34388
rect 1670 34348 1676 34360
rect 1728 34348 1734 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 2041 33847 2099 33853
rect 2041 33813 2053 33847
rect 2087 33844 2099 33847
rect 2130 33844 2136 33856
rect 2087 33816 2136 33844
rect 2087 33813 2099 33816
rect 2041 33807 2099 33813
rect 2130 33804 2136 33816
rect 2188 33804 2194 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 37476 33476 38025 33504
rect 15838 33260 15844 33312
rect 15896 33300 15902 33312
rect 37476 33309 37504 33476
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 37461 33303 37519 33309
rect 37461 33300 37473 33303
rect 15896 33272 37473 33300
rect 15896 33260 15902 33272
rect 37461 33269 37473 33272
rect 37507 33269 37519 33303
rect 37461 33263 37519 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 32582 32552 32588 32564
rect 32543 32524 32588 32552
rect 32582 32512 32588 32524
rect 32640 32512 32646 32564
rect 1578 32376 1584 32428
rect 1636 32416 1642 32428
rect 1673 32419 1731 32425
rect 1673 32416 1685 32419
rect 1636 32388 1685 32416
rect 1636 32376 1642 32388
rect 1673 32385 1685 32388
rect 1719 32385 1731 32419
rect 1673 32379 1731 32385
rect 27982 32376 27988 32428
rect 28040 32416 28046 32428
rect 32677 32419 32735 32425
rect 32677 32416 32689 32419
rect 28040 32388 32689 32416
rect 28040 32376 28046 32388
rect 32677 32385 32689 32388
rect 32723 32416 32735 32419
rect 33137 32419 33195 32425
rect 33137 32416 33149 32419
rect 32723 32388 33149 32416
rect 32723 32385 32735 32388
rect 32677 32379 32735 32385
rect 33137 32385 33149 32388
rect 33183 32385 33195 32419
rect 33137 32379 33195 32385
rect 29638 32308 29644 32360
rect 29696 32348 29702 32360
rect 38013 32351 38071 32357
rect 38013 32348 38025 32351
rect 29696 32320 38025 32348
rect 29696 32308 29702 32320
rect 38013 32317 38025 32320
rect 38059 32317 38071 32351
rect 38286 32348 38292 32360
rect 38247 32320 38292 32348
rect 38013 32311 38071 32317
rect 38286 32308 38292 32320
rect 38344 32308 38350 32360
rect 1765 32215 1823 32221
rect 1765 32181 1777 32215
rect 1811 32212 1823 32215
rect 21082 32212 21088 32224
rect 1811 32184 21088 32212
rect 1811 32181 1823 32184
rect 1765 32175 1823 32181
rect 21082 32172 21088 32184
rect 21140 32172 21146 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 38286 32008 38292 32020
rect 38247 31980 38292 32008
rect 38286 31968 38292 31980
rect 38344 31968 38350 32020
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 1854 30648 1860 30660
rect 1815 30620 1860 30648
rect 1854 30608 1860 30620
rect 1912 30608 1918 30660
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1670 30376 1676 30388
rect 1631 30348 1676 30376
rect 1670 30336 1676 30348
rect 1728 30336 1734 30388
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30240 11943 30243
rect 38010 30240 38016 30252
rect 11931 30212 12480 30240
rect 37971 30212 38016 30240
rect 11931 30209 11943 30212
rect 11885 30203 11943 30209
rect 4062 30064 4068 30116
rect 4120 30104 4126 30116
rect 11793 30107 11851 30113
rect 11793 30104 11805 30107
rect 4120 30076 11805 30104
rect 4120 30064 4126 30076
rect 11793 30073 11805 30076
rect 11839 30073 11851 30107
rect 11793 30067 11851 30073
rect 12452 30048 12480 30212
rect 38010 30200 38016 30212
rect 38068 30200 38074 30252
rect 12434 30036 12440 30048
rect 12395 30008 12440 30036
rect 12434 29996 12440 30008
rect 12492 29996 12498 30048
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 22186 29792 22192 29844
rect 22244 29832 22250 29844
rect 22373 29835 22431 29841
rect 22373 29832 22385 29835
rect 22244 29804 22385 29832
rect 22244 29792 22250 29804
rect 22373 29801 22385 29804
rect 22419 29832 22431 29835
rect 23106 29832 23112 29844
rect 22419 29804 23112 29832
rect 22419 29801 22431 29804
rect 22373 29795 22431 29801
rect 23106 29792 23112 29804
rect 23164 29792 23170 29844
rect 38010 29832 38016 29844
rect 37971 29804 38016 29832
rect 38010 29792 38016 29804
rect 38068 29792 38074 29844
rect 37826 29628 37832 29640
rect 37787 29600 37832 29628
rect 37826 29588 37832 29600
rect 37884 29588 37890 29640
rect 20073 29563 20131 29569
rect 20073 29529 20085 29563
rect 20119 29560 20131 29563
rect 20625 29563 20683 29569
rect 20625 29560 20637 29563
rect 20119 29532 20637 29560
rect 20119 29529 20131 29532
rect 20073 29523 20131 29529
rect 20625 29529 20637 29532
rect 20671 29560 20683 29563
rect 20714 29560 20720 29572
rect 20671 29532 20720 29560
rect 20671 29529 20683 29532
rect 20625 29523 20683 29529
rect 20714 29520 20720 29532
rect 20772 29520 20778 29572
rect 20809 29563 20867 29569
rect 20809 29529 20821 29563
rect 20855 29560 20867 29563
rect 20855 29532 26234 29560
rect 20855 29529 20867 29532
rect 20809 29523 20867 29529
rect 26206 29492 26234 29532
rect 36722 29492 36728 29504
rect 26206 29464 36728 29492
rect 36722 29452 36728 29464
rect 36780 29452 36786 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1578 29112 1584 29164
rect 1636 29152 1642 29164
rect 1673 29155 1731 29161
rect 1673 29152 1685 29155
rect 1636 29124 1685 29152
rect 1636 29112 1642 29124
rect 1673 29121 1685 29124
rect 1719 29121 1731 29155
rect 22186 29152 22192 29164
rect 22147 29124 22192 29152
rect 1673 29115 1731 29121
rect 22186 29112 22192 29124
rect 22244 29112 22250 29164
rect 22278 29112 22284 29164
rect 22336 29152 22342 29164
rect 22649 29155 22707 29161
rect 22649 29152 22661 29155
rect 22336 29124 22661 29152
rect 22336 29112 22342 29124
rect 22649 29121 22661 29124
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 12434 29044 12440 29096
rect 12492 29084 12498 29096
rect 23750 29084 23756 29096
rect 12492 29056 23756 29084
rect 12492 29044 12498 29056
rect 23750 29044 23756 29056
rect 23808 29044 23814 29096
rect 1857 29019 1915 29025
rect 1857 28985 1869 29019
rect 1903 29016 1915 29019
rect 20714 29016 20720 29028
rect 1903 28988 20720 29016
rect 1903 28985 1915 28988
rect 1857 28979 1915 28985
rect 20714 28976 20720 28988
rect 20772 28976 20778 29028
rect 22097 29019 22155 29025
rect 22097 28985 22109 29019
rect 22143 29016 22155 29019
rect 22186 29016 22192 29028
rect 22143 28988 22192 29016
rect 22143 28985 22155 28988
rect 22097 28979 22155 28985
rect 22186 28976 22192 28988
rect 22244 28976 22250 29028
rect 22741 29019 22799 29025
rect 22741 28985 22753 29019
rect 22787 29016 22799 29019
rect 23566 29016 23572 29028
rect 22787 28988 23572 29016
rect 22787 28985 22799 28988
rect 22741 28979 22799 28985
rect 23566 28976 23572 28988
rect 23624 28976 23630 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 21174 28744 21180 28756
rect 21135 28716 21180 28744
rect 21174 28704 21180 28716
rect 21232 28704 21238 28756
rect 1578 28676 1584 28688
rect 1539 28648 1584 28676
rect 1578 28636 1584 28648
rect 1636 28636 1642 28688
rect 21269 28475 21327 28481
rect 21269 28441 21281 28475
rect 21315 28441 21327 28475
rect 21269 28435 21327 28441
rect 21284 28404 21312 28435
rect 21913 28407 21971 28413
rect 21913 28404 21925 28407
rect 21284 28376 21925 28404
rect 21913 28373 21925 28376
rect 21959 28404 21971 28407
rect 23382 28404 23388 28416
rect 21959 28376 23388 28404
rect 21959 28373 21971 28376
rect 21913 28367 21971 28373
rect 23382 28364 23388 28376
rect 23440 28364 23446 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 15930 28064 15936 28076
rect 15891 28036 15936 28064
rect 15930 28024 15936 28036
rect 15988 28024 15994 28076
rect 38013 28067 38071 28073
rect 38013 28064 38025 28067
rect 37476 28036 38025 28064
rect 16025 27863 16083 27869
rect 16025 27829 16037 27863
rect 16071 27860 16083 27863
rect 16114 27860 16120 27872
rect 16071 27832 16120 27860
rect 16071 27829 16083 27832
rect 16025 27823 16083 27829
rect 16114 27820 16120 27832
rect 16172 27820 16178 27872
rect 20622 27820 20628 27872
rect 20680 27860 20686 27872
rect 37476 27869 37504 28036
rect 38013 28033 38025 28036
rect 38059 28033 38071 28067
rect 38013 28027 38071 28033
rect 38194 27928 38200 27940
rect 38155 27900 38200 27928
rect 38194 27888 38200 27900
rect 38252 27888 38258 27940
rect 37461 27863 37519 27869
rect 37461 27860 37473 27863
rect 20680 27832 37473 27860
rect 20680 27820 20686 27832
rect 37461 27829 37473 27832
rect 37507 27829 37519 27863
rect 37461 27823 37519 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 23382 27616 23388 27668
rect 23440 27656 23446 27668
rect 38010 27656 38016 27668
rect 23440 27628 38016 27656
rect 23440 27616 23446 27628
rect 38010 27616 38016 27628
rect 38068 27616 38074 27668
rect 30742 27452 30748 27464
rect 30703 27424 30748 27452
rect 30742 27412 30748 27424
rect 30800 27412 30806 27464
rect 27798 27276 27804 27328
rect 27856 27316 27862 27328
rect 30653 27319 30711 27325
rect 30653 27316 30665 27319
rect 27856 27288 30665 27316
rect 27856 27276 27862 27288
rect 30653 27285 30665 27288
rect 30699 27285 30711 27319
rect 30653 27279 30711 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 19613 27115 19671 27121
rect 19613 27081 19625 27115
rect 19659 27112 19671 27115
rect 20622 27112 20628 27124
rect 19659 27084 20628 27112
rect 19659 27081 19671 27084
rect 19613 27075 19671 27081
rect 20622 27072 20628 27084
rect 20680 27072 20686 27124
rect 38010 27044 38016 27056
rect 37971 27016 38016 27044
rect 38010 27004 38016 27016
rect 38068 27004 38074 27056
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26976 1915 26979
rect 6822 26976 6828 26988
rect 1903 26948 6828 26976
rect 1903 26945 1915 26948
rect 1857 26939 1915 26945
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 19429 26979 19487 26985
rect 19429 26976 19441 26979
rect 16546 26948 19441 26976
rect 2038 26868 2044 26920
rect 2096 26908 2102 26920
rect 16546 26908 16574 26948
rect 19429 26945 19441 26948
rect 19475 26976 19487 26979
rect 20070 26976 20076 26988
rect 19475 26948 20076 26976
rect 19475 26945 19487 26948
rect 19429 26939 19487 26945
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 37553 26979 37611 26985
rect 37553 26945 37565 26979
rect 37599 26976 37611 26979
rect 38194 26976 38200 26988
rect 37599 26948 38200 26976
rect 37599 26945 37611 26948
rect 37553 26939 37611 26945
rect 38194 26936 38200 26948
rect 38252 26936 38258 26988
rect 2096 26880 16574 26908
rect 2096 26868 2102 26880
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1762 26024 1768 26036
rect 1723 25996 1768 26024
rect 1762 25984 1768 25996
rect 1820 25984 1826 26036
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25888 2007 25891
rect 2038 25888 2044 25900
rect 1995 25860 2044 25888
rect 1995 25857 2007 25860
rect 1949 25851 2007 25857
rect 2038 25848 2044 25860
rect 2096 25888 2102 25900
rect 2409 25891 2467 25897
rect 2409 25888 2421 25891
rect 2096 25860 2421 25888
rect 2096 25848 2102 25860
rect 2409 25857 2421 25860
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 21082 25440 21088 25492
rect 21140 25480 21146 25492
rect 21177 25483 21235 25489
rect 21177 25480 21189 25483
rect 21140 25452 21189 25480
rect 21140 25440 21146 25452
rect 21177 25449 21189 25452
rect 21223 25449 21235 25483
rect 21177 25443 21235 25449
rect 28353 25483 28411 25489
rect 28353 25449 28365 25483
rect 28399 25480 28411 25483
rect 29638 25480 29644 25492
rect 28399 25452 29644 25480
rect 28399 25449 28411 25452
rect 28353 25443 28411 25449
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 1946 25276 1952 25288
rect 1903 25248 1952 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 1946 25236 1952 25248
rect 2004 25236 2010 25288
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25276 20775 25279
rect 21082 25276 21088 25288
rect 20763 25248 21088 25276
rect 20763 25245 20775 25248
rect 20717 25239 20775 25245
rect 21082 25236 21088 25248
rect 21140 25236 21146 25288
rect 27801 25279 27859 25285
rect 27801 25245 27813 25279
rect 27847 25276 27859 25279
rect 28368 25276 28396 25443
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 27847 25248 28396 25276
rect 32125 25279 32183 25285
rect 27847 25245 27859 25248
rect 27801 25239 27859 25245
rect 32125 25245 32137 25279
rect 32171 25276 32183 25279
rect 37826 25276 37832 25288
rect 32171 25248 37832 25276
rect 32171 25245 32183 25248
rect 32125 25239 32183 25245
rect 37826 25236 37832 25248
rect 37884 25236 37890 25288
rect 20530 25100 20536 25152
rect 20588 25140 20594 25152
rect 20625 25143 20683 25149
rect 20625 25140 20637 25143
rect 20588 25112 20637 25140
rect 20588 25100 20594 25112
rect 20625 25109 20637 25112
rect 20671 25109 20683 25143
rect 20625 25103 20683 25109
rect 26694 25100 26700 25152
rect 26752 25140 26758 25152
rect 27709 25143 27767 25149
rect 27709 25140 27721 25143
rect 26752 25112 27721 25140
rect 26752 25100 26758 25112
rect 27709 25109 27721 25112
rect 27755 25109 27767 25143
rect 32030 25140 32036 25152
rect 31991 25112 32036 25140
rect 27709 25103 27767 25109
rect 32030 25100 32036 25112
rect 32088 25100 32094 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24769 25835 24803
rect 38010 24800 38016 24812
rect 37971 24772 38016 24800
rect 25777 24763 25835 24769
rect 25792 24596 25820 24763
rect 38010 24760 38016 24772
rect 38068 24760 38074 24812
rect 25961 24667 26019 24673
rect 25961 24633 25973 24667
rect 26007 24664 26019 24667
rect 27154 24664 27160 24676
rect 26007 24636 27160 24664
rect 26007 24633 26019 24636
rect 25961 24627 26019 24633
rect 27154 24624 27160 24636
rect 27212 24624 27218 24676
rect 26513 24599 26571 24605
rect 26513 24596 26525 24599
rect 25792 24568 26525 24596
rect 26513 24565 26525 24568
rect 26559 24596 26571 24599
rect 29914 24596 29920 24608
rect 26559 24568 29920 24596
rect 26559 24565 26571 24568
rect 26513 24559 26571 24565
rect 29914 24556 29920 24568
rect 29972 24556 29978 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 11974 24080 11980 24132
rect 12032 24120 12038 24132
rect 21266 24120 21272 24132
rect 12032 24092 21272 24120
rect 12032 24080 12038 24092
rect 21266 24080 21272 24092
rect 21324 24080 21330 24132
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1857 23715 1915 23721
rect 1857 23681 1869 23715
rect 1903 23712 1915 23715
rect 2866 23712 2872 23724
rect 1903 23684 2872 23712
rect 1903 23681 1915 23684
rect 1857 23675 1915 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 1670 23508 1676 23520
rect 1631 23480 1676 23508
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 20070 22720 20076 22772
rect 20128 22760 20134 22772
rect 20257 22763 20315 22769
rect 20257 22760 20269 22763
rect 20128 22732 20269 22760
rect 20128 22720 20134 22732
rect 20257 22729 20269 22732
rect 20303 22729 20315 22763
rect 20257 22723 20315 22729
rect 19613 22627 19671 22633
rect 19613 22593 19625 22627
rect 19659 22624 19671 22627
rect 20088 22624 20116 22720
rect 19659 22596 20116 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 34054 22584 34060 22636
rect 34112 22624 34118 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 34112 22596 38025 22624
rect 34112 22584 34118 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 19705 22423 19763 22429
rect 19705 22389 19717 22423
rect 19751 22420 19763 22423
rect 20898 22420 20904 22432
rect 19751 22392 20904 22420
rect 19751 22389 19763 22392
rect 19705 22383 19763 22389
rect 20898 22380 20904 22392
rect 20956 22380 20962 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 20717 21675 20775 21681
rect 20717 21641 20729 21675
rect 20763 21672 20775 21675
rect 20806 21672 20812 21684
rect 20763 21644 20812 21672
rect 20763 21641 20775 21644
rect 20717 21635 20775 21641
rect 20806 21632 20812 21644
rect 20864 21632 20870 21684
rect 1762 21496 1768 21548
rect 1820 21536 1826 21548
rect 1857 21539 1915 21545
rect 1857 21536 1869 21539
rect 1820 21508 1869 21536
rect 1820 21496 1826 21508
rect 1857 21505 1869 21508
rect 1903 21505 1915 21539
rect 20824 21536 20852 21632
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 20824 21508 21189 21536
rect 1857 21499 1915 21505
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 37458 21496 37464 21548
rect 37516 21536 37522 21548
rect 38013 21539 38071 21545
rect 38013 21536 38025 21539
rect 37516 21508 38025 21536
rect 37516 21496 37522 21508
rect 38013 21505 38025 21508
rect 38059 21505 38071 21539
rect 38013 21499 38071 21505
rect 13262 21360 13268 21412
rect 13320 21400 13326 21412
rect 25130 21400 25136 21412
rect 13320 21372 25136 21400
rect 13320 21360 13326 21372
rect 25130 21360 25136 21372
rect 25188 21360 25194 21412
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 21269 21335 21327 21341
rect 21269 21301 21281 21335
rect 21315 21332 21327 21335
rect 22830 21332 22836 21344
rect 21315 21304 22836 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 37458 21332 37464 21344
rect 37419 21304 37464 21332
rect 37458 21292 37464 21304
rect 37516 21292 37522 21344
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1762 21128 1768 21140
rect 1723 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 6822 21088 6828 21140
rect 6880 21128 6886 21140
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 6880 21100 7113 21128
rect 6880 21088 6886 21100
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 1946 20924 1952 20936
rect 1907 20896 1952 20924
rect 1946 20884 1952 20896
rect 2004 20884 2010 20936
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 7331 20896 7880 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 7852 20797 7880 20896
rect 28092 20896 28641 20924
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 8938 20788 8944 20800
rect 7883 20760 8944 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 14458 20788 14464 20800
rect 13504 20760 14464 20788
rect 13504 20748 13510 20760
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 28092 20797 28120 20896
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28077 20791 28135 20797
rect 28077 20788 28089 20791
rect 25372 20760 28089 20788
rect 25372 20748 25378 20760
rect 28077 20757 28089 20760
rect 28123 20757 28135 20791
rect 28077 20751 28135 20757
rect 28813 20791 28871 20797
rect 28813 20757 28825 20791
rect 28859 20788 28871 20791
rect 38010 20788 38016 20800
rect 28859 20760 38016 20788
rect 28859 20757 28871 20760
rect 28813 20751 28871 20757
rect 38010 20748 38016 20760
rect 38068 20748 38074 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 23382 20544 23388 20596
rect 23440 20584 23446 20596
rect 23569 20587 23627 20593
rect 23569 20584 23581 20587
rect 23440 20556 23581 20584
rect 23440 20544 23446 20556
rect 23569 20553 23581 20556
rect 23615 20553 23627 20587
rect 23569 20547 23627 20553
rect 21082 20408 21088 20460
rect 21140 20448 21146 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21140 20420 22017 20448
rect 21140 20408 21146 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20448 22983 20451
rect 23400 20448 23428 20544
rect 22971 20420 23428 20448
rect 25225 20451 25283 20457
rect 22971 20417 22983 20420
rect 22925 20411 22983 20417
rect 25225 20417 25237 20451
rect 25271 20417 25283 20451
rect 25225 20411 25283 20417
rect 23198 20340 23204 20392
rect 23256 20380 23262 20392
rect 25240 20380 25268 20411
rect 25869 20383 25927 20389
rect 25869 20380 25881 20383
rect 23256 20352 25881 20380
rect 23256 20340 23262 20352
rect 25869 20349 25881 20352
rect 25915 20349 25927 20383
rect 25869 20343 25927 20349
rect 23017 20315 23075 20321
rect 23017 20281 23029 20315
rect 23063 20312 23075 20315
rect 25038 20312 25044 20324
rect 23063 20284 25044 20312
rect 23063 20281 23075 20284
rect 23017 20275 23075 20281
rect 25038 20272 25044 20284
rect 25096 20272 25102 20324
rect 25317 20315 25375 20321
rect 25317 20281 25329 20315
rect 25363 20312 25375 20315
rect 27522 20312 27528 20324
rect 25363 20284 27528 20312
rect 25363 20281 25375 20284
rect 25317 20275 25375 20281
rect 27522 20272 27528 20284
rect 27580 20272 27586 20324
rect 1854 20204 1860 20256
rect 1912 20244 1918 20256
rect 19797 20247 19855 20253
rect 19797 20244 19809 20247
rect 1912 20216 19809 20244
rect 1912 20204 1918 20216
rect 19797 20213 19809 20216
rect 19843 20244 19855 20247
rect 19978 20244 19984 20256
rect 19843 20216 19984 20244
rect 19843 20213 19855 20216
rect 19797 20207 19855 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 22462 20244 22468 20256
rect 22143 20216 22468 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 24394 20204 24400 20256
rect 24452 20244 24458 20256
rect 24489 20247 24547 20253
rect 24489 20244 24501 20247
rect 24452 20216 24501 20244
rect 24452 20204 24458 20216
rect 24489 20213 24501 20216
rect 24535 20213 24547 20247
rect 24489 20207 24547 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 25777 20043 25835 20049
rect 25777 20009 25789 20043
rect 25823 20040 25835 20043
rect 28442 20040 28448 20052
rect 25823 20012 28448 20040
rect 25823 20009 25835 20012
rect 25777 20003 25835 20009
rect 28442 20000 28448 20012
rect 28500 20000 28506 20052
rect 20898 19864 20904 19916
rect 20956 19904 20962 19916
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 20956 19876 22017 19904
rect 20956 19864 20962 19876
rect 22005 19873 22017 19876
rect 22051 19873 22063 19907
rect 22005 19867 22063 19873
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 37458 19904 37464 19916
rect 26936 19876 37464 19904
rect 26936 19864 26942 19876
rect 37458 19864 37464 19876
rect 37516 19864 37522 19916
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19836 1915 19839
rect 4706 19836 4712 19848
rect 1903 19808 4712 19836
rect 1903 19805 1915 19808
rect 1857 19799 1915 19805
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 21082 19836 21088 19848
rect 21043 19808 21088 19836
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25593 19839 25651 19845
rect 25593 19805 25605 19839
rect 25639 19836 25651 19839
rect 26142 19836 26148 19848
rect 25639 19808 26148 19836
rect 25639 19805 25651 19808
rect 25593 19799 25651 19805
rect 22094 19728 22100 19780
rect 22152 19768 22158 19780
rect 22646 19768 22652 19780
rect 22152 19740 22197 19768
rect 22607 19740 22652 19768
rect 22152 19728 22158 19740
rect 22646 19728 22652 19740
rect 22704 19728 22710 19780
rect 24964 19768 24992 19799
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 26786 19768 26792 19780
rect 24964 19740 26792 19768
rect 26786 19728 26792 19740
rect 26844 19728 26850 19780
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19613 19703 19671 19709
rect 19613 19700 19625 19703
rect 19392 19672 19625 19700
rect 19392 19660 19398 19672
rect 19613 19669 19625 19672
rect 19659 19669 19671 19703
rect 20254 19700 20260 19712
rect 20215 19672 20260 19700
rect 19613 19663 19671 19669
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 20993 19703 21051 19709
rect 20993 19700 21005 19703
rect 20772 19672 21005 19700
rect 20772 19660 20778 19672
rect 20993 19669 21005 19672
rect 21039 19669 21051 19703
rect 23198 19700 23204 19712
rect 23159 19672 23204 19700
rect 20993 19663 21051 19669
rect 23198 19660 23204 19672
rect 23256 19660 23262 19712
rect 24029 19703 24087 19709
rect 24029 19669 24041 19703
rect 24075 19700 24087 19703
rect 24118 19700 24124 19712
rect 24075 19672 24124 19700
rect 24075 19669 24087 19672
rect 24029 19663 24087 19669
rect 24118 19660 24124 19672
rect 24176 19660 24182 19712
rect 24857 19703 24915 19709
rect 24857 19669 24869 19703
rect 24903 19700 24915 19703
rect 25590 19700 25596 19712
rect 24903 19672 25596 19700
rect 24903 19669 24915 19672
rect 24857 19663 24915 19669
rect 25590 19660 25596 19672
rect 25648 19660 25654 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19496 20223 19499
rect 26878 19496 26884 19508
rect 20211 19468 26884 19496
rect 20211 19465 20223 19468
rect 20165 19459 20223 19465
rect 26878 19456 26884 19468
rect 26936 19456 26942 19508
rect 34054 19496 34060 19508
rect 34015 19468 34060 19496
rect 34054 19456 34060 19468
rect 34112 19456 34118 19508
rect 18690 19388 18696 19440
rect 18748 19428 18754 19440
rect 18877 19431 18935 19437
rect 18877 19428 18889 19431
rect 18748 19400 18889 19428
rect 18748 19388 18754 19400
rect 18877 19397 18889 19400
rect 18923 19397 18935 19431
rect 18877 19391 18935 19397
rect 18969 19431 19027 19437
rect 18969 19397 18981 19431
rect 19015 19428 19027 19431
rect 20530 19428 20536 19440
rect 19015 19400 20536 19428
rect 19015 19397 19027 19400
rect 18969 19391 19027 19397
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 20806 19428 20812 19440
rect 20767 19400 20812 19428
rect 20806 19388 20812 19400
rect 20864 19388 20870 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 22066 19400 22385 19428
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 21726 19320 21732 19372
rect 21784 19360 21790 19372
rect 22066 19360 22094 19400
rect 22373 19397 22385 19400
rect 22419 19397 22431 19431
rect 22373 19391 22431 19397
rect 22462 19388 22468 19440
rect 22520 19428 22526 19440
rect 22520 19400 22565 19428
rect 22520 19388 22526 19400
rect 23750 19388 23756 19440
rect 23808 19428 23814 19440
rect 23937 19431 23995 19437
rect 23937 19428 23949 19431
rect 23808 19400 23949 19428
rect 23808 19388 23814 19400
rect 23937 19397 23949 19400
rect 23983 19397 23995 19431
rect 23937 19391 23995 19397
rect 24857 19431 24915 19437
rect 24857 19397 24869 19431
rect 24903 19428 24915 19431
rect 25866 19428 25872 19440
rect 24903 19400 25872 19428
rect 24903 19397 24915 19400
rect 24857 19391 24915 19397
rect 25866 19388 25872 19400
rect 25924 19388 25930 19440
rect 26050 19428 26056 19440
rect 26011 19400 26056 19428
rect 26050 19388 26056 19400
rect 26108 19388 26114 19440
rect 26145 19431 26203 19437
rect 26145 19397 26157 19431
rect 26191 19428 26203 19431
rect 26694 19428 26700 19440
rect 26191 19400 26700 19428
rect 26191 19397 26203 19400
rect 26145 19391 26203 19397
rect 26694 19388 26700 19400
rect 26752 19388 26758 19440
rect 21784 19332 22094 19360
rect 21784 19320 21790 19332
rect 29178 19320 29184 19372
rect 29236 19360 29242 19372
rect 33965 19363 34023 19369
rect 33965 19360 33977 19363
rect 29236 19332 33977 19360
rect 29236 19320 29242 19332
rect 33965 19329 33977 19332
rect 34011 19329 34023 19363
rect 38010 19360 38016 19372
rect 37971 19332 38016 19360
rect 33965 19323 34023 19329
rect 38010 19320 38016 19332
rect 38068 19320 38074 19372
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 20898 19292 20904 19304
rect 20763 19264 20904 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 23017 19295 23075 19301
rect 23017 19261 23029 19295
rect 23063 19292 23075 19295
rect 24762 19292 24768 19304
rect 23063 19264 24768 19292
rect 23063 19261 23075 19264
rect 23017 19255 23075 19261
rect 19429 19227 19487 19233
rect 19429 19193 19441 19227
rect 19475 19224 19487 19227
rect 21008 19224 21036 19255
rect 24762 19252 24768 19264
rect 24820 19292 24826 19304
rect 24949 19295 25007 19301
rect 24949 19292 24961 19295
rect 24820 19264 24961 19292
rect 24820 19252 24826 19264
rect 24949 19261 24961 19264
rect 24995 19261 25007 19295
rect 24949 19255 25007 19261
rect 25406 19252 25412 19304
rect 25464 19292 25470 19304
rect 25501 19295 25559 19301
rect 25501 19292 25513 19295
rect 25464 19264 25513 19292
rect 25464 19252 25470 19264
rect 25501 19261 25513 19264
rect 25547 19261 25559 19295
rect 25501 19255 25559 19261
rect 19475 19196 21036 19224
rect 19475 19193 19487 19196
rect 19429 19187 19487 19193
rect 20916 19168 20944 19196
rect 20898 19116 20904 19168
rect 20956 19116 20962 19168
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 4706 18952 4712 18964
rect 4667 18924 4712 18952
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 19613 18955 19671 18961
rect 19613 18921 19625 18955
rect 19659 18952 19671 18955
rect 20806 18952 20812 18964
rect 19659 18924 20812 18952
rect 19659 18921 19671 18924
rect 19613 18915 19671 18921
rect 20806 18912 20812 18924
rect 20864 18912 20870 18964
rect 21453 18955 21511 18961
rect 21453 18921 21465 18955
rect 21499 18952 21511 18955
rect 22094 18952 22100 18964
rect 21499 18924 22100 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 22094 18912 22100 18924
rect 22152 18912 22158 18964
rect 25498 18912 25504 18964
rect 25556 18952 25562 18964
rect 30926 18952 30932 18964
rect 25556 18924 30932 18952
rect 25556 18912 25562 18924
rect 30926 18912 30932 18924
rect 30984 18912 30990 18964
rect 19536 18856 23888 18884
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 18233 18751 18291 18757
rect 4939 18720 5488 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 5460 18621 5488 18720
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18693 18751 18751 18757
rect 18693 18748 18705 18751
rect 18279 18720 18705 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18693 18717 18705 18720
rect 18739 18748 18751 18751
rect 18966 18748 18972 18760
rect 18739 18720 18972 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 18966 18708 18972 18720
rect 19024 18748 19030 18760
rect 19536 18757 19564 18856
rect 20254 18816 20260 18828
rect 20215 18788 20260 18816
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 22097 18819 22155 18825
rect 22097 18785 22109 18819
rect 22143 18816 22155 18819
rect 22186 18816 22192 18828
rect 22143 18788 22192 18816
rect 22143 18785 22155 18788
rect 22097 18779 22155 18785
rect 22186 18776 22192 18788
rect 22244 18776 22250 18828
rect 22370 18816 22376 18828
rect 22331 18788 22376 18816
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19024 18720 19533 18748
rect 19024 18708 19030 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 21082 18708 21088 18760
rect 21140 18748 21146 18760
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 21140 18720 21373 18748
rect 21140 18708 21146 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18748 23443 18751
rect 23658 18748 23664 18760
rect 23431 18720 23664 18748
rect 23431 18717 23443 18720
rect 23385 18711 23443 18717
rect 20349 18683 20407 18689
rect 20349 18649 20361 18683
rect 20395 18680 20407 18683
rect 20714 18680 20720 18692
rect 20395 18652 20720 18680
rect 20395 18649 20407 18652
rect 20349 18643 20407 18649
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 20898 18680 20904 18692
rect 20859 18652 20904 18680
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 5445 18615 5503 18621
rect 5445 18581 5457 18615
rect 5491 18612 5503 18615
rect 8018 18612 8024 18624
rect 5491 18584 8024 18612
rect 5491 18581 5503 18584
rect 5445 18575 5503 18581
rect 8018 18572 8024 18584
rect 8076 18612 8082 18624
rect 12894 18612 12900 18624
rect 8076 18584 12900 18612
rect 8076 18572 8082 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 18785 18615 18843 18621
rect 18785 18581 18797 18615
rect 18831 18612 18843 18615
rect 19426 18612 19432 18624
rect 18831 18584 19432 18612
rect 18831 18581 18843 18584
rect 18785 18575 18843 18581
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 21376 18612 21404 18711
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 23860 18757 23888 18856
rect 24026 18844 24032 18896
rect 24084 18884 24090 18896
rect 26789 18887 26847 18893
rect 26789 18884 26801 18887
rect 24084 18856 26801 18884
rect 24084 18844 24090 18856
rect 26789 18853 26801 18856
rect 26835 18884 26847 18887
rect 27154 18884 27160 18896
rect 26835 18856 27160 18884
rect 26835 18853 26847 18856
rect 26789 18847 26847 18853
rect 27154 18844 27160 18856
rect 27212 18844 27218 18896
rect 23937 18819 23995 18825
rect 23937 18785 23949 18819
rect 23983 18816 23995 18819
rect 26237 18819 26295 18825
rect 23983 18788 25820 18816
rect 23983 18785 23995 18788
rect 23937 18779 23995 18785
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 24118 18748 24124 18760
rect 23891 18720 24124 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 24118 18708 24124 18720
rect 24176 18708 24182 18760
rect 22186 18640 22192 18692
rect 22244 18680 22250 18692
rect 22244 18652 22289 18680
rect 22664 18652 23704 18680
rect 22244 18640 22250 18652
rect 22664 18624 22692 18652
rect 22554 18612 22560 18624
rect 21376 18584 22560 18612
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 22646 18572 22652 18624
rect 22704 18572 22710 18624
rect 23293 18615 23351 18621
rect 23293 18581 23305 18615
rect 23339 18612 23351 18615
rect 23382 18612 23388 18624
rect 23339 18584 23388 18612
rect 23339 18581 23351 18584
rect 23293 18575 23351 18581
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 23676 18612 23704 18652
rect 23750 18640 23756 18692
rect 23808 18680 23814 18692
rect 24581 18683 24639 18689
rect 24581 18680 24593 18683
rect 23808 18652 24593 18680
rect 23808 18640 23814 18652
rect 24581 18649 24593 18652
rect 24627 18649 24639 18683
rect 25498 18680 25504 18692
rect 25459 18652 25504 18680
rect 24581 18643 24639 18649
rect 25498 18640 25504 18652
rect 25556 18640 25562 18692
rect 25593 18683 25651 18689
rect 25593 18649 25605 18683
rect 25639 18649 25651 18683
rect 25792 18680 25820 18788
rect 26237 18785 26249 18819
rect 26283 18816 26295 18819
rect 26694 18816 26700 18828
rect 26283 18788 26700 18816
rect 26283 18785 26295 18788
rect 26237 18779 26295 18785
rect 26694 18776 26700 18788
rect 26752 18776 26758 18828
rect 26329 18683 26387 18689
rect 26329 18680 26341 18683
rect 25792 18652 26341 18680
rect 25593 18643 25651 18649
rect 26329 18649 26341 18652
rect 26375 18649 26387 18683
rect 26329 18643 26387 18649
rect 25608 18612 25636 18643
rect 23676 18584 25636 18612
rect 25682 18572 25688 18624
rect 25740 18612 25746 18624
rect 27341 18615 27399 18621
rect 27341 18612 27353 18615
rect 25740 18584 27353 18612
rect 25740 18572 25746 18584
rect 27341 18581 27353 18584
rect 27387 18581 27399 18615
rect 27341 18575 27399 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 15838 18408 15844 18420
rect 15799 18380 15844 18408
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 19702 18408 19708 18420
rect 19306 18380 19708 18408
rect 1857 18343 1915 18349
rect 1857 18309 1869 18343
rect 1903 18340 1915 18343
rect 1903 18312 12434 18340
rect 1903 18309 1915 18312
rect 1857 18303 1915 18309
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1673 18275 1731 18281
rect 1673 18272 1685 18275
rect 1636 18244 1685 18272
rect 1636 18232 1642 18244
rect 1673 18241 1685 18244
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 2004 18244 9689 18272
rect 2004 18232 2010 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 12406 18204 12434 18312
rect 17678 18300 17684 18352
rect 17736 18340 17742 18352
rect 19306 18340 19334 18380
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 20530 18368 20536 18420
rect 20588 18408 20594 18420
rect 20717 18411 20775 18417
rect 20717 18408 20729 18411
rect 20588 18380 20729 18408
rect 20588 18368 20594 18380
rect 20717 18377 20729 18380
rect 20763 18377 20775 18411
rect 20717 18371 20775 18377
rect 22097 18411 22155 18417
rect 22097 18377 22109 18411
rect 22143 18408 22155 18411
rect 22186 18408 22192 18420
rect 22143 18380 22192 18408
rect 22143 18377 22155 18380
rect 22097 18371 22155 18377
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 25774 18408 25780 18420
rect 22848 18380 25780 18408
rect 17736 18312 19334 18340
rect 17736 18300 17742 18312
rect 19518 18300 19524 18352
rect 19576 18340 19582 18352
rect 22848 18349 22876 18380
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 37553 18411 37611 18417
rect 37553 18377 37565 18411
rect 37599 18408 37611 18411
rect 38010 18408 38016 18420
rect 37599 18380 38016 18408
rect 37599 18377 37611 18380
rect 37553 18371 37611 18377
rect 38010 18368 38016 18380
rect 38068 18368 38074 18420
rect 19613 18343 19671 18349
rect 19613 18340 19625 18343
rect 19576 18312 19625 18340
rect 19576 18300 19582 18312
rect 19613 18309 19625 18312
rect 19659 18309 19671 18343
rect 22833 18343 22891 18349
rect 19613 18303 19671 18309
rect 20824 18312 22600 18340
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15470 18272 15476 18284
rect 15243 18244 15476 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 15470 18232 15476 18244
rect 15528 18272 15534 18284
rect 20824 18281 20852 18312
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15528 18244 15761 18272
rect 15528 18232 15534 18244
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 21358 18272 21364 18284
rect 21315 18244 21364 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 22020 18281 22048 18312
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18272 22063 18275
rect 22186 18272 22192 18284
rect 22051 18244 22192 18272
rect 22051 18241 22063 18244
rect 22005 18235 22063 18241
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 12406 18176 18368 18204
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 16482 18136 16488 18148
rect 9815 18108 16488 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 16482 18096 16488 18108
rect 16540 18096 16546 18148
rect 18340 18068 18368 18176
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 19392 18176 19533 18204
rect 19392 18164 19398 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 19521 18167 19579 18173
rect 19702 18164 19708 18216
rect 19760 18204 19766 18216
rect 19797 18207 19855 18213
rect 19797 18204 19809 18207
rect 19760 18176 19809 18204
rect 19760 18164 19766 18176
rect 19797 18173 19809 18176
rect 19843 18204 19855 18207
rect 22370 18204 22376 18216
rect 19843 18176 22376 18204
rect 19843 18173 19855 18176
rect 19797 18167 19855 18173
rect 22370 18164 22376 18176
rect 22428 18164 22434 18216
rect 18417 18139 18475 18145
rect 18417 18105 18429 18139
rect 18463 18136 18475 18139
rect 19978 18136 19984 18148
rect 18463 18108 19984 18136
rect 18463 18105 18475 18108
rect 18417 18099 18475 18105
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 21542 18136 21548 18148
rect 21284 18108 21548 18136
rect 21284 18068 21312 18108
rect 21542 18096 21548 18108
rect 21600 18096 21606 18148
rect 22572 18136 22600 18312
rect 22833 18309 22845 18343
rect 22879 18309 22891 18343
rect 23750 18340 23756 18352
rect 23711 18312 23756 18340
rect 22833 18303 22891 18309
rect 23750 18300 23756 18312
rect 23808 18300 23814 18352
rect 25590 18340 25596 18352
rect 25551 18312 25596 18340
rect 25590 18300 25596 18312
rect 25648 18300 25654 18352
rect 25682 18300 25688 18352
rect 25740 18340 25746 18352
rect 27154 18340 27160 18352
rect 25740 18312 25785 18340
rect 27115 18312 27160 18340
rect 25740 18300 25746 18312
rect 27154 18300 27160 18312
rect 27212 18300 27218 18352
rect 27522 18300 27528 18352
rect 27580 18340 27586 18352
rect 27709 18343 27767 18349
rect 27709 18340 27721 18343
rect 27580 18312 27721 18340
rect 27580 18300 27586 18312
rect 27709 18309 27721 18312
rect 27755 18309 27767 18343
rect 27709 18303 27767 18309
rect 27798 18300 27804 18352
rect 27856 18340 27862 18352
rect 27856 18312 27901 18340
rect 27856 18300 27862 18312
rect 24394 18272 24400 18284
rect 24355 18244 24400 18272
rect 24394 18232 24400 18244
rect 24452 18232 24458 18284
rect 26237 18275 26295 18281
rect 26237 18272 26249 18275
rect 26068 18244 26249 18272
rect 22738 18204 22744 18216
rect 22699 18176 22744 18204
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 24912 18176 25053 18204
rect 24912 18164 24918 18176
rect 25041 18173 25053 18176
rect 25087 18173 25099 18207
rect 25041 18167 25099 18173
rect 23198 18136 23204 18148
rect 22572 18108 23204 18136
rect 23198 18096 23204 18108
rect 23256 18096 23262 18148
rect 23658 18096 23664 18148
rect 23716 18136 23722 18148
rect 26068 18136 26096 18244
rect 26237 18241 26249 18244
rect 26283 18241 26295 18275
rect 26237 18235 26295 18241
rect 28902 18232 28908 18284
rect 28960 18272 28966 18284
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 28960 18244 37473 18272
rect 28960 18232 28966 18244
rect 37461 18241 37473 18244
rect 37507 18241 37519 18275
rect 37461 18235 37519 18241
rect 26602 18136 26608 18148
rect 23716 18108 26096 18136
rect 26160 18108 26608 18136
rect 23716 18096 23722 18108
rect 18340 18040 21312 18068
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 22462 18068 22468 18080
rect 21407 18040 22468 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 23750 18028 23756 18080
rect 23808 18068 23814 18080
rect 24305 18071 24363 18077
rect 24305 18068 24317 18071
rect 23808 18040 24317 18068
rect 23808 18028 23814 18040
rect 24305 18037 24317 18040
rect 24351 18037 24363 18071
rect 24305 18031 24363 18037
rect 24394 18028 24400 18080
rect 24452 18068 24458 18080
rect 26160 18068 26188 18108
rect 26602 18096 26608 18108
rect 26660 18136 26666 18148
rect 28353 18139 28411 18145
rect 28353 18136 28365 18139
rect 26660 18108 28365 18136
rect 26660 18096 26666 18108
rect 28353 18105 28365 18108
rect 28399 18105 28411 18139
rect 28353 18099 28411 18105
rect 26326 18068 26332 18080
rect 24452 18040 26188 18068
rect 26287 18040 26332 18068
rect 24452 18028 24458 18040
rect 26326 18028 26332 18040
rect 26384 18028 26390 18080
rect 28368 18068 28396 18099
rect 28994 18068 29000 18080
rect 28368 18040 29000 18068
rect 28994 18028 29000 18040
rect 29052 18028 29058 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 20898 17824 20904 17876
rect 20956 17864 20962 17876
rect 20956 17836 22784 17864
rect 20956 17824 20962 17836
rect 22756 17808 22784 17836
rect 23290 17824 23296 17876
rect 23348 17864 23354 17876
rect 25958 17864 25964 17876
rect 23348 17836 25964 17864
rect 23348 17824 23354 17836
rect 25958 17824 25964 17836
rect 26016 17824 26022 17876
rect 26050 17824 26056 17876
rect 26108 17864 26114 17876
rect 26513 17867 26571 17873
rect 26513 17864 26525 17867
rect 26108 17836 26525 17864
rect 26108 17824 26114 17836
rect 26513 17833 26525 17836
rect 26559 17833 26571 17867
rect 26513 17827 26571 17833
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 19150 17796 19156 17808
rect 17972 17768 19156 17796
rect 17972 17669 18000 17768
rect 19150 17756 19156 17768
rect 19208 17756 19214 17808
rect 20257 17799 20315 17805
rect 20257 17765 20269 17799
rect 20303 17796 20315 17799
rect 21726 17796 21732 17808
rect 20303 17768 21732 17796
rect 20303 17765 20315 17768
rect 20257 17759 20315 17765
rect 21726 17756 21732 17768
rect 21784 17756 21790 17808
rect 21821 17799 21879 17805
rect 21821 17765 21833 17799
rect 21867 17796 21879 17799
rect 22186 17796 22192 17808
rect 21867 17768 22192 17796
rect 21867 17765 21879 17768
rect 21821 17759 21879 17765
rect 22186 17756 22192 17768
rect 22244 17756 22250 17808
rect 22738 17756 22744 17808
rect 22796 17796 22802 17808
rect 22925 17799 22983 17805
rect 22925 17796 22937 17799
rect 22796 17768 22937 17796
rect 22796 17756 22802 17768
rect 22925 17765 22937 17768
rect 22971 17765 22983 17799
rect 22925 17759 22983 17765
rect 24762 17756 24768 17808
rect 24820 17796 24826 17808
rect 25317 17799 25375 17805
rect 25317 17796 25329 17799
rect 24820 17768 25329 17796
rect 24820 17756 24826 17768
rect 25317 17765 25329 17768
rect 25363 17765 25375 17799
rect 27798 17796 27804 17808
rect 25317 17759 25375 17765
rect 25884 17768 27804 17796
rect 21358 17728 21364 17740
rect 18800 17700 21364 17728
rect 18800 17669 18828 17700
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 25884 17737 25912 17768
rect 26528 17740 26556 17768
rect 27798 17756 27804 17768
rect 27856 17756 27862 17808
rect 25869 17731 25927 17737
rect 25869 17697 25881 17731
rect 25915 17697 25927 17731
rect 25869 17691 25927 17697
rect 26510 17688 26516 17740
rect 26568 17688 26574 17740
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 19521 17663 19579 17669
rect 19521 17660 19533 17663
rect 19208 17632 19533 17660
rect 19208 17620 19214 17632
rect 19521 17629 19533 17632
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 19978 17620 19984 17672
rect 20036 17660 20042 17672
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 20036 17632 20177 17660
rect 20036 17620 20042 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 21082 17660 21088 17672
rect 21043 17632 21088 17660
rect 20165 17623 20223 17629
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 23658 17660 23664 17672
rect 23571 17632 23664 17660
rect 23658 17620 23664 17632
rect 23716 17660 23722 17672
rect 23934 17660 23940 17672
rect 23716 17632 23940 17660
rect 23716 17620 23722 17632
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 24302 17620 24308 17672
rect 24360 17660 24366 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 24360 17632 24593 17660
rect 24360 17620 24366 17632
rect 24581 17629 24593 17632
rect 24627 17629 24639 17663
rect 26602 17660 26608 17672
rect 26563 17632 26608 17660
rect 24581 17623 24639 17629
rect 26602 17620 26608 17632
rect 26660 17620 26666 17672
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 27249 17663 27307 17669
rect 27249 17660 27261 17663
rect 26936 17632 27261 17660
rect 26936 17620 26942 17632
rect 27249 17629 27261 17632
rect 27295 17660 27307 17663
rect 27893 17663 27951 17669
rect 27893 17660 27905 17663
rect 27295 17632 27905 17660
rect 27295 17629 27307 17632
rect 27249 17623 27307 17629
rect 27893 17629 27905 17632
rect 27939 17629 27951 17663
rect 28350 17660 28356 17672
rect 28311 17632 28356 17660
rect 27893 17623 27951 17629
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17592 18107 17595
rect 19426 17592 19432 17604
rect 18095 17564 19432 17592
rect 18095 17561 18107 17564
rect 18049 17555 18107 17561
rect 19426 17552 19432 17564
rect 19484 17552 19490 17604
rect 19613 17595 19671 17601
rect 19613 17561 19625 17595
rect 19659 17592 19671 17595
rect 20990 17592 20996 17604
rect 19659 17564 20996 17592
rect 19659 17561 19671 17564
rect 19613 17555 19671 17561
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 22370 17592 22376 17604
rect 22331 17564 22376 17592
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 22465 17595 22523 17601
rect 22465 17561 22477 17595
rect 22511 17561 22523 17595
rect 22465 17555 22523 17561
rect 25777 17595 25835 17601
rect 25777 17561 25789 17595
rect 25823 17561 25835 17595
rect 25777 17555 25835 17561
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 18564 17496 18705 17524
rect 18564 17484 18570 17496
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 18693 17487 18751 17493
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 22480 17524 22508 17555
rect 23569 17527 23627 17533
rect 23569 17524 23581 17527
rect 22480 17496 23581 17524
rect 23569 17493 23581 17496
rect 23615 17493 23627 17527
rect 23569 17487 23627 17493
rect 24673 17527 24731 17533
rect 24673 17493 24685 17527
rect 24719 17524 24731 17527
rect 24946 17524 24952 17536
rect 24719 17496 24952 17524
rect 24719 17493 24731 17496
rect 24673 17487 24731 17493
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 25792 17524 25820 17555
rect 26234 17552 26240 17604
rect 26292 17592 26298 17604
rect 27157 17595 27215 17601
rect 27157 17592 27169 17595
rect 26292 17564 27169 17592
rect 26292 17552 26298 17564
rect 27157 17561 27169 17564
rect 27203 17561 27215 17595
rect 27157 17555 27215 17561
rect 26326 17524 26332 17536
rect 25792 17496 26332 17524
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 27614 17484 27620 17536
rect 27672 17524 27678 17536
rect 27801 17527 27859 17533
rect 27801 17524 27813 17527
rect 27672 17496 27813 17524
rect 27672 17484 27678 17496
rect 27801 17493 27813 17496
rect 27847 17493 27859 17527
rect 28442 17524 28448 17536
rect 28403 17496 28448 17524
rect 27801 17487 27859 17493
rect 28442 17484 28448 17496
rect 28500 17484 28506 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 18690 17320 18696 17332
rect 17512 17292 18696 17320
rect 17402 17252 17408 17264
rect 17363 17224 17408 17252
rect 17402 17212 17408 17224
rect 17460 17212 17466 17264
rect 17512 17261 17540 17292
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 23290 17320 23296 17332
rect 21008 17292 23296 17320
rect 17497 17255 17555 17261
rect 17497 17221 17509 17255
rect 17543 17221 17555 17255
rect 18506 17252 18512 17264
rect 18467 17224 18512 17252
rect 17497 17215 17555 17221
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 19061 17255 19119 17261
rect 19061 17221 19073 17255
rect 19107 17252 19119 17255
rect 20898 17252 20904 17264
rect 19107 17224 20904 17252
rect 19107 17221 19119 17224
rect 19061 17215 19119 17221
rect 20898 17212 20904 17224
rect 20956 17212 20962 17264
rect 20254 17184 20260 17196
rect 20215 17156 20260 17184
rect 20254 17144 20260 17156
rect 20312 17184 20318 17196
rect 21008 17184 21036 17292
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 26329 17323 26387 17329
rect 26329 17320 26341 17323
rect 23532 17292 26341 17320
rect 23532 17280 23538 17292
rect 26329 17289 26341 17292
rect 26375 17289 26387 17323
rect 26329 17283 26387 17289
rect 21174 17212 21180 17264
rect 21232 17252 21238 17264
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 21232 17224 22201 17252
rect 21232 17212 21238 17224
rect 22189 17221 22201 17224
rect 22235 17221 22247 17255
rect 23750 17252 23756 17264
rect 23711 17224 23756 17252
rect 22189 17215 22247 17221
rect 23750 17212 23756 17224
rect 23808 17212 23814 17264
rect 24946 17252 24952 17264
rect 24907 17224 24952 17252
rect 24946 17212 24952 17224
rect 25004 17212 25010 17264
rect 25038 17212 25044 17264
rect 25096 17252 25102 17264
rect 25682 17252 25688 17264
rect 25096 17224 25688 17252
rect 25096 17212 25102 17224
rect 25682 17212 25688 17224
rect 25740 17212 25746 17264
rect 26050 17212 26056 17264
rect 26108 17252 26114 17264
rect 26108 17224 27384 17252
rect 26108 17212 26114 17224
rect 20312 17156 21036 17184
rect 20312 17144 20318 17156
rect 21082 17144 21088 17196
rect 21140 17184 21146 17196
rect 25590 17184 25596 17196
rect 21140 17156 21185 17184
rect 25551 17156 25596 17184
rect 21140 17144 21146 17156
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 25958 17144 25964 17196
rect 26016 17184 26022 17196
rect 26421 17187 26479 17193
rect 26421 17184 26433 17187
rect 26016 17156 26433 17184
rect 26016 17144 26022 17156
rect 26421 17153 26433 17156
rect 26467 17184 26479 17187
rect 27154 17184 27160 17196
rect 26467 17156 27160 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 27154 17144 27160 17156
rect 27212 17144 27218 17196
rect 27356 17193 27384 17224
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17153 27399 17187
rect 27982 17184 27988 17196
rect 27943 17156 27988 17184
rect 27341 17147 27399 17153
rect 27982 17144 27988 17156
rect 28040 17184 28046 17196
rect 28997 17187 29055 17193
rect 28997 17184 29009 17187
rect 28040 17156 29009 17184
rect 28040 17144 28046 17156
rect 28997 17153 29009 17156
rect 29043 17153 29055 17187
rect 28997 17147 29055 17153
rect 37553 17187 37611 17193
rect 37553 17153 37565 17187
rect 37599 17184 37611 17187
rect 38194 17184 38200 17196
rect 37599 17156 38200 17184
rect 37599 17153 37611 17156
rect 37553 17147 37611 17153
rect 38194 17144 38200 17156
rect 38252 17144 38258 17196
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17116 17279 17119
rect 17862 17116 17868 17128
rect 17267 17088 17868 17116
rect 17267 17085 17279 17088
rect 17221 17079 17279 17085
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 18414 17116 18420 17128
rect 18375 17088 18420 17116
rect 18414 17076 18420 17088
rect 18472 17076 18478 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 22097 17119 22155 17125
rect 22097 17116 22109 17119
rect 19392 17088 22109 17116
rect 19392 17076 19398 17088
rect 22097 17085 22109 17088
rect 22143 17085 22155 17119
rect 23201 17119 23259 17125
rect 23201 17116 23213 17119
rect 22097 17079 22155 17085
rect 22572 17088 23213 17116
rect 15286 17008 15292 17060
rect 15344 17048 15350 17060
rect 22572 17048 22600 17088
rect 23201 17085 23213 17088
rect 23247 17085 23259 17119
rect 23201 17079 23259 17085
rect 23566 17076 23572 17128
rect 23624 17116 23630 17128
rect 23845 17119 23903 17125
rect 23845 17116 23857 17119
rect 23624 17088 23857 17116
rect 23624 17076 23630 17088
rect 23845 17085 23857 17088
rect 23891 17085 23903 17119
rect 24854 17116 24860 17128
rect 23845 17079 23903 17085
rect 24412 17088 24860 17116
rect 15344 17020 22600 17048
rect 22649 17051 22707 17057
rect 15344 17008 15350 17020
rect 22649 17017 22661 17051
rect 22695 17048 22707 17051
rect 24412 17048 24440 17088
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 25498 17076 25504 17128
rect 25556 17116 25562 17128
rect 27249 17119 27307 17125
rect 27249 17116 27261 17119
rect 25556 17088 27261 17116
rect 25556 17076 25562 17088
rect 27249 17085 27261 17088
rect 27295 17085 27307 17119
rect 27249 17079 27307 17085
rect 22695 17020 24440 17048
rect 24489 17051 24547 17057
rect 22695 17017 22707 17020
rect 22649 17011 22707 17017
rect 24489 17017 24501 17051
rect 24535 17017 24547 17051
rect 24872 17048 24900 17076
rect 24872 17020 26372 17048
rect 24489 17011 24547 17017
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 20254 16980 20260 16992
rect 19843 16952 20260 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20622 16980 20628 16992
rect 20395 16952 20628 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 20993 16983 21051 16989
rect 20993 16949 21005 16983
rect 21039 16980 21051 16983
rect 21910 16980 21916 16992
rect 21039 16952 21916 16980
rect 21039 16949 21051 16952
rect 20993 16943 21051 16949
rect 21910 16940 21916 16952
rect 21968 16940 21974 16992
rect 22002 16940 22008 16992
rect 22060 16980 22066 16992
rect 24504 16980 24532 17011
rect 22060 16952 24532 16980
rect 22060 16940 22066 16952
rect 25130 16940 25136 16992
rect 25188 16980 25194 16992
rect 25685 16983 25743 16989
rect 25685 16980 25697 16983
rect 25188 16952 25697 16980
rect 25188 16940 25194 16952
rect 25685 16949 25697 16952
rect 25731 16949 25743 16983
rect 26344 16980 26372 17020
rect 26418 17008 26424 17060
rect 26476 17048 26482 17060
rect 27893 17051 27951 17057
rect 27893 17048 27905 17051
rect 26476 17020 27905 17048
rect 26476 17008 26482 17020
rect 27893 17017 27905 17020
rect 27939 17017 27951 17051
rect 38010 17048 38016 17060
rect 37971 17020 38016 17048
rect 27893 17011 27951 17017
rect 38010 17008 38016 17020
rect 38068 17008 38074 17060
rect 27062 16980 27068 16992
rect 26344 16952 27068 16980
rect 25685 16943 25743 16949
rect 27062 16940 27068 16952
rect 27120 16940 27126 16992
rect 27154 16940 27160 16992
rect 27212 16980 27218 16992
rect 28537 16983 28595 16989
rect 28537 16980 28549 16983
rect 27212 16952 28549 16980
rect 27212 16940 27218 16952
rect 28537 16949 28549 16952
rect 28583 16980 28595 16983
rect 29270 16980 29276 16992
rect 28583 16952 29276 16980
rect 28583 16949 28595 16952
rect 28537 16943 28595 16949
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 17494 16776 17500 16788
rect 17455 16748 17500 16776
rect 17494 16736 17500 16748
rect 17552 16776 17558 16788
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 17552 16748 18061 16776
rect 17552 16736 17558 16748
rect 18049 16745 18061 16748
rect 18095 16745 18107 16779
rect 22738 16776 22744 16788
rect 18049 16739 18107 16745
rect 22296 16748 22744 16776
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 12952 16612 13645 16640
rect 12952 16600 12958 16612
rect 13004 16581 13032 16612
rect 13633 16609 13645 16612
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 14642 16600 14648 16652
rect 14700 16640 14706 16652
rect 15933 16643 15991 16649
rect 15933 16640 15945 16643
rect 14700 16612 15945 16640
rect 14700 16600 14706 16612
rect 15304 16581 15332 16612
rect 15933 16609 15945 16612
rect 15979 16609 15991 16643
rect 18064 16640 18092 16739
rect 20438 16668 20444 16720
rect 20496 16708 20502 16720
rect 20496 16680 20576 16708
rect 20496 16668 20502 16680
rect 20548 16649 20576 16680
rect 21082 16668 21088 16720
rect 21140 16708 21146 16720
rect 22002 16708 22008 16720
rect 21140 16680 22008 16708
rect 21140 16668 21146 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 20533 16643 20591 16649
rect 18064 16612 18828 16640
rect 15933 16603 15991 16609
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 12989 16575 13047 16581
rect 3099 16544 4108 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 2866 16436 2872 16448
rect 2827 16408 2872 16436
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 4080 16445 4108 16544
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16572 15439 16575
rect 17402 16572 17408 16584
rect 15427 16544 17408 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 18690 16572 18696 16584
rect 18651 16544 18696 16572
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 18800 16581 18828 16612
rect 20533 16609 20545 16643
rect 20579 16609 20591 16643
rect 21174 16640 21180 16652
rect 21135 16612 21180 16640
rect 20533 16603 20591 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 22296 16640 22324 16748
rect 22738 16736 22744 16748
rect 22796 16776 22802 16788
rect 22796 16748 23060 16776
rect 22796 16736 22802 16748
rect 22646 16668 22652 16720
rect 22704 16708 22710 16720
rect 22925 16711 22983 16717
rect 22925 16708 22937 16711
rect 22704 16680 22937 16708
rect 22704 16668 22710 16680
rect 22925 16677 22937 16680
rect 22971 16677 22983 16711
rect 23032 16708 23060 16748
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 26050 16776 26056 16788
rect 24360 16748 26056 16776
rect 24360 16736 24366 16748
rect 26050 16736 26056 16748
rect 26108 16736 26114 16788
rect 26142 16736 26148 16788
rect 26200 16776 26206 16788
rect 26200 16748 26924 16776
rect 26200 16736 26206 16748
rect 25590 16708 25596 16720
rect 23032 16680 25596 16708
rect 22925 16671 22983 16677
rect 25590 16668 25596 16680
rect 25648 16668 25654 16720
rect 26326 16668 26332 16720
rect 26384 16708 26390 16720
rect 26421 16711 26479 16717
rect 26421 16708 26433 16711
rect 26384 16680 26433 16708
rect 26384 16668 26390 16680
rect 26421 16677 26433 16680
rect 26467 16677 26479 16711
rect 26421 16671 26479 16677
rect 21416 16612 22324 16640
rect 22373 16643 22431 16649
rect 21416 16600 21422 16612
rect 22373 16609 22385 16643
rect 22419 16640 22431 16643
rect 23658 16640 23664 16652
rect 22419 16612 23664 16640
rect 22419 16609 22431 16612
rect 22373 16603 22431 16609
rect 23658 16600 23664 16612
rect 23716 16600 23722 16652
rect 24762 16640 24768 16652
rect 24723 16612 24768 16640
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 25222 16640 25228 16652
rect 25135 16612 25228 16640
rect 25222 16600 25228 16612
rect 25280 16640 25286 16652
rect 25280 16612 26556 16640
rect 25280 16600 25286 16612
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16572 18843 16575
rect 19242 16572 19248 16584
rect 18831 16544 19248 16572
rect 18831 16541 18843 16544
rect 18785 16535 18843 16541
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20070 16572 20076 16584
rect 19843 16544 20076 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 20070 16532 20076 16544
rect 20128 16532 20134 16584
rect 26528 16572 26556 16612
rect 26896 16574 26924 16748
rect 27816 16680 28856 16708
rect 27816 16581 27844 16680
rect 28828 16652 28856 16680
rect 28350 16640 28356 16652
rect 28311 16612 28356 16640
rect 28350 16600 28356 16612
rect 28408 16600 28414 16652
rect 28810 16640 28816 16652
rect 28771 16612 28816 16640
rect 28810 16600 28816 16612
rect 28868 16600 28874 16652
rect 26973 16575 27031 16581
rect 26973 16574 26985 16575
rect 26528 16544 26740 16572
rect 26896 16546 26985 16574
rect 13081 16507 13139 16513
rect 13081 16473 13093 16507
rect 13127 16504 13139 16507
rect 19334 16504 19340 16516
rect 13127 16476 19340 16504
rect 13127 16473 13139 16476
rect 13081 16467 13139 16473
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 20622 16464 20628 16516
rect 20680 16504 20686 16516
rect 21726 16504 21732 16516
rect 20680 16476 20725 16504
rect 21687 16476 21732 16504
rect 20680 16464 20686 16476
rect 21726 16464 21732 16476
rect 21784 16464 21790 16516
rect 21821 16507 21879 16513
rect 21821 16473 21833 16507
rect 21867 16504 21879 16507
rect 22370 16504 22376 16516
rect 21867 16476 22376 16504
rect 21867 16473 21879 16476
rect 21821 16467 21879 16473
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 23382 16504 23388 16516
rect 23343 16476 23388 16504
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 23477 16507 23535 16513
rect 23477 16473 23489 16507
rect 23523 16504 23535 16507
rect 24946 16504 24952 16516
rect 23523 16476 24952 16504
rect 23523 16473 23535 16476
rect 23477 16467 23535 16473
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 25130 16504 25136 16516
rect 25091 16476 25136 16504
rect 25130 16464 25136 16476
rect 25188 16464 25194 16516
rect 25682 16464 25688 16516
rect 25740 16504 25746 16516
rect 25869 16507 25927 16513
rect 25869 16504 25881 16507
rect 25740 16476 25881 16504
rect 25740 16464 25746 16476
rect 25869 16473 25881 16476
rect 25915 16473 25927 16507
rect 25869 16467 25927 16473
rect 25961 16507 26019 16513
rect 25961 16473 25973 16507
rect 26007 16504 26019 16507
rect 26602 16504 26608 16516
rect 26007 16476 26608 16504
rect 26007 16473 26019 16476
rect 25961 16467 26019 16473
rect 26602 16464 26608 16476
rect 26660 16464 26666 16516
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16436 4123 16439
rect 4614 16436 4620 16448
rect 4111 16408 4620 16436
rect 4111 16405 4123 16408
rect 4065 16399 4123 16405
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 15746 16396 15752 16448
rect 15804 16436 15810 16448
rect 17037 16439 17095 16445
rect 17037 16436 17049 16439
rect 15804 16408 17049 16436
rect 15804 16396 15810 16408
rect 17037 16405 17049 16408
rect 17083 16436 17095 16439
rect 18046 16436 18052 16448
rect 17083 16408 18052 16436
rect 17083 16405 17095 16408
rect 17037 16399 17095 16405
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 19889 16439 19947 16445
rect 19889 16405 19901 16439
rect 19935 16436 19947 16439
rect 21910 16436 21916 16448
rect 19935 16408 21916 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 21910 16396 21916 16408
rect 21968 16396 21974 16448
rect 26712 16436 26740 16544
rect 26973 16541 26985 16546
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 26786 16464 26792 16516
rect 26844 16504 26850 16516
rect 27614 16504 27620 16516
rect 26844 16476 27620 16504
rect 26844 16464 26850 16476
rect 27614 16464 27620 16476
rect 27672 16464 27678 16516
rect 27065 16439 27123 16445
rect 27065 16436 27077 16439
rect 26712 16408 27077 16436
rect 27065 16405 27077 16408
rect 27111 16405 27123 16439
rect 27065 16399 27123 16405
rect 27154 16396 27160 16448
rect 27212 16436 27218 16448
rect 27709 16439 27767 16445
rect 27709 16436 27721 16439
rect 27212 16408 27721 16436
rect 27212 16396 27218 16408
rect 27709 16405 27721 16408
rect 27755 16405 27767 16439
rect 27709 16399 27767 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 19981 16235 20039 16241
rect 19981 16232 19993 16235
rect 6886 16204 19993 16232
rect 2130 16124 2136 16176
rect 2188 16164 2194 16176
rect 6886 16164 6914 16204
rect 19981 16201 19993 16204
rect 20027 16201 20039 16235
rect 25498 16232 25504 16244
rect 19981 16195 20039 16201
rect 23768 16204 25504 16232
rect 15746 16164 15752 16176
rect 2188 16136 6914 16164
rect 15707 16136 15752 16164
rect 2188 16124 2194 16136
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 17221 16167 17279 16173
rect 17221 16164 17233 16167
rect 17184 16136 17233 16164
rect 17184 16124 17190 16136
rect 17221 16133 17233 16136
rect 17267 16133 17279 16167
rect 17221 16127 17279 16133
rect 18601 16167 18659 16173
rect 18601 16133 18613 16167
rect 18647 16164 18659 16167
rect 21177 16167 21235 16173
rect 21177 16164 21189 16167
rect 18647 16136 21189 16164
rect 18647 16133 18659 16136
rect 18601 16127 18659 16133
rect 21177 16133 21189 16136
rect 21223 16133 21235 16167
rect 21177 16127 21235 16133
rect 22182 16167 22240 16173
rect 22182 16133 22194 16167
rect 22228 16164 22240 16167
rect 22462 16164 22468 16176
rect 22228 16136 22468 16164
rect 22228 16133 22240 16136
rect 22182 16127 22240 16133
rect 22462 16124 22468 16136
rect 22520 16124 22526 16176
rect 23768 16173 23796 16204
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 23753 16167 23811 16173
rect 23753 16133 23765 16167
rect 23799 16133 23811 16167
rect 23753 16127 23811 16133
rect 23842 16124 23848 16176
rect 23900 16164 23906 16176
rect 24949 16167 25007 16173
rect 23900 16136 23945 16164
rect 23900 16124 23906 16136
rect 24949 16133 24961 16167
rect 24995 16164 25007 16167
rect 26234 16164 26240 16176
rect 24995 16136 26240 16164
rect 24995 16133 25007 16136
rect 24949 16127 25007 16133
rect 26234 16124 26240 16136
rect 26292 16124 26298 16176
rect 26418 16164 26424 16176
rect 26379 16136 26424 16164
rect 26418 16124 26424 16136
rect 26476 16124 26482 16176
rect 26510 16124 26516 16176
rect 26568 16164 26574 16176
rect 27341 16167 27399 16173
rect 26568 16136 26613 16164
rect 26568 16124 26574 16136
rect 27341 16133 27353 16167
rect 27387 16164 27399 16167
rect 28718 16164 28724 16176
rect 27387 16136 28724 16164
rect 27387 16133 27399 16136
rect 27341 16127 27399 16133
rect 28718 16124 28724 16136
rect 28776 16124 28782 16176
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 10594 16096 10600 16108
rect 1903 16068 10600 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16065 18567 16099
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 18509 16059 18567 16065
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 10560 16000 17141 16028
rect 10560 15988 10566 16000
rect 17129 15997 17141 16000
rect 17175 16028 17187 16031
rect 18414 16028 18420 16040
rect 17175 16000 18420 16028
rect 17175 15997 17187 16000
rect 17129 15991 17187 15997
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 16942 15920 16948 15972
rect 17000 15960 17006 15972
rect 17678 15960 17684 15972
rect 17000 15932 17684 15960
rect 17000 15920 17006 15932
rect 17678 15920 17684 15932
rect 17736 15920 17742 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16390 15892 16396 15904
rect 16347 15864 16396 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 18524 15892 18552 16059
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 20073 16099 20131 16105
rect 20073 16065 20085 16099
rect 20119 16096 20131 16099
rect 20622 16096 20628 16108
rect 20119 16068 20628 16096
rect 20119 16065 20131 16068
rect 20073 16059 20131 16065
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 28905 16099 28963 16105
rect 28905 16065 28917 16099
rect 28951 16096 28963 16099
rect 31386 16096 31392 16108
rect 28951 16068 31392 16096
rect 28951 16065 28963 16068
rect 28905 16059 28963 16065
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 37553 16099 37611 16105
rect 37553 16065 37565 16099
rect 37599 16096 37611 16099
rect 38194 16096 38200 16108
rect 37599 16068 38200 16096
rect 37599 16065 37611 16068
rect 37553 16059 37611 16065
rect 38194 16056 38200 16068
rect 38252 16056 38258 16108
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 16028 19487 16031
rect 21269 16031 21327 16037
rect 19475 16000 20852 16028
rect 19475 15997 19487 16000
rect 19429 15991 19487 15997
rect 18598 15920 18604 15972
rect 18656 15960 18662 15972
rect 20714 15960 20720 15972
rect 18656 15932 20720 15960
rect 18656 15920 18662 15932
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 20824 15960 20852 16000
rect 21269 15997 21281 16031
rect 21315 16028 21327 16031
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 21315 16000 22109 16028
rect 21315 15997 21327 16000
rect 21269 15991 21327 15997
rect 22097 15997 22109 16000
rect 22143 16028 22155 16031
rect 22186 16028 22192 16040
rect 22143 16000 22192 16028
rect 22143 15997 22155 16000
rect 22097 15991 22155 15997
rect 22186 15988 22192 16000
rect 22244 15988 22250 16040
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 23201 16031 23259 16037
rect 23201 16028 23213 16031
rect 23072 16000 23213 16028
rect 23072 15988 23078 16000
rect 23201 15997 23213 16000
rect 23247 15997 23259 16031
rect 23201 15991 23259 15997
rect 23658 15988 23664 16040
rect 23716 16028 23722 16040
rect 24762 16028 24768 16040
rect 23716 16000 24768 16028
rect 23716 15988 23722 16000
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 24946 15988 24952 16040
rect 25004 16028 25010 16040
rect 25041 16031 25099 16037
rect 25041 16028 25053 16031
rect 25004 16000 25053 16028
rect 25004 15988 25010 16000
rect 25041 15997 25053 16000
rect 25087 16028 25099 16031
rect 25406 16028 25412 16040
rect 25087 16000 25412 16028
rect 25087 15997 25099 16000
rect 25041 15991 25099 15997
rect 25406 15988 25412 16000
rect 25464 16028 25470 16040
rect 25464 16000 26096 16028
rect 25464 15988 25470 16000
rect 22646 15960 22652 15972
rect 20824 15932 22508 15960
rect 22607 15932 22652 15960
rect 22186 15892 22192 15904
rect 17276 15864 22192 15892
rect 17276 15852 17282 15864
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 22480 15892 22508 15932
rect 22646 15920 22652 15932
rect 22704 15920 22710 15972
rect 25498 15960 25504 15972
rect 22756 15932 25504 15960
rect 22756 15892 22784 15932
rect 25498 15920 25504 15932
rect 25556 15920 25562 15972
rect 25958 15960 25964 15972
rect 25919 15932 25964 15960
rect 25958 15920 25964 15932
rect 26016 15920 26022 15972
rect 26068 15960 26096 16000
rect 26234 15988 26240 16040
rect 26292 16028 26298 16040
rect 27062 16028 27068 16040
rect 26292 16000 27068 16028
rect 26292 15988 26298 16000
rect 27062 15988 27068 16000
rect 27120 16028 27126 16040
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 27120 16000 27261 16028
rect 27120 15988 27126 16000
rect 27249 15997 27261 16000
rect 27295 15997 27307 16031
rect 28074 16028 28080 16040
rect 28035 16000 28080 16028
rect 27249 15991 27307 15997
rect 28074 15988 28080 16000
rect 28132 15988 28138 16040
rect 29546 15960 29552 15972
rect 26068 15932 29552 15960
rect 29546 15920 29552 15932
rect 29604 15920 29610 15972
rect 22480 15864 22784 15892
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 26970 15892 26976 15904
rect 24820 15864 26976 15892
rect 24820 15852 24826 15864
rect 26970 15852 26976 15864
rect 27028 15852 27034 15904
rect 27614 15852 27620 15904
rect 27672 15892 27678 15904
rect 28813 15895 28871 15901
rect 28813 15892 28825 15895
rect 27672 15864 28825 15892
rect 27672 15852 27678 15864
rect 28813 15861 28825 15864
rect 28859 15861 28871 15895
rect 28813 15855 28871 15861
rect 28994 15852 29000 15904
rect 29052 15892 29058 15904
rect 29454 15892 29460 15904
rect 29052 15864 29460 15892
rect 29052 15852 29058 15864
rect 29454 15852 29460 15864
rect 29512 15852 29518 15904
rect 38102 15892 38108 15904
rect 38063 15864 38108 15892
rect 38102 15852 38108 15864
rect 38160 15852 38166 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 10502 15688 10508 15700
rect 10463 15660 10508 15688
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 17126 15688 17132 15700
rect 17087 15660 17132 15688
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 21634 15688 21640 15700
rect 18104 15660 21640 15688
rect 18104 15648 18110 15660
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 25682 15688 25688 15700
rect 25056 15660 25688 15688
rect 15378 15620 15384 15632
rect 15291 15592 15384 15620
rect 15378 15580 15384 15592
rect 15436 15620 15442 15632
rect 17310 15620 17316 15632
rect 15436 15592 17316 15620
rect 15436 15580 15442 15592
rect 17310 15580 17316 15592
rect 17368 15620 17374 15632
rect 17368 15592 22140 15620
rect 17368 15580 17374 15592
rect 17678 15552 17684 15564
rect 16408 15524 17684 15552
rect 16408 15496 16436 15524
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18187 15524 19380 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 4672 15456 10425 15484
rect 4672 15444 4678 15456
rect 10413 15453 10425 15456
rect 10459 15484 10471 15487
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10459 15456 11069 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 11057 15453 11069 15456
rect 11103 15453 11115 15487
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 11057 15447 11115 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 17218 15484 17224 15496
rect 17179 15456 17224 15484
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 18046 15484 18052 15496
rect 18007 15456 18052 15484
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15453 18935 15487
rect 19352 15484 19380 15524
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19889 15555 19947 15561
rect 19889 15552 19901 15555
rect 19484 15524 19901 15552
rect 19484 15512 19490 15524
rect 19889 15521 19901 15524
rect 19935 15521 19947 15555
rect 19889 15515 19947 15521
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 20438 15552 20444 15564
rect 20119 15524 20444 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 20990 15552 20996 15564
rect 20951 15524 20996 15552
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 21177 15555 21235 15561
rect 21177 15521 21189 15555
rect 21223 15552 21235 15555
rect 21450 15552 21456 15564
rect 21223 15524 21456 15552
rect 21223 15521 21235 15524
rect 21177 15515 21235 15521
rect 21450 15512 21456 15524
rect 21508 15512 21514 15564
rect 22112 15552 22140 15592
rect 22186 15580 22192 15632
rect 22244 15620 22250 15632
rect 25056 15620 25084 15660
rect 25682 15648 25688 15660
rect 25740 15648 25746 15700
rect 25774 15648 25780 15700
rect 25832 15688 25838 15700
rect 25869 15691 25927 15697
rect 25869 15688 25881 15691
rect 25832 15660 25881 15688
rect 25832 15648 25838 15660
rect 25869 15657 25881 15660
rect 25915 15657 25927 15691
rect 25869 15651 25927 15657
rect 26050 15648 26056 15700
rect 26108 15688 26114 15700
rect 29733 15691 29791 15697
rect 29733 15688 29745 15691
rect 26108 15660 29745 15688
rect 26108 15648 26114 15660
rect 29733 15657 29745 15660
rect 29779 15688 29791 15691
rect 36814 15688 36820 15700
rect 29779 15660 36820 15688
rect 29779 15657 29791 15660
rect 29733 15651 29791 15657
rect 36814 15648 36820 15660
rect 36872 15648 36878 15700
rect 22244 15592 25084 15620
rect 25148 15592 25452 15620
rect 22244 15580 22250 15592
rect 25148 15552 25176 15592
rect 22112 15524 25176 15552
rect 25222 15512 25228 15564
rect 25280 15552 25286 15564
rect 25424 15552 25452 15592
rect 25590 15580 25596 15632
rect 25648 15620 25654 15632
rect 29089 15623 29147 15629
rect 29089 15620 29101 15623
rect 25648 15592 29101 15620
rect 25648 15580 25654 15592
rect 29089 15589 29101 15592
rect 29135 15589 29147 15623
rect 29089 15583 29147 15589
rect 38102 15552 38108 15564
rect 25280 15524 25325 15552
rect 25424 15524 38108 15552
rect 25280 15512 25286 15524
rect 38102 15512 38108 15524
rect 38160 15512 38166 15564
rect 21358 15484 21364 15496
rect 19352 15456 21364 15484
rect 18877 15447 18935 15453
rect 15933 15419 15991 15425
rect 15933 15385 15945 15419
rect 15979 15416 15991 15419
rect 18892 15416 18920 15447
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 25774 15444 25780 15496
rect 25832 15484 25838 15496
rect 25961 15487 26019 15493
rect 25961 15484 25973 15487
rect 25832 15456 25973 15484
rect 25832 15444 25838 15456
rect 25961 15453 25973 15456
rect 26007 15484 26019 15487
rect 26050 15484 26056 15496
rect 26007 15456 26056 15484
rect 26007 15453 26019 15456
rect 25961 15447 26019 15453
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 28629 15487 28687 15493
rect 27908 15456 28580 15484
rect 21726 15416 21732 15428
rect 15979 15388 20668 15416
rect 21687 15388 21732 15416
rect 15979 15385 15991 15388
rect 15933 15379 15991 15385
rect 14826 15348 14832 15360
rect 14787 15320 14832 15348
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 16485 15351 16543 15357
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16666 15348 16672 15360
rect 16531 15320 16672 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 18564 15320 18797 15348
rect 18564 15308 18570 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 19150 15308 19156 15360
rect 19208 15348 19214 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 19208 15320 19441 15348
rect 19208 15308 19214 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 20530 15348 20536 15360
rect 20491 15320 20536 15348
rect 19429 15311 19487 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 20640 15348 20668 15388
rect 21726 15376 21732 15388
rect 21784 15376 21790 15428
rect 21821 15419 21879 15425
rect 21821 15385 21833 15419
rect 21867 15416 21879 15419
rect 21910 15416 21916 15428
rect 21867 15388 21916 15416
rect 21867 15385 21879 15388
rect 21821 15379 21879 15385
rect 21910 15376 21916 15388
rect 21968 15376 21974 15428
rect 22373 15419 22431 15425
rect 22373 15385 22385 15419
rect 22419 15385 22431 15419
rect 22373 15379 22431 15385
rect 22278 15348 22284 15360
rect 20640 15320 22284 15348
rect 22278 15308 22284 15320
rect 22336 15308 22342 15360
rect 22388 15348 22416 15379
rect 22830 15376 22836 15428
rect 22888 15416 22894 15428
rect 23385 15419 23443 15425
rect 23385 15416 23397 15419
rect 22888 15388 23397 15416
rect 22888 15376 22894 15388
rect 23385 15385 23397 15388
rect 23431 15385 23443 15419
rect 23385 15379 23443 15385
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 24029 15419 24087 15425
rect 23532 15388 23577 15416
rect 23532 15376 23538 15388
rect 24029 15385 24041 15419
rect 24075 15416 24087 15419
rect 24486 15416 24492 15428
rect 24075 15388 24492 15416
rect 24075 15385 24087 15388
rect 24029 15379 24087 15385
rect 24486 15376 24492 15388
rect 24544 15376 24550 15428
rect 24581 15419 24639 15425
rect 24581 15385 24593 15419
rect 24627 15385 24639 15419
rect 24581 15379 24639 15385
rect 25140 15419 25198 15425
rect 25140 15385 25152 15419
rect 25186 15385 25198 15419
rect 26970 15416 26976 15428
rect 25140 15379 25198 15385
rect 25332 15388 26832 15416
rect 26931 15388 26976 15416
rect 23566 15348 23572 15360
rect 22388 15320 23572 15348
rect 23566 15308 23572 15320
rect 23624 15348 23630 15360
rect 24596 15348 24624 15379
rect 23624 15320 24624 15348
rect 25148 15348 25176 15379
rect 25332 15348 25360 15388
rect 25148 15320 25360 15348
rect 23624 15308 23630 15320
rect 25682 15308 25688 15360
rect 25740 15348 25746 15360
rect 26694 15348 26700 15360
rect 25740 15320 26700 15348
rect 25740 15308 25746 15320
rect 26694 15308 26700 15320
rect 26752 15308 26758 15360
rect 26804 15348 26832 15388
rect 26970 15376 26976 15388
rect 27028 15376 27034 15428
rect 27065 15419 27123 15425
rect 27065 15385 27077 15419
rect 27111 15416 27123 15419
rect 27908 15416 27936 15456
rect 27111 15388 27936 15416
rect 27985 15419 28043 15425
rect 27111 15385 27123 15388
rect 27065 15379 27123 15385
rect 27985 15385 27997 15419
rect 28031 15416 28043 15419
rect 28074 15416 28080 15428
rect 28031 15388 28080 15416
rect 28031 15385 28043 15388
rect 27985 15379 28043 15385
rect 28074 15376 28080 15388
rect 28132 15376 28138 15428
rect 28552 15416 28580 15456
rect 28629 15453 28641 15487
rect 28675 15484 28687 15487
rect 29730 15484 29736 15496
rect 28675 15456 29736 15484
rect 28675 15453 28687 15456
rect 28629 15447 28687 15453
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 30190 15416 30196 15428
rect 28552 15388 30196 15416
rect 30190 15376 30196 15388
rect 30248 15376 30254 15428
rect 28537 15351 28595 15357
rect 28537 15348 28549 15351
rect 26804 15320 28549 15348
rect 28537 15317 28549 15320
rect 28583 15317 28595 15351
rect 30374 15348 30380 15360
rect 30335 15320 30380 15348
rect 28537 15311 28595 15317
rect 30374 15308 30380 15320
rect 30432 15348 30438 15360
rect 31294 15348 31300 15360
rect 30432 15320 31300 15348
rect 30432 15308 30438 15320
rect 31294 15308 31300 15320
rect 31352 15308 31358 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 15657 15147 15715 15153
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 15703 15116 19656 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 13630 15036 13636 15088
rect 13688 15076 13694 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 13688 15048 15884 15076
rect 13688 15036 13694 15048
rect 14642 15008 14648 15020
rect 14108 14980 14648 15008
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 14108 14813 14136 14980
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 14737 14875 14795 14881
rect 14737 14841 14749 14875
rect 14783 14872 14795 14875
rect 15746 14872 15752 14884
rect 14783 14844 15752 14872
rect 14783 14841 14795 14844
rect 14737 14835 14795 14841
rect 15746 14832 15752 14844
rect 15804 14832 15810 14884
rect 15856 14872 15884 15048
rect 16776 15048 17049 15076
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16574 15008 16580 15020
rect 16347 14980 16580 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 16776 15008 16804 15048
rect 17037 15045 17049 15048
rect 17083 15045 17095 15079
rect 17037 15039 17095 15045
rect 18325 15079 18383 15085
rect 18325 15045 18337 15079
rect 18371 15076 18383 15079
rect 18506 15076 18512 15088
rect 18371 15048 18512 15076
rect 18371 15045 18383 15048
rect 18325 15039 18383 15045
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 19518 15076 19524 15088
rect 19479 15048 19524 15076
rect 19518 15036 19524 15048
rect 19576 15036 19582 15088
rect 19628 15076 19656 15116
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20404 15116 21496 15144
rect 20404 15104 20410 15116
rect 21269 15079 21327 15085
rect 21269 15076 21281 15079
rect 19628 15048 21281 15076
rect 21269 15045 21281 15048
rect 21315 15076 21327 15079
rect 21468 15076 21496 15116
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 25222 15144 25228 15156
rect 22152 15116 22197 15144
rect 22848 15116 25228 15144
rect 22152 15104 22158 15116
rect 22741 15079 22799 15085
rect 22741 15076 22753 15079
rect 21315 15048 21404 15076
rect 21468 15048 22753 15076
rect 21315 15045 21327 15048
rect 21269 15039 21327 15045
rect 16724 14980 16804 15008
rect 21376 15008 21404 15048
rect 22741 15045 22753 15048
rect 22787 15045 22799 15079
rect 22741 15039 22799 15045
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21376 14980 22201 15008
rect 16724 14968 16730 14980
rect 22189 14977 22201 14980
rect 22235 15008 22247 15011
rect 22848 15008 22876 15116
rect 25222 15104 25228 15116
rect 25280 15104 25286 15156
rect 28442 15144 28448 15156
rect 26436 15116 28448 15144
rect 24394 15076 24400 15088
rect 24355 15048 24400 15076
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 24489 15079 24547 15085
rect 24489 15045 24501 15079
rect 24535 15076 24547 15079
rect 25130 15076 25136 15088
rect 24535 15048 25136 15076
rect 24535 15045 24547 15048
rect 24489 15039 24547 15045
rect 25130 15036 25136 15048
rect 25188 15036 25194 15088
rect 26436 15085 26464 15116
rect 28442 15104 28448 15116
rect 28500 15104 28506 15156
rect 29454 15144 29460 15156
rect 28828 15116 29460 15144
rect 26421 15079 26479 15085
rect 26421 15045 26433 15079
rect 26467 15045 26479 15079
rect 26421 15039 26479 15045
rect 27062 15036 27068 15088
rect 27120 15076 27126 15088
rect 27249 15079 27307 15085
rect 27249 15076 27261 15079
rect 27120 15048 27261 15076
rect 27120 15036 27126 15048
rect 27249 15045 27261 15048
rect 27295 15045 27307 15079
rect 27249 15039 27307 15045
rect 27341 15079 27399 15085
rect 27341 15045 27353 15079
rect 27387 15076 27399 15079
rect 28534 15076 28540 15088
rect 27387 15048 28540 15076
rect 27387 15045 27399 15048
rect 27341 15039 27399 15045
rect 28534 15036 28540 15048
rect 28592 15036 28598 15088
rect 22235 14980 22876 15008
rect 22925 15011 22983 15017
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22925 14977 22937 15011
rect 22971 15008 22983 15011
rect 25038 15008 25044 15020
rect 22971 14980 23888 15008
rect 24999 14980 25044 15008
rect 22971 14977 22983 14980
rect 22925 14971 22983 14977
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 16540 14912 16957 14940
rect 16540 14900 16546 14912
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 17310 14940 17316 14952
rect 17271 14912 17316 14940
rect 16945 14903 17003 14909
rect 16960 14872 16988 14903
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 18233 14943 18291 14949
rect 18233 14928 18245 14943
rect 18156 14909 18245 14928
rect 18279 14909 18291 14943
rect 18156 14903 18291 14909
rect 18156 14900 18276 14903
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 19242 14940 19248 14952
rect 18380 14912 19248 14940
rect 18380 14900 18386 14912
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19426 14940 19432 14952
rect 19387 14912 19432 14940
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 23658 14940 23664 14952
rect 19812 14912 23664 14940
rect 18156 14872 18184 14900
rect 15856 14844 16804 14872
rect 16960 14844 18184 14872
rect 18785 14875 18843 14881
rect 14093 14807 14151 14813
rect 14093 14804 14105 14807
rect 13964 14776 14105 14804
rect 13964 14764 13970 14776
rect 14093 14773 14105 14776
rect 14139 14773 14151 14807
rect 14093 14767 14151 14773
rect 16209 14807 16267 14813
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 16666 14804 16672 14816
rect 16255 14776 16672 14804
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 16776 14804 16804 14844
rect 18785 14841 18797 14875
rect 18831 14872 18843 14875
rect 19812 14872 19840 14912
rect 23658 14900 23664 14912
rect 23716 14900 23722 14952
rect 23860 14940 23888 14980
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 25225 15011 25283 15017
rect 25225 14977 25237 15011
rect 25271 14977 25283 15011
rect 28828 15008 28856 15116
rect 29454 15104 29460 15116
rect 29512 15104 29518 15156
rect 29914 15104 29920 15156
rect 29972 15144 29978 15156
rect 31205 15147 31263 15153
rect 31205 15144 31217 15147
rect 29972 15116 31217 15144
rect 29972 15104 29978 15116
rect 31205 15113 31217 15116
rect 31251 15113 31263 15147
rect 31205 15107 31263 15113
rect 28905 15011 28963 15017
rect 28905 15008 28917 15011
rect 28828 14980 28917 15008
rect 25225 14971 25283 14977
rect 28905 14977 28917 14980
rect 28951 14977 28963 15011
rect 28905 14971 28963 14977
rect 25130 14940 25136 14952
rect 23860 14912 25136 14940
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 19978 14872 19984 14884
rect 18831 14844 19840 14872
rect 19939 14844 19984 14872
rect 18831 14841 18843 14844
rect 18785 14835 18843 14841
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 23937 14875 23995 14881
rect 23937 14841 23949 14875
rect 23983 14872 23995 14875
rect 24026 14872 24032 14884
rect 23983 14844 24032 14872
rect 23983 14841 23995 14844
rect 23937 14835 23995 14841
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 19334 14804 19340 14816
rect 16776 14776 19340 14804
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 20622 14804 20628 14816
rect 20583 14776 20628 14804
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 21177 14807 21235 14813
rect 21177 14773 21189 14807
rect 21223 14804 21235 14807
rect 21266 14804 21272 14816
rect 21223 14776 21272 14804
rect 21223 14773 21235 14776
rect 21177 14767 21235 14773
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 25240 14804 25268 14971
rect 28994 14968 29000 15020
rect 29052 15008 29058 15020
rect 29362 15008 29368 15020
rect 29052 14980 29368 15008
rect 29052 14968 29058 14980
rect 29362 14968 29368 14980
rect 29420 15008 29426 15020
rect 29549 15011 29607 15017
rect 29549 15008 29561 15011
rect 29420 14980 29561 15008
rect 29420 14968 29426 14980
rect 29549 14977 29561 14980
rect 29595 14977 29607 15011
rect 29549 14971 29607 14977
rect 30098 14968 30104 15020
rect 30156 15008 30162 15020
rect 30193 15011 30251 15017
rect 30193 15008 30205 15011
rect 30156 14980 30205 15008
rect 30156 14968 30162 14980
rect 30193 14977 30205 14980
rect 30239 14977 30251 15011
rect 30193 14971 30251 14977
rect 25590 14900 25596 14952
rect 25648 14940 25654 14952
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25648 14912 25881 14940
rect 25648 14900 25654 14912
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 26510 14940 26516 14952
rect 26423 14912 26516 14940
rect 25869 14903 25927 14909
rect 25884 14872 25912 14903
rect 26510 14900 26516 14912
rect 26568 14940 26574 14952
rect 27338 14940 27344 14952
rect 26568 14912 27344 14940
rect 26568 14900 26574 14912
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 28074 14940 28080 14952
rect 28035 14912 28080 14940
rect 28074 14900 28080 14912
rect 28132 14900 28138 14952
rect 28350 14900 28356 14952
rect 28408 14940 28414 14952
rect 30374 14940 30380 14952
rect 28408 14912 30380 14940
rect 28408 14900 28414 14912
rect 30374 14900 30380 14912
rect 30432 14900 30438 14952
rect 26326 14872 26332 14884
rect 25884 14844 26332 14872
rect 26326 14832 26332 14844
rect 26384 14872 26390 14884
rect 27062 14872 27068 14884
rect 26384 14844 27068 14872
rect 26384 14832 26390 14844
rect 27062 14832 27068 14844
rect 27120 14832 27126 14884
rect 27798 14872 27804 14884
rect 27632 14844 27804 14872
rect 27632 14804 27660 14844
rect 27798 14832 27804 14844
rect 27856 14832 27862 14884
rect 27890 14832 27896 14884
rect 27948 14872 27954 14884
rect 29457 14875 29515 14881
rect 29457 14872 29469 14875
rect 27948 14844 29469 14872
rect 27948 14832 27954 14844
rect 29457 14841 29469 14844
rect 29503 14841 29515 14875
rect 29457 14835 29515 14841
rect 29546 14832 29552 14884
rect 29604 14872 29610 14884
rect 30101 14875 30159 14881
rect 30101 14872 30113 14875
rect 29604 14844 30113 14872
rect 29604 14832 29610 14844
rect 30101 14841 30113 14844
rect 30147 14841 30159 14875
rect 30101 14835 30159 14841
rect 25240 14776 27660 14804
rect 27706 14764 27712 14816
rect 27764 14804 27770 14816
rect 28813 14807 28871 14813
rect 28813 14804 28825 14807
rect 27764 14776 28825 14804
rect 27764 14764 27770 14776
rect 28813 14773 28825 14776
rect 28859 14773 28871 14807
rect 28813 14767 28871 14773
rect 30282 14764 30288 14816
rect 30340 14804 30346 14816
rect 30653 14807 30711 14813
rect 30653 14804 30665 14807
rect 30340 14776 30665 14804
rect 30340 14764 30346 14776
rect 30653 14773 30665 14776
rect 30699 14773 30711 14807
rect 31220 14804 31248 15107
rect 31294 15104 31300 15156
rect 31352 15144 31358 15156
rect 33962 15144 33968 15156
rect 31352 15116 33968 15144
rect 31352 15104 31358 15116
rect 33962 15104 33968 15116
rect 34020 15104 34026 15156
rect 38102 14804 38108 14816
rect 31220 14776 38108 14804
rect 30653 14767 30711 14773
rect 38102 14764 38108 14776
rect 38160 14764 38166 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13725 14603 13783 14609
rect 13725 14600 13737 14603
rect 13219 14572 13737 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13725 14569 13737 14572
rect 13771 14600 13783 14603
rect 14182 14600 14188 14612
rect 13771 14572 14188 14600
rect 13771 14569 13783 14572
rect 13725 14563 13783 14569
rect 14182 14560 14188 14572
rect 14240 14600 14246 14612
rect 18690 14600 18696 14612
rect 14240 14572 18696 14600
rect 14240 14560 14246 14572
rect 9217 14535 9275 14541
rect 9217 14501 9229 14535
rect 9263 14532 9275 14535
rect 15378 14532 15384 14544
rect 9263 14504 15384 14532
rect 9263 14501 9275 14504
rect 9217 14495 9275 14501
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 8297 14399 8355 14405
rect 1903 14368 6914 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 6886 14260 6914 14368
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 9232 14396 9260 14495
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 8343 14368 9260 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 14884 14368 15485 14396
rect 14884 14356 14890 14368
rect 15473 14365 15485 14368
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 16592 14405 16620 14572
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 19518 14600 19524 14612
rect 19479 14572 19524 14600
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 23842 14600 23848 14612
rect 20036 14572 23848 14600
rect 20036 14560 20042 14572
rect 23842 14560 23848 14572
rect 23900 14560 23906 14612
rect 24394 14560 24400 14612
rect 24452 14600 24458 14612
rect 27065 14603 27123 14609
rect 27065 14600 27077 14603
rect 24452 14572 27077 14600
rect 24452 14560 24458 14572
rect 27065 14569 27077 14572
rect 27111 14569 27123 14603
rect 27065 14563 27123 14569
rect 27338 14560 27344 14612
rect 27396 14600 27402 14612
rect 29825 14603 29883 14609
rect 29825 14600 29837 14603
rect 27396 14572 29837 14600
rect 27396 14560 27402 14572
rect 29825 14569 29837 14572
rect 29871 14569 29883 14603
rect 29825 14563 29883 14569
rect 16669 14535 16727 14541
rect 16669 14501 16681 14535
rect 16715 14532 16727 14535
rect 20070 14532 20076 14544
rect 16715 14504 20076 14532
rect 16715 14501 16727 14504
rect 16669 14495 16727 14501
rect 20070 14492 20076 14504
rect 20128 14492 20134 14544
rect 20346 14532 20352 14544
rect 20180 14504 20352 14532
rect 18049 14467 18107 14473
rect 18049 14464 18061 14467
rect 17052 14436 18061 14464
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15896 14368 15945 14396
rect 15896 14356 15902 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 17052 14328 17080 14436
rect 18049 14433 18061 14436
rect 18095 14433 18107 14467
rect 18049 14427 18107 14433
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 19426 14464 19432 14476
rect 18196 14436 19432 14464
rect 18196 14424 18202 14436
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 20180 14464 20208 14504
rect 20346 14492 20352 14504
rect 20404 14492 20410 14544
rect 25038 14532 25044 14544
rect 22664 14504 25044 14532
rect 19720 14436 20208 14464
rect 17218 14396 17224 14408
rect 17179 14368 17224 14396
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17460 14368 17877 14396
rect 17460 14356 17466 14368
rect 17865 14365 17877 14368
rect 17911 14396 17923 14399
rect 19610 14396 19616 14408
rect 17911 14368 19334 14396
rect 19571 14368 19616 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 16040 14300 17080 14328
rect 17313 14331 17371 14337
rect 8113 14263 8171 14269
rect 8113 14260 8125 14263
rect 6886 14232 8125 14260
rect 8113 14229 8125 14232
rect 8159 14229 8171 14263
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 8113 14223 8171 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 15378 14260 15384 14272
rect 15339 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 16040 14269 16068 14300
rect 17313 14297 17325 14331
rect 17359 14328 17371 14331
rect 18322 14328 18328 14340
rect 17359 14300 18328 14328
rect 17359 14297 17371 14300
rect 17313 14291 17371 14297
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 18509 14331 18567 14337
rect 18509 14297 18521 14331
rect 18555 14328 18567 14331
rect 19150 14328 19156 14340
rect 18555 14300 19156 14328
rect 18555 14297 18567 14300
rect 18509 14291 18567 14297
rect 19150 14288 19156 14300
rect 19208 14288 19214 14340
rect 19306 14328 19334 14368
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 19720 14328 19748 14436
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 21453 14467 21511 14473
rect 21453 14464 21465 14467
rect 20312 14436 21465 14464
rect 20312 14424 20318 14436
rect 21453 14433 21465 14436
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 20254 14328 20260 14340
rect 19306 14300 19748 14328
rect 20215 14300 20260 14328
rect 20254 14288 20260 14300
rect 20312 14288 20318 14340
rect 20349 14331 20407 14337
rect 20349 14297 20361 14331
rect 20395 14297 20407 14331
rect 20898 14328 20904 14340
rect 20859 14300 20904 14328
rect 20349 14291 20407 14297
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14229 16083 14263
rect 16025 14223 16083 14229
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 20364 14260 20392 14291
rect 20898 14288 20904 14300
rect 20956 14288 20962 14340
rect 18012 14232 20392 14260
rect 18012 14220 18018 14232
rect 20438 14220 20444 14272
rect 20496 14260 20502 14272
rect 21266 14260 21272 14272
rect 20496 14232 21272 14260
rect 20496 14220 20502 14232
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 21468 14260 21496 14427
rect 21542 14356 21548 14408
rect 21600 14396 21606 14408
rect 21600 14368 21645 14396
rect 21600 14356 21606 14368
rect 21818 14356 21824 14408
rect 21876 14396 21882 14408
rect 22005 14399 22063 14405
rect 22005 14396 22017 14399
rect 21876 14368 22017 14396
rect 21876 14356 21882 14368
rect 22005 14365 22017 14368
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 21560 14328 21588 14356
rect 22664 14328 22692 14504
rect 25038 14492 25044 14504
rect 25096 14532 25102 14544
rect 25314 14532 25320 14544
rect 25096 14504 25320 14532
rect 25096 14492 25102 14504
rect 25314 14492 25320 14504
rect 25372 14492 25378 14544
rect 26050 14492 26056 14544
rect 26108 14532 26114 14544
rect 28997 14535 29055 14541
rect 28997 14532 29009 14535
rect 26108 14504 27660 14532
rect 26108 14492 26114 14504
rect 23014 14464 23020 14476
rect 22975 14436 23020 14464
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 25774 14464 25780 14476
rect 24044 14436 25780 14464
rect 24044 14405 24072 14436
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 26142 14464 26148 14476
rect 26103 14436 26148 14464
rect 26142 14424 26148 14436
rect 26200 14424 26206 14476
rect 26234 14424 26240 14476
rect 26292 14464 26298 14476
rect 27154 14464 27160 14476
rect 26292 14436 27160 14464
rect 26292 14424 26298 14436
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 27632 14473 27660 14504
rect 27724 14504 29009 14532
rect 27617 14467 27675 14473
rect 27617 14433 27629 14467
rect 27663 14433 27675 14467
rect 27617 14427 27675 14433
rect 24029 14399 24087 14405
rect 24029 14365 24041 14399
rect 24075 14365 24087 14399
rect 24029 14359 24087 14365
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14396 24823 14399
rect 25682 14396 25688 14408
rect 24811 14368 25688 14396
rect 24811 14365 24823 14368
rect 24765 14359 24823 14365
rect 25682 14356 25688 14368
rect 25740 14356 25746 14408
rect 26694 14356 26700 14408
rect 26752 14396 26758 14408
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26752 14368 26985 14396
rect 26752 14356 26758 14368
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 21560 14300 22692 14328
rect 23201 14331 23259 14337
rect 23201 14297 23213 14331
rect 23247 14297 23259 14331
rect 23201 14291 23259 14297
rect 22002 14260 22008 14272
rect 21468 14232 22008 14260
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 22097 14263 22155 14269
rect 22097 14229 22109 14263
rect 22143 14260 22155 14263
rect 23216 14260 23244 14291
rect 23290 14288 23296 14340
rect 23348 14328 23354 14340
rect 23348 14300 23393 14328
rect 23348 14288 23354 14300
rect 23842 14288 23848 14340
rect 23900 14328 23906 14340
rect 26142 14328 26148 14340
rect 23900 14300 26148 14328
rect 23900 14288 23906 14300
rect 26142 14288 26148 14300
rect 26200 14288 26206 14340
rect 26234 14288 26240 14340
rect 26292 14328 26298 14340
rect 26329 14331 26387 14337
rect 26329 14328 26341 14331
rect 26292 14300 26341 14328
rect 26292 14288 26298 14300
rect 26329 14297 26341 14300
rect 26375 14297 26387 14331
rect 26329 14291 26387 14297
rect 26421 14331 26479 14337
rect 26421 14297 26433 14331
rect 26467 14328 26479 14331
rect 27338 14328 27344 14340
rect 26467 14300 27344 14328
rect 26467 14297 26479 14300
rect 26421 14291 26479 14297
rect 27338 14288 27344 14300
rect 27396 14328 27402 14340
rect 27724 14328 27752 14504
rect 28997 14501 29009 14504
rect 29043 14501 29055 14535
rect 28997 14495 29055 14501
rect 29086 14492 29092 14544
rect 29144 14532 29150 14544
rect 30006 14532 30012 14544
rect 29144 14504 30012 14532
rect 29144 14492 29150 14504
rect 30006 14492 30012 14504
rect 30064 14532 30070 14544
rect 30064 14504 30604 14532
rect 30064 14492 30070 14504
rect 28074 14424 28080 14476
rect 28132 14464 28138 14476
rect 30469 14467 30527 14473
rect 30469 14464 30481 14467
rect 28132 14436 30481 14464
rect 28132 14424 28138 14436
rect 30469 14433 30481 14436
rect 30515 14433 30527 14467
rect 30469 14427 30527 14433
rect 27798 14356 27804 14408
rect 27856 14356 27862 14408
rect 28442 14396 28448 14408
rect 28403 14368 28448 14396
rect 28442 14356 28448 14368
rect 28500 14356 28506 14408
rect 29089 14399 29147 14405
rect 29089 14365 29101 14399
rect 29135 14365 29147 14399
rect 29914 14396 29920 14408
rect 29875 14368 29920 14396
rect 29089 14359 29147 14365
rect 27396 14300 27752 14328
rect 27816 14328 27844 14356
rect 29104 14328 29132 14359
rect 29914 14356 29920 14368
rect 29972 14356 29978 14408
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30576 14396 30604 14504
rect 30423 14368 30604 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 30282 14328 30288 14340
rect 27816 14300 30288 14328
rect 27396 14288 27402 14300
rect 30282 14288 30288 14300
rect 30340 14328 30346 14340
rect 31573 14331 31631 14337
rect 31573 14328 31585 14331
rect 30340 14300 31585 14328
rect 30340 14288 30346 14300
rect 31573 14297 31585 14300
rect 31619 14328 31631 14331
rect 31619 14300 31754 14328
rect 31619 14297 31631 14300
rect 31573 14291 31631 14297
rect 22143 14232 23244 14260
rect 22143 14229 22155 14232
rect 22097 14223 22155 14229
rect 23382 14220 23388 14272
rect 23440 14260 23446 14272
rect 23937 14263 23995 14269
rect 23937 14260 23949 14263
rect 23440 14232 23949 14260
rect 23440 14220 23446 14232
rect 23937 14229 23949 14232
rect 23983 14229 23995 14263
rect 24670 14260 24676 14272
rect 24631 14232 24676 14260
rect 23937 14223 23995 14229
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 25222 14260 25228 14272
rect 25183 14232 25228 14260
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 25314 14220 25320 14272
rect 25372 14260 25378 14272
rect 26050 14260 26056 14272
rect 25372 14232 26056 14260
rect 25372 14220 25378 14232
rect 26050 14220 26056 14232
rect 26108 14220 26114 14272
rect 27798 14220 27804 14272
rect 27856 14260 27862 14272
rect 28353 14263 28411 14269
rect 28353 14260 28365 14263
rect 27856 14232 28365 14260
rect 27856 14220 27862 14232
rect 28353 14229 28365 14232
rect 28399 14229 28411 14263
rect 28353 14223 28411 14229
rect 29730 14220 29736 14272
rect 29788 14260 29794 14272
rect 30374 14260 30380 14272
rect 29788 14232 30380 14260
rect 29788 14220 29794 14232
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 31113 14263 31171 14269
rect 31113 14229 31125 14263
rect 31159 14260 31171 14263
rect 31202 14260 31208 14272
rect 31159 14232 31208 14260
rect 31159 14229 31171 14232
rect 31113 14223 31171 14229
rect 31202 14220 31208 14232
rect 31260 14220 31266 14272
rect 31726 14260 31754 14300
rect 36814 14260 36820 14272
rect 31726 14232 36820 14260
rect 36814 14220 36820 14232
rect 36872 14220 36878 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14056 16267 14059
rect 17402 14056 17408 14068
rect 16255 14028 17408 14056
rect 16255 14025 16267 14028
rect 16209 14019 16267 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 19981 14059 20039 14065
rect 17543 14028 19196 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 19168 14000 19196 14028
rect 19981 14025 19993 14059
rect 20027 14056 20039 14059
rect 22094 14056 22100 14068
rect 20027 14028 22100 14056
rect 20027 14025 20039 14028
rect 19981 14019 20039 14025
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 22186 14016 22192 14068
rect 22244 14056 22250 14068
rect 22244 14028 27200 14056
rect 22244 14016 22250 14028
rect 13354 13948 13360 14000
rect 13412 13988 13418 14000
rect 13630 13988 13636 14000
rect 13412 13960 13636 13988
rect 13412 13948 13418 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 14274 13988 14280 14000
rect 14235 13960 14280 13988
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 18138 13988 18144 14000
rect 18099 13960 18144 13988
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 19058 13988 19064 14000
rect 19019 13960 19064 13988
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 19150 13948 19156 14000
rect 19208 13988 19214 14000
rect 19208 13960 19253 13988
rect 19208 13948 19214 13960
rect 20346 13948 20352 14000
rect 20404 13988 20410 14000
rect 20625 13991 20683 13997
rect 20625 13988 20637 13991
rect 20404 13960 20637 13988
rect 20404 13948 20410 13960
rect 20625 13957 20637 13960
rect 20671 13957 20683 13991
rect 20625 13951 20683 13957
rect 20717 13991 20775 13997
rect 20717 13957 20729 13991
rect 20763 13988 20775 13991
rect 23382 13988 23388 14000
rect 20763 13960 23388 13988
rect 20763 13957 20775 13960
rect 20717 13951 20775 13957
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 23937 13991 23995 13997
rect 23937 13957 23949 13991
rect 23983 13988 23995 13991
rect 24670 13988 24676 14000
rect 23983 13960 24676 13988
rect 23983 13957 23995 13960
rect 23937 13951 23995 13957
rect 24670 13948 24676 13960
rect 24728 13948 24734 14000
rect 24762 13948 24768 14000
rect 24820 13988 24826 14000
rect 25777 13991 25835 13997
rect 25777 13988 25789 13991
rect 24820 13960 25789 13988
rect 24820 13948 24826 13960
rect 25777 13957 25789 13960
rect 25823 13957 25835 13991
rect 26326 13988 26332 14000
rect 26287 13960 26332 13988
rect 25777 13951 25835 13957
rect 14182 13920 14188 13932
rect 14143 13892 14188 13920
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15470 13920 15476 13932
rect 14292 13892 15476 13920
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 12621 13855 12679 13861
rect 12621 13852 12633 13855
rect 4120 13824 12633 13852
rect 4120 13812 4126 13824
rect 12621 13821 12633 13824
rect 12667 13852 12679 13855
rect 14292 13852 14320 13892
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 16117 13926 16175 13929
rect 16117 13923 16252 13926
rect 16117 13889 16129 13923
rect 16163 13898 16252 13923
rect 16163 13889 16175 13898
rect 16117 13883 16175 13889
rect 15010 13852 15016 13864
rect 12667 13824 14320 13852
rect 14971 13824 15016 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 16224 13852 16252 13898
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16850 13920 16856 13932
rect 16632 13892 16856 13920
rect 16632 13880 16638 13892
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17034 13920 17040 13932
rect 16995 13892 17040 13920
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 19889 13923 19947 13929
rect 19889 13920 19901 13923
rect 19392 13892 19901 13920
rect 19392 13880 19398 13892
rect 19889 13889 19901 13892
rect 19935 13920 19947 13923
rect 20438 13920 20444 13932
rect 19935 13892 20444 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 21358 13880 21364 13932
rect 21416 13920 21422 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21416 13892 22201 13920
rect 21416 13880 21422 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 24578 13920 24584 13932
rect 24539 13892 24584 13920
rect 22189 13883 22247 13889
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 25038 13880 25044 13932
rect 25096 13920 25102 13932
rect 25225 13923 25283 13929
rect 25225 13920 25237 13923
rect 25096 13892 25237 13920
rect 25096 13880 25102 13892
rect 25225 13889 25237 13892
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 16298 13852 16304 13864
rect 16224 13824 16304 13852
rect 16298 13812 16304 13824
rect 16356 13852 16362 13864
rect 16758 13852 16764 13864
rect 16356 13824 16764 13852
rect 16356 13812 16362 13824
rect 16758 13812 16764 13824
rect 16816 13852 16822 13864
rect 18138 13852 18144 13864
rect 16816 13824 18144 13852
rect 16816 13812 16822 13824
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 18380 13824 22017 13852
rect 18380 13812 18386 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 23753 13855 23811 13861
rect 23753 13821 23765 13855
rect 23799 13852 23811 13855
rect 23842 13852 23848 13864
rect 23799 13824 23848 13852
rect 23799 13821 23811 13824
rect 23753 13815 23811 13821
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13852 24087 13855
rect 25314 13852 25320 13864
rect 24075 13824 25320 13852
rect 24075 13821 24087 13824
rect 24029 13815 24087 13821
rect 25314 13812 25320 13824
rect 25372 13812 25378 13864
rect 25792 13852 25820 13951
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 26418 13948 26424 14000
rect 26476 13988 26482 14000
rect 27062 13988 27068 14000
rect 26476 13960 27068 13988
rect 26476 13948 26482 13960
rect 27062 13948 27068 13960
rect 27120 13948 27126 14000
rect 27172 13997 27200 14028
rect 27246 14016 27252 14068
rect 27304 14056 27310 14068
rect 27304 14028 29868 14056
rect 27304 14016 27310 14028
rect 27157 13991 27215 13997
rect 27157 13957 27169 13991
rect 27203 13957 27215 13991
rect 27706 13988 27712 14000
rect 27667 13960 27712 13988
rect 27157 13951 27215 13957
rect 27706 13948 27712 13960
rect 27764 13948 27770 14000
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 28537 13991 28595 13997
rect 27856 13960 27901 13988
rect 27856 13948 27862 13960
rect 28537 13957 28549 13991
rect 28583 13988 28595 13991
rect 28583 13960 29500 13988
rect 28583 13957 28595 13960
rect 28537 13951 28595 13957
rect 26421 13855 26479 13861
rect 25792 13824 26390 13852
rect 13170 13784 13176 13796
rect 13131 13756 13176 13784
rect 13170 13744 13176 13756
rect 13228 13744 13234 13796
rect 14734 13744 14740 13796
rect 14792 13784 14798 13796
rect 18046 13784 18052 13796
rect 14792 13756 18052 13784
rect 14792 13744 14798 13756
rect 18046 13744 18052 13756
rect 18104 13744 18110 13796
rect 21082 13784 21088 13796
rect 20456 13756 21088 13784
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 20456 13716 20484 13756
rect 21082 13744 21088 13756
rect 21140 13744 21146 13796
rect 21174 13744 21180 13796
rect 21232 13784 21238 13796
rect 23382 13784 23388 13796
rect 21232 13756 23388 13784
rect 21232 13744 21238 13756
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 23658 13744 23664 13796
rect 23716 13784 23722 13796
rect 23934 13784 23940 13796
rect 23716 13756 23940 13784
rect 23716 13744 23722 13756
rect 23934 13744 23940 13756
rect 23992 13744 23998 13796
rect 24578 13744 24584 13796
rect 24636 13784 24642 13796
rect 26362 13784 26390 13824
rect 26421 13821 26433 13855
rect 26467 13852 26479 13855
rect 27798 13852 27804 13864
rect 26467 13824 27804 13852
rect 26467 13821 26479 13824
rect 26421 13815 26479 13821
rect 27798 13812 27804 13824
rect 27856 13812 27862 13864
rect 28074 13812 28080 13864
rect 28132 13852 28138 13864
rect 28445 13855 28503 13861
rect 28445 13852 28457 13855
rect 28132 13824 28457 13852
rect 28132 13812 28138 13824
rect 28445 13821 28457 13824
rect 28491 13821 28503 13855
rect 28902 13852 28908 13864
rect 28863 13824 28908 13852
rect 28445 13815 28503 13821
rect 28902 13812 28908 13824
rect 28960 13812 28966 13864
rect 27154 13784 27160 13796
rect 24636 13756 25820 13784
rect 26362 13756 27160 13784
rect 24636 13744 24642 13756
rect 14240 13688 20484 13716
rect 14240 13676 14246 13688
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 22373 13719 22431 13725
rect 22373 13716 22385 13719
rect 20588 13688 22385 13716
rect 20588 13676 20594 13688
rect 22373 13685 22385 13688
rect 22419 13685 22431 13719
rect 22373 13679 22431 13685
rect 24673 13719 24731 13725
rect 24673 13685 24685 13719
rect 24719 13716 24731 13719
rect 24762 13716 24768 13728
rect 24719 13688 24768 13716
rect 24719 13685 24731 13688
rect 24673 13679 24731 13685
rect 24762 13676 24768 13688
rect 24820 13676 24826 13728
rect 25792 13716 25820 13756
rect 27154 13744 27160 13756
rect 27212 13744 27218 13796
rect 28258 13744 28264 13796
rect 28316 13784 28322 13796
rect 29178 13784 29184 13796
rect 28316 13756 29184 13784
rect 28316 13744 28322 13756
rect 29178 13744 29184 13756
rect 29236 13744 29242 13796
rect 29472 13784 29500 13960
rect 29730 13920 29736 13932
rect 29691 13892 29736 13920
rect 29730 13880 29736 13892
rect 29788 13880 29794 13932
rect 29840 13920 29868 14028
rect 30190 14016 30196 14068
rect 30248 14056 30254 14068
rect 30285 14059 30343 14065
rect 30285 14056 30297 14059
rect 30248 14028 30297 14056
rect 30248 14016 30254 14028
rect 30285 14025 30297 14028
rect 30331 14025 30343 14059
rect 30285 14019 30343 14025
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 31481 14059 31539 14065
rect 31481 14056 31493 14059
rect 30524 14028 31493 14056
rect 30524 14016 30530 14028
rect 31481 14025 31493 14028
rect 31527 14025 31539 14059
rect 31481 14019 31539 14025
rect 29914 13948 29920 14000
rect 29972 13988 29978 14000
rect 29972 13960 30880 13988
rect 29972 13948 29978 13960
rect 30852 13929 30880 13960
rect 30193 13923 30251 13929
rect 30193 13920 30205 13923
rect 29840 13892 30205 13920
rect 30193 13889 30205 13892
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 30837 13923 30895 13929
rect 30837 13889 30849 13923
rect 30883 13889 30895 13923
rect 30837 13883 30895 13889
rect 29638 13852 29644 13864
rect 29599 13824 29644 13852
rect 29638 13812 29644 13824
rect 29696 13812 29702 13864
rect 29822 13812 29828 13864
rect 29880 13852 29886 13864
rect 30929 13855 30987 13861
rect 30929 13852 30941 13855
rect 29880 13824 30941 13852
rect 29880 13812 29886 13824
rect 30929 13821 30941 13824
rect 30975 13821 30987 13855
rect 31570 13852 31576 13864
rect 30929 13815 30987 13821
rect 31036 13824 31576 13852
rect 31036 13784 31064 13824
rect 31570 13812 31576 13824
rect 31628 13812 31634 13864
rect 33134 13812 33140 13864
rect 33192 13852 33198 13864
rect 38013 13855 38071 13861
rect 38013 13852 38025 13855
rect 33192 13824 38025 13852
rect 33192 13812 33198 13824
rect 38013 13821 38025 13824
rect 38059 13821 38071 13855
rect 38286 13852 38292 13864
rect 38247 13824 38292 13852
rect 38013 13815 38071 13821
rect 38286 13812 38292 13824
rect 38344 13812 38350 13864
rect 29472 13756 31064 13784
rect 29730 13716 29736 13728
rect 25792 13688 29736 13716
rect 29730 13676 29736 13688
rect 29788 13676 29794 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 10594 13512 10600 13524
rect 10555 13484 10600 13512
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 10704 13484 14872 13512
rect 10704 13317 10732 13484
rect 13633 13447 13691 13453
rect 13633 13413 13645 13447
rect 13679 13444 13691 13447
rect 14734 13444 14740 13456
rect 13679 13416 14740 13444
rect 13679 13413 13691 13416
rect 13633 13407 13691 13413
rect 14734 13404 14740 13416
rect 14792 13404 14798 13456
rect 14844 13444 14872 13484
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16850 13512 16856 13524
rect 15528 13484 16856 13512
rect 15528 13472 15534 13484
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 16945 13515 17003 13521
rect 16945 13481 16957 13515
rect 16991 13512 17003 13515
rect 17954 13512 17960 13524
rect 16991 13484 17960 13512
rect 16991 13481 17003 13484
rect 16945 13475 17003 13481
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 19242 13472 19248 13524
rect 19300 13512 19306 13524
rect 19300 13484 20300 13512
rect 19300 13472 19306 13484
rect 17218 13444 17224 13456
rect 14844 13416 17224 13444
rect 17218 13404 17224 13416
rect 17276 13404 17282 13456
rect 20162 13444 20168 13456
rect 18708 13416 20168 13444
rect 14366 13376 14372 13388
rect 14327 13348 14372 13376
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 16114 13376 16120 13388
rect 15703 13348 16120 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 16114 13336 16120 13348
rect 16172 13376 16178 13388
rect 16172 13348 17264 13376
rect 16172 13336 16178 13348
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15286 13308 15292 13320
rect 15059 13280 15292 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13308 16911 13311
rect 17126 13308 17132 13320
rect 16899 13280 17132 13308
rect 16899 13277 16911 13280
rect 16853 13271 16911 13277
rect 12069 13243 12127 13249
rect 12069 13209 12081 13243
rect 12115 13240 12127 13243
rect 13173 13243 13231 13249
rect 13173 13240 13185 13243
rect 12115 13212 13185 13240
rect 12115 13209 12127 13212
rect 12069 13203 12127 13209
rect 13173 13209 13185 13212
rect 13219 13240 13231 13243
rect 14366 13240 14372 13252
rect 13219 13212 14372 13240
rect 13219 13209 13231 13212
rect 13173 13203 13231 13209
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13209 14519 13243
rect 14461 13203 14519 13209
rect 12621 13175 12679 13181
rect 12621 13141 12633 13175
rect 12667 13172 12679 13175
rect 13354 13172 13360 13184
rect 12667 13144 13360 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 14476 13172 14504 13203
rect 15746 13200 15752 13252
rect 15804 13240 15810 13252
rect 16316 13240 16344 13271
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17236 13240 17264 13348
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18708 13376 18736 13416
rect 20162 13404 20168 13416
rect 20220 13404 20226 13456
rect 20272 13444 20300 13484
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 20404 13484 21864 13512
rect 20404 13472 20410 13484
rect 20438 13444 20444 13456
rect 20272 13416 20444 13444
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 20898 13404 20904 13456
rect 20956 13444 20962 13456
rect 21634 13444 21640 13456
rect 20956 13416 21640 13444
rect 20956 13404 20962 13416
rect 21634 13404 21640 13416
rect 21692 13444 21698 13456
rect 21729 13447 21787 13453
rect 21729 13444 21741 13447
rect 21692 13416 21741 13444
rect 21692 13404 21698 13416
rect 21729 13413 21741 13416
rect 21775 13413 21787 13447
rect 21836 13444 21864 13484
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22554 13512 22560 13524
rect 22060 13484 22560 13512
rect 22060 13472 22066 13484
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 28442 13512 28448 13524
rect 23308 13484 28448 13512
rect 23308 13444 23336 13484
rect 28442 13472 28448 13484
rect 28500 13472 28506 13524
rect 28626 13472 28632 13524
rect 28684 13512 28690 13524
rect 31110 13512 31116 13524
rect 28684 13484 29960 13512
rect 31071 13484 31116 13512
rect 28684 13472 28690 13484
rect 21836 13416 23336 13444
rect 21729 13407 21787 13413
rect 23382 13404 23388 13456
rect 23440 13444 23446 13456
rect 23440 13416 27384 13444
rect 23440 13404 23446 13416
rect 18104 13348 18736 13376
rect 18104 13336 18110 13348
rect 18708 13317 18736 13348
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19484 13348 19901 13376
rect 19484 13336 19490 13348
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 20588 13348 21128 13376
rect 20588 13336 20594 13348
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 17589 13243 17647 13249
rect 17589 13240 17601 13243
rect 15804 13212 15849 13240
rect 16316 13212 17172 13240
rect 17236 13212 17601 13240
rect 15804 13200 15810 13212
rect 15378 13172 15384 13184
rect 14476 13144 15384 13172
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 17144 13172 17172 13212
rect 17589 13209 17601 13212
rect 17635 13209 17647 13243
rect 17589 13203 17647 13209
rect 17681 13243 17739 13249
rect 17681 13209 17693 13243
rect 17727 13240 17739 13243
rect 18046 13240 18052 13252
rect 17727 13212 18052 13240
rect 17727 13209 17739 13212
rect 17681 13203 17739 13209
rect 18046 13200 18052 13212
rect 18104 13200 18110 13252
rect 18233 13243 18291 13249
rect 18233 13209 18245 13243
rect 18279 13240 18291 13243
rect 18966 13240 18972 13252
rect 18279 13212 18972 13240
rect 18279 13209 18291 13212
rect 18233 13203 18291 13209
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 20809 13243 20867 13249
rect 20809 13240 20821 13243
rect 20772 13212 20821 13240
rect 20772 13200 20778 13212
rect 20809 13209 20821 13212
rect 20855 13209 20867 13243
rect 20809 13203 20867 13209
rect 20901 13243 20959 13249
rect 20901 13209 20913 13243
rect 20947 13240 20959 13243
rect 21100 13240 21128 13348
rect 21266 13336 21272 13388
rect 21324 13376 21330 13388
rect 21324 13348 22600 13376
rect 21324 13336 21330 13348
rect 20947 13212 21128 13240
rect 20947 13209 20959 13212
rect 20901 13203 20959 13209
rect 22094 13200 22100 13252
rect 22152 13240 22158 13252
rect 22189 13243 22247 13249
rect 22189 13240 22201 13243
rect 22152 13212 22201 13240
rect 22152 13200 22158 13212
rect 22189 13209 22201 13212
rect 22235 13209 22247 13243
rect 22189 13203 22247 13209
rect 22278 13200 22284 13252
rect 22336 13240 22342 13252
rect 22572 13240 22600 13348
rect 22738 13336 22744 13388
rect 22796 13376 22802 13388
rect 23106 13376 23112 13388
rect 22796 13348 23112 13376
rect 22796 13336 22802 13348
rect 23106 13336 23112 13348
rect 23164 13336 23170 13388
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13376 25375 13379
rect 25590 13376 25596 13388
rect 25363 13348 25596 13376
rect 25363 13345 25375 13348
rect 25317 13339 25375 13345
rect 25590 13336 25596 13348
rect 25648 13336 25654 13388
rect 25682 13336 25688 13388
rect 25740 13376 25746 13388
rect 25958 13376 25964 13388
rect 25740 13348 25964 13376
rect 25740 13336 25746 13348
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 27356 13385 27384 13416
rect 27522 13404 27528 13456
rect 27580 13444 27586 13456
rect 29086 13444 29092 13456
rect 27580 13416 29092 13444
rect 27580 13404 27586 13416
rect 29086 13404 29092 13416
rect 29144 13404 29150 13456
rect 26605 13379 26663 13385
rect 26605 13376 26617 13379
rect 26568 13348 26617 13376
rect 26568 13336 26574 13348
rect 26605 13345 26617 13348
rect 26651 13345 26663 13379
rect 26605 13339 26663 13345
rect 27341 13379 27399 13385
rect 27341 13345 27353 13379
rect 27387 13345 27399 13379
rect 27341 13339 27399 13345
rect 27430 13336 27436 13388
rect 27488 13376 27494 13388
rect 29825 13379 29883 13385
rect 29825 13376 29837 13379
rect 27488 13348 29837 13376
rect 27488 13336 27494 13348
rect 29825 13345 29837 13348
rect 29871 13345 29883 13379
rect 29825 13339 29883 13345
rect 29932 13376 29960 13484
rect 31110 13472 31116 13484
rect 31168 13472 31174 13524
rect 38286 13512 38292 13524
rect 38247 13484 38292 13512
rect 38286 13472 38292 13484
rect 38344 13472 38350 13524
rect 31202 13376 31208 13388
rect 29932 13348 31208 13376
rect 27985 13311 28043 13317
rect 27985 13277 27997 13311
rect 28031 13308 28043 13311
rect 28258 13308 28264 13320
rect 28031 13280 28264 13308
rect 28031 13277 28043 13280
rect 27985 13271 28043 13277
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 29178 13268 29184 13320
rect 29236 13308 29242 13320
rect 29932 13317 29960 13348
rect 31202 13336 31208 13348
rect 31260 13376 31266 13388
rect 31757 13379 31815 13385
rect 31757 13376 31769 13379
rect 31260 13348 31769 13376
rect 31260 13336 31266 13348
rect 31757 13345 31769 13348
rect 31803 13376 31815 13379
rect 37090 13376 37096 13388
rect 31803 13348 37096 13376
rect 31803 13345 31815 13348
rect 31757 13339 31815 13345
rect 37090 13336 37096 13348
rect 37148 13336 37154 13388
rect 29917 13311 29975 13317
rect 29236 13280 29281 13308
rect 29236 13268 29242 13280
rect 29917 13277 29929 13311
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 30561 13311 30619 13317
rect 30561 13277 30573 13311
rect 30607 13277 30619 13311
rect 30561 13271 30619 13277
rect 22830 13240 22836 13252
rect 22336 13212 22381 13240
rect 22572 13212 22692 13240
rect 22791 13212 22836 13240
rect 22336 13200 22342 13212
rect 18506 13172 18512 13184
rect 17144 13144 18512 13172
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 18785 13175 18843 13181
rect 18785 13141 18797 13175
rect 18831 13172 18843 13175
rect 22554 13172 22560 13184
rect 18831 13144 22560 13172
rect 18831 13141 18843 13144
rect 18785 13135 18843 13141
rect 22554 13132 22560 13144
rect 22612 13132 22618 13184
rect 22664 13172 22692 13212
rect 22830 13200 22836 13212
rect 22888 13200 22894 13252
rect 23385 13243 23443 13249
rect 23385 13209 23397 13243
rect 23431 13209 23443 13243
rect 23385 13203 23443 13209
rect 23477 13243 23535 13249
rect 23477 13209 23489 13243
rect 23523 13240 23535 13243
rect 24673 13243 24731 13249
rect 24673 13240 24685 13243
rect 23523 13212 24685 13240
rect 23523 13209 23535 13212
rect 23477 13203 23535 13209
rect 24673 13209 24685 13212
rect 24719 13209 24731 13243
rect 24673 13203 24731 13209
rect 23400 13172 23428 13203
rect 22664 13144 23428 13172
rect 24688 13172 24716 13203
rect 24762 13200 24768 13252
rect 24820 13240 24826 13252
rect 24820 13212 24865 13240
rect 24820 13200 24826 13212
rect 24946 13200 24952 13252
rect 25004 13240 25010 13252
rect 25958 13240 25964 13252
rect 25004 13212 25964 13240
rect 25004 13200 25010 13212
rect 25958 13200 25964 13212
rect 26016 13200 26022 13252
rect 26513 13243 26571 13249
rect 26513 13209 26525 13243
rect 26559 13209 26571 13243
rect 26513 13203 26571 13209
rect 27433 13243 27491 13249
rect 27433 13209 27445 13243
rect 27479 13240 27491 13243
rect 27614 13240 27620 13252
rect 27479 13212 27620 13240
rect 27479 13209 27491 13212
rect 27433 13203 27491 13209
rect 26418 13172 26424 13184
rect 24688 13144 26424 13172
rect 26418 13132 26424 13144
rect 26476 13132 26482 13184
rect 26528 13172 26556 13203
rect 27614 13200 27620 13212
rect 27672 13200 27678 13252
rect 27706 13200 27712 13252
rect 27764 13240 27770 13252
rect 28537 13243 28595 13249
rect 28537 13240 28549 13243
rect 27764 13212 28549 13240
rect 27764 13200 27770 13212
rect 28537 13209 28549 13212
rect 28583 13209 28595 13243
rect 28537 13203 28595 13209
rect 28629 13243 28687 13249
rect 28629 13209 28641 13243
rect 28675 13240 28687 13243
rect 28902 13240 28908 13252
rect 28675 13212 28908 13240
rect 28675 13209 28687 13212
rect 28629 13203 28687 13209
rect 28902 13200 28908 13212
rect 28960 13200 28966 13252
rect 30576 13240 30604 13271
rect 30742 13268 30748 13320
rect 30800 13308 30806 13320
rect 31021 13311 31079 13317
rect 31021 13308 31033 13311
rect 30800 13280 31033 13308
rect 30800 13268 30806 13280
rect 31021 13277 31033 13280
rect 31067 13277 31079 13311
rect 31021 13271 31079 13277
rect 30576 13212 32352 13240
rect 27890 13172 27896 13184
rect 26528 13144 27896 13172
rect 27890 13132 27896 13144
rect 27948 13132 27954 13184
rect 28166 13132 28172 13184
rect 28224 13172 28230 13184
rect 30190 13172 30196 13184
rect 28224 13144 30196 13172
rect 28224 13132 28230 13144
rect 30190 13132 30196 13144
rect 30248 13132 30254 13184
rect 30466 13172 30472 13184
rect 30427 13144 30472 13172
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 32324 13181 32352 13212
rect 32309 13175 32367 13181
rect 32309 13141 32321 13175
rect 32355 13172 32367 13175
rect 37918 13172 37924 13184
rect 32355 13144 37924 13172
rect 32355 13141 32367 13144
rect 32309 13135 32367 13141
rect 37918 13132 37924 13144
rect 37976 13132 37982 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 13078 12968 13084 12980
rect 12483 12940 13084 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 13078 12928 13084 12940
rect 13136 12968 13142 12980
rect 15565 12971 15623 12977
rect 13136 12940 14872 12968
rect 13136 12928 13142 12940
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 11931 12872 14228 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 14200 12844 14228 12872
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 10962 12832 10968 12844
rect 1903 12804 10968 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12912 12764 12940 12795
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 13412 12804 13553 12832
rect 13412 12792 13418 12804
rect 13541 12801 13553 12804
rect 13587 12801 13599 12835
rect 14182 12832 14188 12844
rect 14143 12804 14188 12832
rect 13541 12795 13599 12801
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 14844 12841 14872 12940
rect 15565 12937 15577 12971
rect 15611 12968 15623 12971
rect 15611 12940 18920 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 14921 12903 14979 12909
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 17681 12903 17739 12909
rect 17681 12900 17693 12903
rect 14967 12872 17693 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 17681 12869 17693 12872
rect 17727 12869 17739 12903
rect 17681 12863 17739 12869
rect 17954 12860 17960 12912
rect 18012 12900 18018 12912
rect 18892 12909 18920 12940
rect 22554 12928 22560 12980
rect 22612 12968 22618 12980
rect 22612 12940 24624 12968
rect 22612 12928 22618 12940
rect 18785 12903 18843 12909
rect 18785 12900 18797 12903
rect 18012 12872 18797 12900
rect 18012 12860 18018 12872
rect 18785 12869 18797 12872
rect 18831 12869 18843 12903
rect 18785 12863 18843 12869
rect 18877 12903 18935 12909
rect 18877 12869 18889 12903
rect 18923 12869 18935 12903
rect 18877 12863 18935 12869
rect 18966 12860 18972 12912
rect 19024 12900 19030 12912
rect 19518 12900 19524 12912
rect 19024 12872 19524 12900
rect 19024 12860 19030 12872
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 21085 12903 21143 12909
rect 19812 12872 20944 12900
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15470 12832 15476 12844
rect 14875 12804 15476 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 15620 12804 16129 12832
rect 15620 12792 15626 12804
rect 16117 12801 16129 12804
rect 16163 12832 16175 12835
rect 16390 12832 16396 12844
rect 16163 12804 16396 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17402 12832 17408 12844
rect 17083 12804 17408 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 14366 12764 14372 12776
rect 12912 12736 14372 12764
rect 14366 12724 14372 12736
rect 14424 12764 14430 12776
rect 14424 12736 15608 12764
rect 14424 12724 14430 12736
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12696 13047 12699
rect 14182 12696 14188 12708
rect 13035 12668 14188 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 14277 12699 14335 12705
rect 14277 12665 14289 12699
rect 14323 12696 14335 12699
rect 15470 12696 15476 12708
rect 14323 12668 15476 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 15580 12696 15608 12736
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 17589 12767 17647 12773
rect 17589 12764 17601 12767
rect 16816 12736 17601 12764
rect 16816 12724 16822 12736
rect 17589 12733 17601 12736
rect 17635 12733 17647 12767
rect 17589 12727 17647 12733
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 19812 12764 19840 12872
rect 20070 12832 20076 12844
rect 20031 12804 20076 12832
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 20530 12832 20536 12844
rect 20491 12804 20536 12832
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 18279 12736 19840 12764
rect 19889 12767 19947 12773
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20254 12764 20260 12776
rect 19935 12736 20260 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20806 12764 20812 12776
rect 20364 12736 20812 12764
rect 17126 12696 17132 12708
rect 15580 12668 17132 12696
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 19337 12699 19395 12705
rect 19337 12665 19349 12699
rect 19383 12696 19395 12699
rect 20364 12696 20392 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 20916 12764 20944 12872
rect 21085 12869 21097 12903
rect 21131 12900 21143 12903
rect 22189 12903 22247 12909
rect 22189 12900 22201 12903
rect 21131 12872 22201 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 22189 12869 22201 12872
rect 22235 12869 22247 12903
rect 22189 12863 22247 12869
rect 22278 12860 22284 12912
rect 22336 12900 22342 12912
rect 24596 12909 24624 12940
rect 26418 12928 26424 12980
rect 26476 12968 26482 12980
rect 27522 12968 27528 12980
rect 26476 12940 27528 12968
rect 26476 12928 26482 12940
rect 27522 12928 27528 12940
rect 27580 12928 27586 12980
rect 28994 12968 29000 12980
rect 27724 12940 29000 12968
rect 23753 12903 23811 12909
rect 23753 12900 23765 12903
rect 22336 12872 23765 12900
rect 22336 12860 22342 12872
rect 23753 12869 23765 12872
rect 23799 12869 23811 12903
rect 23753 12863 23811 12869
rect 24581 12903 24639 12909
rect 24581 12869 24593 12903
rect 24627 12869 24639 12903
rect 25590 12900 25596 12912
rect 25551 12872 25596 12900
rect 24581 12863 24639 12869
rect 25590 12860 25596 12872
rect 25648 12860 25654 12912
rect 27724 12909 27752 12940
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 29086 12928 29092 12980
rect 29144 12968 29150 12980
rect 29641 12971 29699 12977
rect 29641 12968 29653 12971
rect 29144 12940 29653 12968
rect 29144 12928 29150 12940
rect 29641 12937 29653 12940
rect 29687 12937 29699 12971
rect 29641 12931 29699 12937
rect 30374 12928 30380 12980
rect 30432 12928 30438 12980
rect 30926 12968 30932 12980
rect 30887 12940 30932 12968
rect 30926 12928 30932 12940
rect 30984 12928 30990 12980
rect 38010 12968 38016 12980
rect 35866 12940 38016 12968
rect 26145 12903 26203 12909
rect 26145 12869 26157 12903
rect 26191 12900 26203 12903
rect 27716 12903 27774 12909
rect 26191 12872 27200 12900
rect 26191 12869 26203 12872
rect 26145 12863 26203 12869
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21174 12832 21180 12844
rect 21039 12804 21180 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 21174 12792 21180 12804
rect 21232 12832 21238 12844
rect 21450 12832 21456 12844
rect 21232 12804 21456 12832
rect 21232 12792 21238 12804
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 22097 12767 22155 12773
rect 20916 12736 22048 12764
rect 21174 12696 21180 12708
rect 19383 12668 20392 12696
rect 20456 12668 21180 12696
rect 19383 12665 19395 12668
rect 19337 12659 19395 12665
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 13630 12628 13636 12640
rect 13591 12600 13636 12628
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 15930 12628 15936 12640
rect 15344 12600 15936 12628
rect 15344 12588 15350 12600
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16209 12631 16267 12637
rect 16209 12597 16221 12631
rect 16255 12628 16267 12631
rect 16482 12628 16488 12640
rect 16255 12600 16488 12628
rect 16255 12597 16267 12600
rect 16209 12591 16267 12597
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 16945 12631 17003 12637
rect 16945 12597 16957 12631
rect 16991 12628 17003 12631
rect 20456 12628 20484 12668
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 22020 12696 22048 12736
rect 22097 12733 22109 12767
rect 22143 12764 22155 12767
rect 22186 12764 22192 12776
rect 22143 12736 22192 12764
rect 22143 12733 22155 12736
rect 22097 12727 22155 12733
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 22738 12764 22744 12776
rect 22699 12736 22744 12764
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 23845 12767 23903 12773
rect 23216 12736 23796 12764
rect 23216 12696 23244 12736
rect 22020 12668 23244 12696
rect 23293 12699 23351 12705
rect 23293 12665 23305 12699
rect 23339 12665 23351 12699
rect 23768 12696 23796 12736
rect 23845 12733 23857 12767
rect 23891 12764 23903 12767
rect 24118 12764 24124 12776
rect 23891 12736 24124 12764
rect 23891 12733 23903 12736
rect 23845 12727 23903 12733
rect 24118 12724 24124 12736
rect 24176 12724 24182 12776
rect 24486 12764 24492 12776
rect 24447 12736 24492 12764
rect 24486 12724 24492 12736
rect 24544 12724 24550 12776
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12733 24823 12767
rect 24765 12727 24823 12733
rect 26237 12767 26295 12773
rect 26237 12733 26249 12767
rect 26283 12764 26295 12767
rect 26510 12764 26516 12776
rect 26283 12736 26516 12764
rect 26283 12733 26295 12736
rect 26237 12727 26295 12733
rect 24780 12696 24808 12727
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 27172 12764 27200 12872
rect 27716 12869 27728 12903
rect 27762 12869 27774 12903
rect 28442 12900 28448 12912
rect 28403 12872 28448 12900
rect 27716 12863 27774 12869
rect 28442 12860 28448 12872
rect 28500 12860 28506 12912
rect 28537 12903 28595 12909
rect 28537 12869 28549 12903
rect 28583 12900 28595 12903
rect 29822 12900 29828 12912
rect 28583 12872 29828 12900
rect 28583 12869 28595 12872
rect 28537 12863 28595 12869
rect 29822 12860 29828 12872
rect 29880 12860 29886 12912
rect 30392 12900 30420 12928
rect 31294 12900 31300 12912
rect 30392 12872 31300 12900
rect 29730 12832 29736 12844
rect 29691 12804 29736 12832
rect 29730 12792 29736 12804
rect 29788 12792 29794 12844
rect 30392 12841 30420 12872
rect 31294 12860 31300 12872
rect 31352 12860 31358 12912
rect 35866 12900 35894 12940
rect 38010 12928 38016 12940
rect 38068 12928 38074 12980
rect 31496 12872 35894 12900
rect 30377 12835 30435 12841
rect 30377 12801 30389 12835
rect 30423 12801 30435 12835
rect 30377 12795 30435 12801
rect 31021 12835 31079 12841
rect 31021 12801 31033 12835
rect 31067 12832 31079 12835
rect 31202 12832 31208 12844
rect 31067 12804 31208 12832
rect 31067 12801 31079 12804
rect 31021 12795 31079 12801
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 27172 12736 27752 12764
rect 27249 12699 27307 12705
rect 27249 12696 27261 12699
rect 23768 12668 27261 12696
rect 23293 12659 23351 12665
rect 27249 12665 27261 12668
rect 27295 12696 27307 12699
rect 27614 12696 27620 12708
rect 27295 12668 27620 12696
rect 27295 12665 27307 12668
rect 27249 12659 27307 12665
rect 16991 12600 20484 12628
rect 16991 12597 17003 12600
rect 16945 12591 17003 12597
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 23308 12628 23336 12659
rect 27614 12656 27620 12668
rect 27672 12656 27678 12708
rect 27724 12696 27752 12736
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28166 12764 28172 12776
rect 27856 12736 28172 12764
rect 27856 12724 27862 12736
rect 28166 12724 28172 12736
rect 28224 12724 28230 12776
rect 28810 12764 28816 12776
rect 28771 12736 28816 12764
rect 28810 12724 28816 12736
rect 28868 12724 28874 12776
rect 29454 12764 29460 12776
rect 28920 12736 29460 12764
rect 28920 12696 28948 12736
rect 29454 12724 29460 12736
rect 29512 12724 29518 12776
rect 29748 12764 29776 12792
rect 31496 12773 31524 12872
rect 33226 12832 33232 12844
rect 33187 12804 33232 12832
rect 33226 12792 33232 12804
rect 33284 12792 33290 12844
rect 31481 12767 31539 12773
rect 31481 12764 31493 12767
rect 29748 12736 31493 12764
rect 31481 12733 31493 12736
rect 31527 12733 31539 12767
rect 31481 12727 31539 12733
rect 30285 12699 30343 12705
rect 30285 12696 30297 12699
rect 27724 12668 28948 12696
rect 29104 12668 30297 12696
rect 21140 12600 23336 12628
rect 21140 12588 21146 12600
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 24670 12628 24676 12640
rect 23532 12600 24676 12628
rect 23532 12588 23538 12600
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 27522 12588 27528 12640
rect 27580 12628 27586 12640
rect 29104 12628 29132 12668
rect 30285 12665 30297 12668
rect 30331 12665 30343 12699
rect 30285 12659 30343 12665
rect 27580 12600 29132 12628
rect 27580 12588 27586 12600
rect 30190 12588 30196 12640
rect 30248 12628 30254 12640
rect 33321 12631 33379 12637
rect 33321 12628 33333 12631
rect 30248 12600 33333 12628
rect 30248 12588 30254 12600
rect 33321 12597 33333 12600
rect 33367 12597 33379 12631
rect 33321 12591 33379 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 13078 12424 13084 12436
rect 13039 12396 13084 12424
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 16482 12384 16488 12436
rect 16540 12424 16546 12436
rect 16540 12396 17356 12424
rect 16540 12384 16546 12396
rect 13633 12359 13691 12365
rect 13633 12325 13645 12359
rect 13679 12356 13691 12359
rect 16850 12356 16856 12368
rect 13679 12328 16856 12356
rect 13679 12325 13691 12328
rect 13633 12319 13691 12325
rect 16850 12316 16856 12328
rect 16908 12316 16914 12368
rect 17328 12356 17356 12396
rect 17402 12384 17408 12436
rect 17460 12424 17466 12436
rect 18322 12424 18328 12436
rect 17460 12396 18328 12424
rect 17460 12384 17466 12396
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 21082 12424 21088 12436
rect 18656 12396 21088 12424
rect 18656 12384 18662 12396
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 21726 12424 21732 12436
rect 21600 12396 21732 12424
rect 21600 12384 21606 12396
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 29638 12424 29644 12436
rect 26914 12396 29644 12424
rect 18966 12356 18972 12368
rect 17328 12328 18972 12356
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 20441 12359 20499 12365
rect 20441 12325 20453 12359
rect 20487 12356 20499 12359
rect 22738 12356 22744 12368
rect 20487 12328 22744 12356
rect 20487 12325 20499 12328
rect 20441 12319 20499 12325
rect 22738 12316 22744 12328
rect 22796 12356 22802 12368
rect 22833 12359 22891 12365
rect 22833 12356 22845 12359
rect 22796 12328 22845 12356
rect 22796 12316 22802 12328
rect 22833 12325 22845 12328
rect 22879 12356 22891 12359
rect 25958 12356 25964 12368
rect 22879 12328 25964 12356
rect 22879 12325 22891 12328
rect 22833 12319 22891 12325
rect 25958 12316 25964 12328
rect 26016 12316 26022 12368
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 15068 12260 16589 12288
rect 15068 12248 15074 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 18230 12288 18236 12300
rect 18191 12260 18236 12288
rect 16577 12251 16635 12257
rect 18230 12248 18236 12260
rect 18288 12288 18294 12300
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 18288 12260 19901 12288
rect 18288 12248 18294 12260
rect 19889 12257 19901 12260
rect 19935 12257 19947 12291
rect 21542 12288 21548 12300
rect 19889 12251 19947 12257
rect 20548 12260 21548 12288
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 12575 12192 13553 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 13541 12189 13553 12192
rect 13587 12220 13599 12223
rect 14090 12220 14096 12232
rect 13587 12192 14096 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14642 12220 14648 12232
rect 14603 12192 14648 12220
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 15378 12152 15384 12164
rect 13780 12124 15384 12152
rect 13780 12112 13786 12124
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 15470 12112 15476 12164
rect 15528 12152 15534 12164
rect 16025 12155 16083 12161
rect 15528 12124 15573 12152
rect 15528 12112 15534 12124
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16298 12152 16304 12164
rect 16071 12124 16304 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 16666 12112 16672 12164
rect 16724 12152 16730 12164
rect 17221 12155 17279 12161
rect 16724 12124 16769 12152
rect 16724 12112 16730 12124
rect 17221 12121 17233 12155
rect 17267 12152 17279 12155
rect 17310 12152 17316 12164
rect 17267 12124 17316 12152
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 18325 12155 18383 12161
rect 18325 12121 18337 12155
rect 18371 12121 18383 12155
rect 18325 12115 18383 12121
rect 18877 12155 18935 12161
rect 18877 12121 18889 12155
rect 18923 12121 18935 12155
rect 18877 12115 18935 12121
rect 14737 12087 14795 12093
rect 14737 12053 14749 12087
rect 14783 12084 14795 12087
rect 18340 12084 18368 12115
rect 14783 12056 18368 12084
rect 18892 12084 18920 12115
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 19981 12155 20039 12161
rect 19981 12152 19993 12155
rect 19024 12124 19993 12152
rect 19024 12112 19030 12124
rect 19981 12121 19993 12124
rect 20027 12121 20039 12155
rect 19981 12115 20039 12121
rect 20162 12084 20168 12096
rect 18892 12056 20168 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 20162 12044 20168 12056
rect 20220 12084 20226 12096
rect 20548 12084 20576 12260
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 22002 12248 22008 12300
rect 22060 12288 22066 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 22060 12260 22293 12288
rect 22060 12248 22066 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 23290 12248 23296 12300
rect 23348 12288 23354 12300
rect 23385 12291 23443 12297
rect 23385 12288 23397 12291
rect 23348 12260 23397 12288
rect 23348 12248 23354 12260
rect 23385 12257 23397 12260
rect 23431 12257 23443 12291
rect 23385 12251 23443 12257
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25406 12288 25412 12300
rect 25271 12260 25412 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 25406 12248 25412 12260
rect 25464 12248 25470 12300
rect 26418 12288 26424 12300
rect 26379 12260 26424 12288
rect 26418 12248 26424 12260
rect 26476 12248 26482 12300
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 23624 12192 24593 12220
rect 23624 12180 23630 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 21085 12155 21143 12161
rect 21085 12121 21097 12155
rect 21131 12121 21143 12155
rect 21085 12115 21143 12121
rect 20220 12056 20576 12084
rect 21100 12084 21128 12115
rect 21174 12112 21180 12164
rect 21232 12152 21238 12164
rect 21232 12124 21277 12152
rect 21232 12112 21238 12124
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 21600 12124 21741 12152
rect 21600 12112 21606 12124
rect 21729 12121 21741 12124
rect 21775 12152 21787 12155
rect 22373 12155 22431 12161
rect 21775 12124 22324 12152
rect 21775 12121 21787 12124
rect 21729 12115 21787 12121
rect 21358 12084 21364 12096
rect 21100 12056 21364 12084
rect 20220 12044 20226 12056
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 22296 12084 22324 12124
rect 22373 12121 22385 12155
rect 22419 12152 22431 12155
rect 23842 12152 23848 12164
rect 22419 12124 23848 12152
rect 22419 12121 22431 12124
rect 22373 12115 22431 12121
rect 23842 12112 23848 12124
rect 23900 12112 23906 12164
rect 25133 12155 25191 12161
rect 25133 12121 25145 12155
rect 25179 12121 25191 12155
rect 25133 12115 25191 12121
rect 22830 12084 22836 12096
rect 22296 12056 22836 12084
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 25148 12084 25176 12115
rect 25774 12112 25780 12164
rect 25832 12152 25838 12164
rect 26329 12155 26387 12161
rect 25832 12124 25877 12152
rect 25832 12112 25838 12124
rect 26329 12121 26341 12155
rect 26375 12152 26387 12155
rect 26914 12152 26942 12396
rect 29638 12384 29644 12396
rect 29696 12384 29702 12436
rect 27062 12356 27068 12368
rect 27023 12328 27068 12356
rect 27062 12316 27068 12328
rect 27120 12316 27126 12368
rect 28810 12356 28816 12368
rect 28771 12328 28816 12356
rect 28810 12316 28816 12328
rect 28868 12316 28874 12368
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 27617 12291 27675 12297
rect 27617 12288 27629 12291
rect 27396 12260 27629 12288
rect 27396 12248 27402 12260
rect 27617 12257 27629 12260
rect 27663 12257 27675 12291
rect 27617 12251 27675 12257
rect 28718 12248 28724 12300
rect 28776 12288 28782 12300
rect 30469 12291 30527 12297
rect 30469 12288 30481 12291
rect 28776 12260 30481 12288
rect 28776 12248 28782 12260
rect 30469 12257 30481 12260
rect 30515 12257 30527 12291
rect 30469 12251 30527 12257
rect 29730 12180 29736 12232
rect 29788 12220 29794 12232
rect 29917 12223 29975 12229
rect 29917 12220 29929 12223
rect 29788 12192 29929 12220
rect 29788 12180 29794 12192
rect 29917 12189 29929 12192
rect 29963 12220 29975 12223
rect 29963 12192 30052 12220
rect 29963 12189 29975 12192
rect 29917 12183 29975 12189
rect 27522 12152 27528 12164
rect 26375 12124 26942 12152
rect 27483 12124 27528 12152
rect 26375 12121 26387 12124
rect 26329 12115 26387 12121
rect 27522 12112 27528 12124
rect 27580 12112 27586 12164
rect 27614 12112 27620 12164
rect 27672 12152 27678 12164
rect 28261 12155 28319 12161
rect 28261 12152 28273 12155
rect 27672 12124 28273 12152
rect 27672 12112 27678 12124
rect 28261 12121 28273 12124
rect 28307 12121 28319 12155
rect 28261 12115 28319 12121
rect 28353 12155 28411 12161
rect 28353 12121 28365 12155
rect 28399 12152 28411 12155
rect 29638 12152 29644 12164
rect 28399 12124 29644 12152
rect 28399 12121 28411 12124
rect 28353 12115 28411 12121
rect 29638 12112 29644 12124
rect 29696 12112 29702 12164
rect 30024 12152 30052 12192
rect 30190 12180 30196 12232
rect 30248 12220 30254 12232
rect 30377 12223 30435 12229
rect 30377 12220 30389 12223
rect 30248 12192 30389 12220
rect 30248 12180 30254 12192
rect 30377 12189 30389 12192
rect 30423 12189 30435 12223
rect 31018 12220 31024 12232
rect 30979 12192 31024 12220
rect 30377 12183 30435 12189
rect 31018 12180 31024 12192
rect 31076 12180 31082 12232
rect 31110 12180 31116 12232
rect 31168 12220 31174 12232
rect 31168 12192 31213 12220
rect 31168 12180 31174 12192
rect 30558 12152 30564 12164
rect 30024 12124 30564 12152
rect 30558 12112 30564 12124
rect 30616 12152 30622 12164
rect 32217 12155 32275 12161
rect 32217 12152 32229 12155
rect 30616 12124 32229 12152
rect 30616 12112 30622 12124
rect 32217 12121 32229 12124
rect 32263 12121 32275 12155
rect 32217 12115 32275 12121
rect 27430 12084 27436 12096
rect 25148 12056 27436 12084
rect 27430 12044 27436 12056
rect 27488 12044 27494 12096
rect 27706 12044 27712 12096
rect 27764 12084 27770 12096
rect 29825 12087 29883 12093
rect 29825 12084 29837 12087
rect 27764 12056 29837 12084
rect 27764 12044 27770 12056
rect 29825 12053 29837 12056
rect 29871 12053 29883 12087
rect 29825 12047 29883 12053
rect 31202 12044 31208 12096
rect 31260 12084 31266 12096
rect 31478 12084 31484 12096
rect 31260 12056 31484 12084
rect 31260 12044 31266 12056
rect 31478 12044 31484 12056
rect 31536 12044 31542 12096
rect 31662 12084 31668 12096
rect 31623 12056 31668 12084
rect 31662 12044 31668 12056
rect 31720 12044 31726 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 13722 11880 13728 11892
rect 13683 11852 13728 11880
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 15013 11883 15071 11889
rect 15013 11849 15025 11883
rect 15059 11880 15071 11883
rect 15059 11852 19012 11880
rect 15059 11849 15071 11852
rect 15013 11843 15071 11849
rect 11974 11812 11980 11824
rect 11887 11784 11980 11812
rect 11974 11772 11980 11784
rect 12032 11812 12038 11824
rect 14369 11815 14427 11821
rect 12032 11784 13492 11812
rect 12032 11772 12038 11784
rect 13464 11756 13492 11784
rect 14369 11781 14381 11815
rect 14415 11812 14427 11815
rect 15749 11815 15807 11821
rect 15749 11812 15761 11815
rect 14415 11784 15761 11812
rect 14415 11781 14427 11784
rect 14369 11775 14427 11781
rect 15749 11781 15761 11784
rect 15795 11781 15807 11815
rect 16298 11812 16304 11824
rect 16259 11784 16304 11812
rect 15749 11775 15807 11781
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 17402 11812 17408 11824
rect 17236 11784 17408 11812
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13188 11676 13216 11707
rect 13446 11704 13452 11756
rect 13504 11744 13510 11756
rect 13633 11747 13691 11753
rect 13633 11744 13645 11747
rect 13504 11716 13645 11744
rect 13504 11704 13510 11716
rect 13633 11713 13645 11716
rect 13679 11713 13691 11747
rect 14458 11744 14464 11756
rect 14419 11716 14464 11744
rect 13633 11707 13691 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11742 14979 11747
rect 17129 11747 17187 11753
rect 14967 11714 15056 11742
rect 14967 11713 14979 11714
rect 14921 11707 14979 11713
rect 14642 11676 14648 11688
rect 13188 11648 14648 11676
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 12529 11611 12587 11617
rect 12529 11577 12541 11611
rect 12575 11608 12587 11611
rect 15028 11608 15056 11714
rect 17129 11713 17141 11747
rect 17175 11742 17187 11747
rect 17236 11742 17264 11784
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 17770 11812 17776 11824
rect 17731 11784 17776 11812
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 18984 11821 19012 11852
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 21542 11880 21548 11892
rect 20312 11852 21548 11880
rect 20312 11840 20318 11852
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 23842 11840 23848 11892
rect 23900 11880 23906 11892
rect 24305 11883 24363 11889
rect 24305 11880 24317 11883
rect 23900 11852 24317 11880
rect 23900 11840 23906 11852
rect 24305 11849 24317 11852
rect 24351 11849 24363 11883
rect 24305 11843 24363 11849
rect 26050 11840 26056 11892
rect 26108 11880 26114 11892
rect 26326 11880 26332 11892
rect 26108 11852 26332 11880
rect 26108 11840 26114 11852
rect 26326 11840 26332 11852
rect 26384 11840 26390 11892
rect 31110 11880 31116 11892
rect 27172 11852 28488 11880
rect 27172 11824 27200 11852
rect 18969 11815 19027 11821
rect 18969 11781 18981 11815
rect 19015 11781 19027 11815
rect 18969 11775 19027 11781
rect 19150 11772 19156 11824
rect 19208 11812 19214 11824
rect 20346 11812 20352 11824
rect 19208 11784 20352 11812
rect 19208 11772 19214 11784
rect 20346 11772 20352 11784
rect 20404 11772 20410 11824
rect 21269 11815 21327 11821
rect 21269 11781 21281 11815
rect 21315 11812 21327 11815
rect 22094 11812 22100 11824
rect 21315 11784 22100 11812
rect 21315 11781 21327 11784
rect 21269 11775 21327 11781
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 22738 11772 22744 11824
rect 22796 11772 22802 11824
rect 23382 11772 23388 11824
rect 23440 11812 23446 11824
rect 23477 11815 23535 11821
rect 23477 11812 23489 11815
rect 23440 11784 23489 11812
rect 23440 11772 23446 11784
rect 23477 11781 23489 11784
rect 23523 11781 23535 11815
rect 23477 11775 23535 11781
rect 24578 11772 24584 11824
rect 24636 11812 24642 11824
rect 27154 11812 27160 11824
rect 24636 11784 25162 11812
rect 27115 11784 27160 11812
rect 24636 11772 24642 11784
rect 27154 11772 27160 11784
rect 27212 11772 27218 11824
rect 28460 11821 28488 11852
rect 28552 11852 31116 11880
rect 28552 11821 28580 11852
rect 31110 11840 31116 11852
rect 31168 11840 31174 11892
rect 31570 11880 31576 11892
rect 31531 11852 31576 11880
rect 31570 11840 31576 11852
rect 31628 11840 31634 11892
rect 27709 11815 27767 11821
rect 27709 11781 27721 11815
rect 27755 11812 27767 11815
rect 28445 11815 28503 11821
rect 27755 11784 28304 11812
rect 27755 11781 27767 11784
rect 27709 11775 27767 11781
rect 24394 11744 24400 11756
rect 17175 11714 17264 11742
rect 24355 11716 24400 11744
rect 17175 11713 17187 11714
rect 17129 11707 17187 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11744 26663 11747
rect 27062 11744 27068 11756
rect 26651 11716 27068 11744
rect 26651 11713 26663 11716
rect 26605 11707 26663 11713
rect 27062 11704 27068 11716
rect 27120 11704 27126 11756
rect 15654 11676 15660 11688
rect 15615 11648 15660 11676
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 17402 11676 17408 11688
rect 15764 11648 17408 11676
rect 15764 11608 15792 11648
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11676 17739 11679
rect 17954 11676 17960 11688
rect 17727 11648 17960 11676
rect 17727 11645 17739 11648
rect 17681 11639 17739 11645
rect 12575 11580 15792 11608
rect 12575 11577 12587 11580
rect 12529 11571 12587 11577
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 17696 11608 17724 11639
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 18966 11676 18972 11688
rect 18923 11648 18972 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 19426 11676 19432 11688
rect 19387 11648 19432 11676
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 21085 11679 21143 11685
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 21174 11676 21180 11688
rect 21131 11648 21180 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 23753 11679 23811 11685
rect 21416 11648 21509 11676
rect 21416 11636 21422 11648
rect 23753 11645 23765 11679
rect 23799 11676 23811 11679
rect 23842 11676 23848 11688
rect 23799 11648 23848 11676
rect 23799 11645 23811 11648
rect 23753 11639 23811 11645
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11676 24915 11679
rect 25038 11676 25044 11688
rect 24903 11648 25044 11676
rect 24903 11645 24915 11648
rect 24857 11639 24915 11645
rect 25038 11636 25044 11648
rect 25096 11676 25102 11688
rect 27798 11676 27804 11688
rect 25096 11648 27292 11676
rect 27759 11648 27804 11676
rect 25096 11636 25102 11648
rect 16632 11580 17724 11608
rect 18233 11611 18291 11617
rect 16632 11568 16638 11580
rect 18233 11577 18245 11611
rect 18279 11608 18291 11611
rect 18598 11608 18604 11620
rect 18279 11580 18604 11608
rect 18279 11577 18291 11580
rect 18233 11571 18291 11577
rect 18598 11568 18604 11580
rect 18656 11568 18662 11620
rect 20714 11608 20720 11620
rect 18800 11580 20720 11608
rect 13081 11543 13139 11549
rect 13081 11509 13093 11543
rect 13127 11540 13139 11543
rect 15102 11540 15108 11552
rect 13127 11512 15108 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11540 17095 11543
rect 18800 11540 18828 11580
rect 20714 11568 20720 11580
rect 20772 11568 20778 11620
rect 21376 11608 21404 11636
rect 27264 11620 27292 11648
rect 27798 11636 27804 11648
rect 27856 11636 27862 11688
rect 21376 11580 22140 11608
rect 17083 11512 18828 11540
rect 17083 11509 17095 11512
rect 17037 11503 17095 11509
rect 18874 11500 18880 11552
rect 18932 11540 18938 11552
rect 21358 11540 21364 11552
rect 18932 11512 21364 11540
rect 18932 11500 18938 11512
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21542 11500 21548 11552
rect 21600 11540 21606 11552
rect 22005 11543 22063 11549
rect 22005 11540 22017 11543
rect 21600 11512 22017 11540
rect 21600 11500 21606 11512
rect 22005 11509 22017 11512
rect 22051 11509 22063 11543
rect 22112 11540 22140 11580
rect 27246 11568 27252 11620
rect 27304 11568 27310 11620
rect 28276 11608 28304 11784
rect 28445 11781 28457 11815
rect 28491 11781 28503 11815
rect 28445 11775 28503 11781
rect 28537 11815 28595 11821
rect 28537 11781 28549 11815
rect 28583 11781 28595 11815
rect 28537 11775 28595 11781
rect 29089 11815 29147 11821
rect 29089 11781 29101 11815
rect 29135 11812 29147 11815
rect 29178 11812 29184 11824
rect 29135 11784 29184 11812
rect 29135 11781 29147 11784
rect 29089 11775 29147 11781
rect 29178 11772 29184 11784
rect 29236 11772 29242 11824
rect 29454 11772 29460 11824
rect 29512 11812 29518 11824
rect 29641 11815 29699 11821
rect 29641 11812 29653 11815
rect 29512 11784 29653 11812
rect 29512 11772 29518 11784
rect 29641 11781 29653 11784
rect 29687 11781 29699 11815
rect 32306 11812 32312 11824
rect 29641 11775 29699 11781
rect 30392 11784 32312 11812
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11744 29607 11747
rect 29730 11744 29736 11756
rect 29595 11716 29736 11744
rect 29595 11713 29607 11716
rect 29549 11707 29607 11713
rect 29730 11704 29736 11716
rect 29788 11704 29794 11756
rect 30392 11753 30420 11784
rect 32306 11772 32312 11784
rect 32364 11772 32370 11824
rect 30377 11747 30435 11753
rect 30377 11713 30389 11747
rect 30423 11713 30435 11747
rect 30926 11744 30932 11756
rect 30887 11716 30932 11744
rect 30377 11707 30435 11713
rect 30926 11704 30932 11716
rect 30984 11704 30990 11756
rect 31021 11747 31079 11753
rect 31021 11713 31033 11747
rect 31067 11744 31079 11747
rect 31202 11744 31208 11756
rect 31067 11716 31208 11744
rect 31067 11713 31079 11716
rect 31021 11707 31079 11713
rect 31202 11704 31208 11716
rect 31260 11704 31266 11756
rect 31665 11747 31723 11753
rect 31665 11713 31677 11747
rect 31711 11713 31723 11747
rect 31665 11707 31723 11713
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11744 37611 11747
rect 38194 11744 38200 11756
rect 37599 11716 38200 11744
rect 37599 11713 37611 11716
rect 37553 11707 37611 11713
rect 28442 11636 28448 11688
rect 28500 11676 28506 11688
rect 30190 11676 30196 11688
rect 28500 11648 30196 11676
rect 28500 11636 28506 11648
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 31110 11636 31116 11688
rect 31168 11676 31174 11688
rect 31680 11676 31708 11707
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 31168 11648 31708 11676
rect 31168 11636 31174 11648
rect 30285 11611 30343 11617
rect 30285 11608 30297 11611
rect 28276 11580 30297 11608
rect 30285 11577 30297 11580
rect 30331 11577 30343 11611
rect 38013 11611 38071 11617
rect 38013 11608 38025 11611
rect 30285 11571 30343 11577
rect 31726 11580 38025 11608
rect 23014 11540 23020 11552
rect 22112 11512 23020 11540
rect 22005 11503 22063 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 26347 11543 26405 11549
rect 26347 11509 26359 11543
rect 26393 11540 26405 11543
rect 28258 11540 28264 11552
rect 26393 11512 28264 11540
rect 26393 11509 26405 11512
rect 26347 11503 26405 11509
rect 28258 11500 28264 11512
rect 28316 11500 28322 11552
rect 29086 11500 29092 11552
rect 29144 11540 29150 11552
rect 31726 11540 31754 11580
rect 38013 11577 38025 11580
rect 38059 11577 38071 11611
rect 38013 11571 38071 11577
rect 32306 11540 32312 11552
rect 29144 11512 31754 11540
rect 32267 11512 32312 11540
rect 29144 11500 29150 11512
rect 32306 11500 32312 11512
rect 32364 11500 32370 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 8996 11308 12173 11336
rect 8996 11296 9002 11308
rect 12161 11305 12173 11308
rect 12207 11305 12219 11339
rect 12161 11299 12219 11305
rect 14369 11339 14427 11345
rect 14369 11305 14381 11339
rect 14415 11336 14427 11339
rect 17770 11336 17776 11348
rect 14415 11308 17776 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 12176 11200 12204 11299
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18141 11339 18199 11345
rect 18141 11336 18153 11339
rect 18104 11308 18153 11336
rect 18104 11296 18110 11308
rect 18141 11305 18153 11308
rect 18187 11305 18199 11339
rect 18141 11299 18199 11305
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 23566 11336 23572 11348
rect 19392 11308 23572 11336
rect 19392 11296 19398 11308
rect 23566 11296 23572 11308
rect 23624 11296 23630 11348
rect 27706 11336 27712 11348
rect 27667 11308 27712 11336
rect 27706 11296 27712 11308
rect 27764 11296 27770 11348
rect 27798 11296 27804 11348
rect 27856 11336 27862 11348
rect 27856 11308 28488 11336
rect 27856 11296 27862 11308
rect 14182 11228 14188 11280
rect 14240 11268 14246 11280
rect 17310 11268 17316 11280
rect 14240 11240 15792 11268
rect 17223 11240 17316 11268
rect 14240 11228 14246 11240
rect 12176 11172 13584 11200
rect 13556 11144 13584 11172
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15764 11209 15792 11240
rect 17310 11228 17316 11240
rect 17368 11268 17374 11280
rect 18966 11268 18972 11280
rect 17368 11240 18972 11268
rect 17368 11228 17374 11240
rect 18966 11228 18972 11240
rect 19024 11268 19030 11280
rect 20257 11271 20315 11277
rect 19024 11240 19840 11268
rect 19024 11228 19030 11240
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15436 11172 15577 11200
rect 15436 11160 15442 11172
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 16758 11200 16764 11212
rect 15749 11163 15807 11169
rect 15856 11172 16764 11200
rect 12894 11132 12900 11144
rect 12855 11104 12900 11132
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13538 11132 13544 11144
rect 13499 11104 13544 11132
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14921 11135 14979 11141
rect 14921 11132 14933 11135
rect 14516 11104 14933 11132
rect 14516 11092 14522 11104
rect 14921 11101 14933 11104
rect 14967 11132 14979 11135
rect 15470 11132 15476 11144
rect 14967 11104 15476 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15856 11132 15884 11172
rect 16758 11160 16764 11172
rect 16816 11160 16822 11212
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 18598 11200 18604 11212
rect 17736 11172 18604 11200
rect 17736 11160 17742 11172
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18708 11172 19012 11200
rect 15764 11104 15884 11132
rect 18233 11135 18291 11141
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 15013 11067 15071 11073
rect 13679 11036 14964 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 12710 10996 12716 11008
rect 12671 10968 12716 10996
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 14936 10996 14964 11036
rect 15013 11033 15025 11067
rect 15059 11064 15071 11067
rect 15378 11064 15384 11076
rect 15059 11036 15384 11064
rect 15059 11033 15071 11036
rect 15013 11027 15071 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 15764 11064 15792 11104
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 18322 11132 18328 11144
rect 18279 11104 18328 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 15488 11036 15792 11064
rect 15488 10996 15516 11036
rect 16390 11024 16396 11076
rect 16448 11064 16454 11076
rect 16448 11036 16804 11064
rect 16448 11024 16454 11036
rect 16206 10996 16212 11008
rect 14936 10968 15516 10996
rect 16167 10968 16212 10996
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16776 10996 16804 11036
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 18708 11064 18736 11172
rect 18874 11132 18880 11144
rect 18835 11104 18880 11132
rect 18874 11092 18880 11104
rect 18932 11092 18938 11144
rect 18984 11132 19012 11172
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 19484 11172 19717 11200
rect 19484 11160 19490 11172
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 19812 11200 19840 11240
rect 20257 11237 20269 11271
rect 20303 11268 20315 11271
rect 20346 11268 20352 11280
rect 20303 11240 20352 11268
rect 20303 11237 20315 11240
rect 20257 11231 20315 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 20438 11228 20444 11280
rect 20496 11268 20502 11280
rect 22002 11268 22008 11280
rect 20496 11240 22008 11268
rect 20496 11228 20502 11240
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 22097 11271 22155 11277
rect 22097 11237 22109 11271
rect 22143 11268 22155 11271
rect 22554 11268 22560 11280
rect 22143 11240 22560 11268
rect 22143 11237 22155 11240
rect 22097 11231 22155 11237
rect 22554 11228 22560 11240
rect 22612 11228 22618 11280
rect 24673 11271 24731 11277
rect 24673 11268 24685 11271
rect 23768 11240 24685 11268
rect 23768 11200 23796 11240
rect 24673 11237 24685 11240
rect 24719 11237 24731 11271
rect 28353 11271 28411 11277
rect 28353 11268 28365 11271
rect 24673 11231 24731 11237
rect 27264 11240 28365 11268
rect 25961 11203 26019 11209
rect 19812 11172 23796 11200
rect 23860 11172 25636 11200
rect 19705 11163 19763 11169
rect 23860 11144 23888 11172
rect 19518 11132 19524 11144
rect 18984 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 20806 11132 20812 11144
rect 20767 11104 20812 11132
rect 20806 11092 20812 11104
rect 20864 11092 20870 11144
rect 23842 11092 23848 11144
rect 23900 11132 23906 11144
rect 25608 11132 25636 11172
rect 25961 11169 25973 11203
rect 26007 11200 26019 11203
rect 26234 11200 26240 11212
rect 26007 11172 26240 11200
rect 26007 11169 26019 11172
rect 25961 11163 26019 11169
rect 25976 11132 26004 11163
rect 26234 11160 26240 11172
rect 26292 11160 26298 11212
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 27264 11200 27292 11240
rect 28353 11237 28365 11240
rect 28399 11237 28411 11271
rect 28460 11268 28488 11308
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29825 11339 29883 11345
rect 29825 11336 29837 11339
rect 29052 11308 29837 11336
rect 29052 11296 29058 11308
rect 29825 11305 29837 11308
rect 29871 11305 29883 11339
rect 29825 11299 29883 11305
rect 29178 11268 29184 11280
rect 28460 11240 29184 11268
rect 28353 11231 28411 11237
rect 29178 11228 29184 11240
rect 29236 11268 29242 11280
rect 30466 11268 30472 11280
rect 29236 11240 30472 11268
rect 29236 11228 29242 11240
rect 30466 11228 30472 11240
rect 30524 11228 30530 11280
rect 33229 11271 33287 11277
rect 33229 11237 33241 11271
rect 33275 11268 33287 11271
rect 33502 11268 33508 11280
rect 33275 11240 33508 11268
rect 33275 11237 33287 11240
rect 33229 11231 33287 11237
rect 33502 11228 33508 11240
rect 33560 11228 33566 11280
rect 32398 11200 32404 11212
rect 26384 11172 27292 11200
rect 27356 11172 29132 11200
rect 26384 11160 26390 11172
rect 23900 11104 23945 11132
rect 25608 11104 26004 11132
rect 27356 11118 27384 11172
rect 29104 11132 29132 11172
rect 29288 11172 32404 11200
rect 29288 11132 29316 11172
rect 32398 11160 32404 11172
rect 32456 11160 32462 11212
rect 29104 11104 29316 11132
rect 23900 11092 23906 11104
rect 29730 11092 29736 11144
rect 29788 11132 29794 11144
rect 29914 11132 29920 11144
rect 29788 11104 29920 11132
rect 29788 11092 29794 11104
rect 29914 11092 29920 11104
rect 29972 11092 29978 11144
rect 30374 11132 30380 11144
rect 30335 11104 30380 11132
rect 30374 11092 30380 11104
rect 30432 11092 30438 11144
rect 33410 11132 33416 11144
rect 33371 11104 33416 11132
rect 33410 11092 33416 11104
rect 33468 11092 33474 11144
rect 16908 11036 16953 11064
rect 17052 11036 18736 11064
rect 18785 11067 18843 11073
rect 16908 11024 16914 11036
rect 17052 10996 17080 11036
rect 18785 11033 18797 11067
rect 18831 11064 18843 11067
rect 19797 11067 19855 11073
rect 18831 11036 19656 11064
rect 18831 11033 18843 11036
rect 18785 11027 18843 11033
rect 16776 10968 17080 10996
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 18598 10996 18604 11008
rect 17184 10968 18604 10996
rect 17184 10956 17190 10968
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 19628 10996 19656 11036
rect 19797 11033 19809 11067
rect 19843 11033 19855 11067
rect 19797 11027 19855 11033
rect 19812 10996 19840 11027
rect 20990 11024 20996 11076
rect 21048 11064 21054 11076
rect 21361 11067 21419 11073
rect 21361 11064 21373 11067
rect 21048 11036 21373 11064
rect 21048 11024 21054 11036
rect 21361 11033 21373 11036
rect 21407 11033 21419 11067
rect 21361 11027 21419 11033
rect 21453 11067 21511 11073
rect 21453 11033 21465 11067
rect 21499 11064 21511 11067
rect 21499 11036 22140 11064
rect 21499 11033 21511 11036
rect 21453 11027 21511 11033
rect 22112 11008 22140 11036
rect 22186 11024 22192 11076
rect 22244 11064 22250 11076
rect 22244 11036 22402 11064
rect 22244 11024 22250 11036
rect 23290 11024 23296 11076
rect 23348 11064 23354 11076
rect 23569 11067 23627 11073
rect 23569 11064 23581 11067
rect 23348 11036 23581 11064
rect 23348 11024 23354 11036
rect 23569 11033 23581 11036
rect 23615 11033 23627 11067
rect 25130 11064 25136 11076
rect 23569 11027 23627 11033
rect 23676 11036 24992 11064
rect 25091 11036 25136 11064
rect 19628 10968 19840 10996
rect 22094 10956 22100 11008
rect 22152 10956 22158 11008
rect 22830 10956 22836 11008
rect 22888 10996 22894 11008
rect 23676 10996 23704 11036
rect 22888 10968 23704 10996
rect 24964 10996 24992 11036
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25222 11024 25228 11076
rect 25280 11064 25286 11076
rect 26237 11067 26295 11073
rect 26237 11064 26249 11067
rect 25280 11036 25325 11064
rect 25976 11036 26249 11064
rect 25280 11024 25286 11036
rect 25976 10996 26004 11036
rect 26237 11033 26249 11036
rect 26283 11033 26295 11067
rect 26237 11027 26295 11033
rect 27522 11024 27528 11076
rect 27580 11064 27586 11076
rect 28813 11067 28871 11073
rect 28813 11064 28825 11067
rect 27580 11036 28825 11064
rect 27580 11024 27586 11036
rect 28813 11033 28825 11036
rect 28859 11033 28871 11067
rect 28813 11027 28871 11033
rect 28905 11067 28963 11073
rect 28905 11033 28917 11067
rect 28951 11064 28963 11067
rect 29178 11064 29184 11076
rect 28951 11036 29184 11064
rect 28951 11033 28963 11036
rect 28905 11027 28963 11033
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 30006 11024 30012 11076
rect 30064 11064 30070 11076
rect 31021 11067 31079 11073
rect 31021 11064 31033 11067
rect 30064 11036 31033 11064
rect 30064 11024 30070 11036
rect 31021 11033 31033 11036
rect 31067 11064 31079 11067
rect 31573 11067 31631 11073
rect 31573 11064 31585 11067
rect 31067 11036 31585 11064
rect 31067 11033 31079 11036
rect 31021 11027 31079 11033
rect 31573 11033 31585 11036
rect 31619 11064 31631 11067
rect 31662 11064 31668 11076
rect 31619 11036 31668 11064
rect 31619 11033 31631 11036
rect 31573 11027 31631 11033
rect 31662 11024 31668 11036
rect 31720 11064 31726 11076
rect 32125 11067 32183 11073
rect 32125 11064 32137 11067
rect 31720 11036 32137 11064
rect 31720 11024 31726 11036
rect 32125 11033 32137 11036
rect 32171 11033 32183 11067
rect 32125 11027 32183 11033
rect 24964 10968 26004 10996
rect 22888 10956 22894 10968
rect 26050 10956 26056 11008
rect 26108 10996 26114 11008
rect 30282 10996 30288 11008
rect 26108 10968 30288 10996
rect 26108 10956 26114 10968
rect 30282 10956 30288 10968
rect 30340 10956 30346 11008
rect 30466 10996 30472 11008
rect 30427 10968 30472 10996
rect 30466 10956 30472 10968
rect 30524 10956 30530 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 12345 10795 12403 10801
rect 12345 10761 12357 10795
rect 12391 10792 12403 10795
rect 12894 10792 12900 10804
rect 12391 10764 12900 10792
rect 12391 10761 12403 10764
rect 12345 10755 12403 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13262 10752 13268 10804
rect 13320 10792 13326 10804
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 13320 10764 13461 10792
rect 13320 10752 13326 10764
rect 13449 10761 13461 10764
rect 13495 10792 13507 10795
rect 16574 10792 16580 10804
rect 13495 10764 16580 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 22094 10792 22100 10804
rect 16991 10764 22100 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22204 10764 23428 10792
rect 12805 10727 12863 10733
rect 12805 10693 12817 10727
rect 12851 10724 12863 10727
rect 14274 10724 14280 10736
rect 12851 10696 14280 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 15378 10684 15384 10736
rect 15436 10724 15442 10736
rect 18877 10727 18935 10733
rect 18877 10724 18889 10727
rect 15436 10696 18889 10724
rect 15436 10684 15442 10696
rect 18877 10693 18889 10696
rect 18923 10693 18935 10727
rect 18877 10687 18935 10693
rect 20441 10727 20499 10733
rect 20441 10693 20453 10727
rect 20487 10724 20499 10727
rect 20806 10724 20812 10736
rect 20487 10696 20812 10724
rect 20487 10693 20499 10696
rect 20441 10687 20499 10693
rect 20806 10684 20812 10696
rect 20864 10684 20870 10736
rect 21266 10724 21272 10736
rect 21227 10696 21272 10724
rect 21266 10684 21272 10696
rect 21324 10684 21330 10736
rect 21450 10684 21456 10736
rect 21508 10724 21514 10736
rect 21634 10724 21640 10736
rect 21508 10696 21640 10724
rect 21508 10684 21514 10696
rect 21634 10684 21640 10696
rect 21692 10724 21698 10736
rect 22204 10724 22232 10764
rect 21692 10696 22232 10724
rect 23400 10724 23428 10764
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 23842 10792 23848 10804
rect 23532 10764 23848 10792
rect 23532 10752 23538 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 24026 10752 24032 10804
rect 24084 10792 24090 10804
rect 26513 10795 26571 10801
rect 24084 10764 26464 10792
rect 24084 10752 24090 10764
rect 23566 10724 23572 10736
rect 23400 10696 23572 10724
rect 21692 10684 21698 10696
rect 23566 10684 23572 10696
rect 23624 10684 23630 10736
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1636 10628 1685 10656
rect 1636 10616 1642 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 9214 10656 9220 10668
rect 9175 10628 9220 10656
rect 1673 10619 1731 10625
rect 9214 10616 9220 10628
rect 9272 10656 9278 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9272 10628 9873 10656
rect 9272 10616 9278 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 13688 10628 14749 10656
rect 13688 10616 13694 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15160 10628 15853 10656
rect 15160 10616 15166 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 16632 10628 17417 10656
rect 16632 10616 16638 10628
rect 17405 10625 17417 10628
rect 17451 10656 17463 10659
rect 17770 10656 17776 10668
rect 17451 10628 17776 10656
rect 17451 10625 17463 10628
rect 17405 10619 17463 10625
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 21358 10656 21364 10668
rect 21223 10628 21364 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 23860 10665 23888 10752
rect 25038 10724 25044 10736
rect 24999 10696 25044 10724
rect 25038 10684 25044 10696
rect 25096 10684 25102 10736
rect 25498 10684 25504 10736
rect 25556 10684 25562 10736
rect 23845 10659 23903 10665
rect 22296 10628 22494 10656
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 14139 10560 14565 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 15654 10588 15660 10600
rect 15567 10560 15660 10588
rect 14553 10551 14611 10557
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 16022 10548 16028 10600
rect 16080 10588 16086 10600
rect 18138 10588 18144 10600
rect 16080 10560 18144 10588
rect 16080 10548 16086 10560
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10520 9367 10523
rect 15672 10520 15700 10548
rect 9355 10492 15700 10520
rect 9355 10489 9367 10492
rect 9309 10483 9367 10489
rect 16666 10480 16672 10532
rect 16724 10520 16730 10532
rect 17862 10520 17868 10532
rect 16724 10492 17868 10520
rect 16724 10480 16730 10492
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 18248 10520 18276 10551
rect 18322 10548 18328 10600
rect 18380 10588 18386 10600
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18380 10560 18797 10588
rect 18380 10548 18386 10560
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 19426 10588 19432 10600
rect 18785 10551 18843 10557
rect 18892 10560 19432 10588
rect 18892 10520 18920 10560
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 20254 10588 20260 10600
rect 19720 10560 20116 10588
rect 20215 10560 20260 10588
rect 18248 10492 18920 10520
rect 19337 10523 19395 10529
rect 19337 10489 19349 10523
rect 19383 10520 19395 10523
rect 19720 10520 19748 10560
rect 19383 10492 19748 10520
rect 19383 10489 19395 10492
rect 19337 10483 19395 10489
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 15194 10452 15200 10464
rect 15155 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10452 15258 10464
rect 16025 10455 16083 10461
rect 16025 10452 16037 10455
rect 15252 10424 16037 10452
rect 15252 10412 15258 10424
rect 16025 10421 16037 10424
rect 16071 10452 16083 10455
rect 16206 10452 16212 10464
rect 16071 10424 16212 10452
rect 16071 10421 16083 10424
rect 16025 10415 16083 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 17497 10455 17555 10461
rect 17497 10421 17509 10455
rect 17543 10452 17555 10455
rect 19610 10452 19616 10464
rect 17543 10424 19616 10452
rect 17543 10421 17555 10424
rect 17497 10415 17555 10421
rect 19610 10412 19616 10424
rect 19668 10412 19674 10464
rect 20088 10452 20116 10560
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 20438 10548 20444 10600
rect 20496 10588 20502 10600
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 20496 10560 20545 10588
rect 20496 10548 20502 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 22094 10588 22100 10600
rect 20533 10551 20591 10557
rect 20824 10560 22100 10588
rect 20824 10452 20852 10560
rect 22094 10548 22100 10560
rect 22152 10548 22158 10600
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 22296 10520 22324 10628
rect 23845 10625 23857 10659
rect 23891 10656 23903 10659
rect 24765 10659 24823 10665
rect 24765 10656 24777 10659
rect 23891 10628 24777 10656
rect 23891 10625 23903 10628
rect 23845 10619 23903 10625
rect 24765 10625 24777 10628
rect 24811 10625 24823 10659
rect 26436 10656 26464 10764
rect 26513 10761 26525 10795
rect 26559 10792 26571 10795
rect 27614 10792 27620 10804
rect 26559 10764 27620 10792
rect 26559 10761 26571 10764
rect 26513 10755 26571 10761
rect 27614 10752 27620 10764
rect 27672 10792 27678 10804
rect 28442 10792 28448 10804
rect 27672 10764 28448 10792
rect 27672 10752 27678 10764
rect 28442 10752 28448 10764
rect 28500 10752 28506 10804
rect 28718 10752 28724 10804
rect 28776 10792 28782 10804
rect 30926 10792 30932 10804
rect 28776 10764 30932 10792
rect 28776 10752 28782 10764
rect 30926 10752 30932 10764
rect 30984 10792 30990 10804
rect 31113 10795 31171 10801
rect 31113 10792 31125 10795
rect 30984 10764 31125 10792
rect 30984 10752 30990 10764
rect 31113 10761 31125 10764
rect 31159 10761 31171 10795
rect 31662 10792 31668 10804
rect 31623 10764 31668 10792
rect 31113 10755 31171 10761
rect 31662 10752 31668 10764
rect 31720 10792 31726 10804
rect 32861 10795 32919 10801
rect 32861 10792 32873 10795
rect 31720 10764 32873 10792
rect 31720 10752 31726 10764
rect 32861 10761 32873 10764
rect 32907 10761 32919 10795
rect 32861 10755 32919 10761
rect 33410 10752 33416 10804
rect 33468 10792 33474 10804
rect 38105 10795 38163 10801
rect 38105 10792 38117 10795
rect 33468 10764 38117 10792
rect 33468 10752 33474 10764
rect 38105 10761 38117 10764
rect 38151 10761 38163 10795
rect 38105 10755 38163 10761
rect 27430 10684 27436 10736
rect 27488 10724 27494 10736
rect 32401 10727 32459 10733
rect 32401 10724 32413 10727
rect 27488 10696 28566 10724
rect 30116 10696 32413 10724
rect 27488 10684 27494 10696
rect 27341 10659 27399 10665
rect 27341 10656 27353 10659
rect 26436 10628 27353 10656
rect 24765 10619 24823 10625
rect 27341 10625 27353 10628
rect 27387 10625 27399 10659
rect 27341 10619 27399 10625
rect 23198 10548 23204 10600
rect 23256 10588 23262 10600
rect 23256 10560 24072 10588
rect 23256 10548 23262 10560
rect 20956 10492 22324 10520
rect 20956 10480 20962 10492
rect 20088 10424 20852 10452
rect 22097 10455 22155 10461
rect 22097 10421 22109 10455
rect 22143 10452 22155 10455
rect 22462 10452 22468 10464
rect 22143 10424 22468 10452
rect 22143 10421 22155 10424
rect 22097 10415 22155 10421
rect 22462 10412 22468 10424
rect 22520 10452 22526 10464
rect 22830 10452 22836 10464
rect 22520 10424 22836 10452
rect 22520 10412 22526 10424
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 24044 10452 24072 10560
rect 24210 10548 24216 10600
rect 24268 10588 24274 10600
rect 27246 10588 27252 10600
rect 24268 10560 27252 10588
rect 24268 10548 24274 10560
rect 27246 10548 27252 10560
rect 27304 10548 27310 10600
rect 27249 10455 27307 10461
rect 27249 10452 27261 10455
rect 24044 10424 27261 10452
rect 27249 10421 27261 10424
rect 27295 10421 27307 10455
rect 27356 10452 27384 10619
rect 27985 10591 28043 10597
rect 27985 10557 27997 10591
rect 28031 10588 28043 10591
rect 28534 10588 28540 10600
rect 28031 10560 28540 10588
rect 28031 10557 28043 10560
rect 27985 10551 28043 10557
rect 28534 10548 28540 10560
rect 28592 10548 28598 10600
rect 29362 10548 29368 10600
rect 29420 10588 29426 10600
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29420 10560 29745 10588
rect 29420 10548 29426 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 30006 10588 30012 10600
rect 29967 10560 30012 10588
rect 29733 10551 29791 10557
rect 30006 10548 30012 10560
rect 30064 10548 30070 10600
rect 30116 10452 30144 10696
rect 32401 10693 32413 10696
rect 32447 10724 32459 10727
rect 33134 10724 33140 10736
rect 32447 10696 33140 10724
rect 32447 10693 32459 10696
rect 32401 10687 32459 10693
rect 33134 10684 33140 10696
rect 33192 10684 33198 10736
rect 30653 10659 30711 10665
rect 30653 10625 30665 10659
rect 30699 10656 30711 10659
rect 33428 10656 33456 10752
rect 30699 10628 33456 10656
rect 37645 10659 37703 10665
rect 30699 10625 30711 10628
rect 30653 10619 30711 10625
rect 37645 10625 37657 10659
rect 37691 10656 37703 10659
rect 38286 10656 38292 10668
rect 37691 10628 38292 10656
rect 37691 10625 37703 10628
rect 37645 10619 37703 10625
rect 38286 10616 38292 10628
rect 38344 10616 38350 10668
rect 27356 10424 30144 10452
rect 27249 10415 27307 10421
rect 30190 10412 30196 10464
rect 30248 10452 30254 10464
rect 30561 10455 30619 10461
rect 30561 10452 30573 10455
rect 30248 10424 30573 10452
rect 30248 10412 30254 10424
rect 30561 10421 30573 10424
rect 30607 10421 30619 10455
rect 30561 10415 30619 10421
rect 30926 10412 30932 10464
rect 30984 10452 30990 10464
rect 32030 10452 32036 10464
rect 30984 10424 32036 10452
rect 30984 10412 30990 10424
rect 32030 10412 32036 10424
rect 32088 10412 32094 10464
rect 33134 10412 33140 10464
rect 33192 10452 33198 10464
rect 33413 10455 33471 10461
rect 33413 10452 33425 10455
rect 33192 10424 33425 10452
rect 33192 10412 33198 10424
rect 33413 10421 33425 10424
rect 33459 10421 33471 10455
rect 33413 10415 33471 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 10962 10248 10968 10260
rect 1820 10220 6914 10248
rect 10923 10220 10968 10248
rect 1820 10208 1826 10220
rect 6886 10180 6914 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 15562 10248 15568 10260
rect 12584 10220 15568 10248
rect 12584 10208 12590 10220
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 20622 10248 20628 10260
rect 16132 10220 20628 10248
rect 13354 10180 13360 10192
rect 6886 10152 13360 10180
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10112 13231 10115
rect 13219 10084 14872 10112
rect 13219 10081 13231 10084
rect 13173 10075 13231 10081
rect 14844 10056 14872 10084
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15436 10084 15481 10112
rect 15436 10072 15442 10084
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 14550 10044 14556 10056
rect 11103 10016 14556 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 14734 10044 14740 10056
rect 14691 10016 14740 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 14884 10016 15301 10044
rect 14884 10004 14890 10016
rect 15289 10013 15301 10016
rect 15335 10044 15347 10047
rect 15470 10044 15476 10056
rect 15335 10016 15476 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 16132 10053 16160 10220
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 20806 10248 20812 10260
rect 20767 10220 20812 10248
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 23658 10208 23664 10260
rect 23716 10248 23722 10260
rect 25409 10251 25467 10257
rect 25409 10248 25421 10251
rect 23716 10220 25421 10248
rect 23716 10208 23722 10220
rect 25409 10217 25421 10220
rect 25455 10217 25467 10251
rect 26786 10248 26792 10260
rect 25409 10211 25467 10217
rect 25884 10220 26792 10248
rect 17218 10180 17224 10192
rect 17179 10152 17224 10180
rect 17218 10140 17224 10152
rect 17276 10140 17282 10192
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 19521 10183 19579 10189
rect 19521 10180 19533 10183
rect 17828 10152 19533 10180
rect 17828 10140 17834 10152
rect 19521 10149 19533 10152
rect 19567 10149 19579 10183
rect 19521 10143 19579 10149
rect 19610 10140 19616 10192
rect 19668 10180 19674 10192
rect 20438 10180 20444 10192
rect 19668 10152 20444 10180
rect 19668 10140 19674 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 25498 10180 25504 10192
rect 23308 10152 25504 10180
rect 18506 10112 18512 10124
rect 18467 10084 18512 10112
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 23308 10112 23336 10152
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 18616 10084 23336 10112
rect 23385 10115 23443 10121
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 13725 9979 13783 9985
rect 13725 9945 13737 9979
rect 13771 9976 13783 9979
rect 16666 9976 16672 9988
rect 13771 9948 16672 9976
rect 13771 9945 13783 9948
rect 13725 9939 13783 9945
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 16758 9936 16764 9988
rect 16816 9976 16822 9988
rect 17862 9976 17868 9988
rect 16816 9948 16861 9976
rect 17823 9948 17868 9976
rect 16816 9936 16822 9948
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 17954 9936 17960 9988
rect 18012 9976 18018 9988
rect 18012 9948 18057 9976
rect 18012 9936 18018 9948
rect 18138 9936 18144 9988
rect 18196 9976 18202 9988
rect 18616 9976 18644 10084
rect 23385 10081 23397 10115
rect 23431 10112 23443 10115
rect 23842 10112 23848 10124
rect 23431 10084 23848 10112
rect 23431 10081 23443 10084
rect 23385 10075 23443 10081
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 24029 10115 24087 10121
rect 24029 10081 24041 10115
rect 24075 10112 24087 10115
rect 24486 10112 24492 10124
rect 24075 10084 24492 10112
rect 24075 10081 24087 10084
rect 24029 10075 24087 10081
rect 24486 10072 24492 10084
rect 24544 10072 24550 10124
rect 25884 10112 25912 10220
rect 26786 10208 26792 10220
rect 26844 10208 26850 10260
rect 26899 10251 26957 10257
rect 26899 10217 26911 10251
rect 26945 10248 26957 10251
rect 27614 10248 27620 10260
rect 26945 10220 27620 10248
rect 26945 10217 26957 10220
rect 26899 10211 26957 10217
rect 27614 10208 27620 10220
rect 27672 10208 27678 10260
rect 27982 10208 27988 10260
rect 28040 10248 28046 10260
rect 28718 10248 28724 10260
rect 28040 10220 28724 10248
rect 28040 10208 28046 10220
rect 28718 10208 28724 10220
rect 28776 10208 28782 10260
rect 28902 10248 28908 10260
rect 28863 10220 28908 10248
rect 28902 10208 28908 10220
rect 28960 10208 28966 10260
rect 30282 10208 30288 10260
rect 30340 10248 30346 10260
rect 31309 10251 31367 10257
rect 31309 10248 31321 10251
rect 30340 10220 31321 10248
rect 30340 10208 30346 10220
rect 31309 10217 31321 10220
rect 31355 10248 31367 10251
rect 32030 10248 32036 10260
rect 31355 10220 31754 10248
rect 31991 10220 32036 10248
rect 31355 10217 31367 10220
rect 31309 10211 31367 10217
rect 27246 10140 27252 10192
rect 27304 10180 27310 10192
rect 30190 10180 30196 10192
rect 27304 10152 30196 10180
rect 27304 10140 27310 10152
rect 24780 10084 25912 10112
rect 20898 10044 20904 10056
rect 20859 10016 20904 10044
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 22002 10004 22008 10056
rect 22060 10004 22066 10056
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 24780 10053 24808 10084
rect 26234 10072 26240 10124
rect 26292 10112 26298 10124
rect 27154 10112 27160 10124
rect 26292 10084 27160 10112
rect 26292 10072 26298 10084
rect 27154 10072 27160 10084
rect 27212 10072 27218 10124
rect 27985 10115 28043 10121
rect 27985 10081 27997 10115
rect 28031 10112 28043 10115
rect 28074 10112 28080 10124
rect 28031 10084 28080 10112
rect 28031 10081 28043 10084
rect 27985 10075 28043 10081
rect 28074 10072 28080 10084
rect 28132 10072 28138 10124
rect 28276 10121 28304 10152
rect 30190 10140 30196 10152
rect 30248 10140 30254 10192
rect 31726 10180 31754 10220
rect 32030 10208 32036 10220
rect 32088 10208 32094 10260
rect 32306 10180 32312 10192
rect 31726 10152 32312 10180
rect 32306 10140 32312 10152
rect 32364 10180 32370 10192
rect 33689 10183 33747 10189
rect 33689 10180 33701 10183
rect 32364 10152 33701 10180
rect 32364 10140 32370 10152
rect 33689 10149 33701 10152
rect 33735 10149 33747 10183
rect 33689 10143 33747 10149
rect 28261 10115 28319 10121
rect 28261 10081 28273 10115
rect 28307 10081 28319 10115
rect 28261 10075 28319 10081
rect 30006 10072 30012 10124
rect 30064 10112 30070 10124
rect 31573 10115 31631 10121
rect 31573 10112 31585 10115
rect 30064 10084 31585 10112
rect 30064 10072 30070 10084
rect 31573 10081 31585 10084
rect 31619 10112 31631 10115
rect 31619 10084 32720 10112
rect 31619 10081 31631 10084
rect 31573 10075 31631 10081
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 23624 10016 24777 10044
rect 23624 10004 23630 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10044 29055 10047
rect 29638 10044 29644 10056
rect 29043 10016 29644 10044
rect 29043 10013 29055 10016
rect 28997 10007 29055 10013
rect 29638 10004 29644 10016
rect 29696 10004 29702 10056
rect 18196 9948 18644 9976
rect 18196 9936 18202 9948
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19610 9976 19616 9988
rect 19392 9948 19616 9976
rect 19392 9936 19398 9948
rect 19610 9936 19616 9948
rect 19668 9936 19674 9988
rect 19978 9976 19984 9988
rect 19939 9948 19984 9976
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 20073 9979 20131 9985
rect 20073 9945 20085 9979
rect 20119 9976 20131 9979
rect 20530 9976 20536 9988
rect 20119 9948 20536 9976
rect 20119 9945 20131 9948
rect 20073 9939 20131 9945
rect 20530 9936 20536 9948
rect 20588 9936 20594 9988
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 21266 9976 21272 9988
rect 20772 9948 21272 9976
rect 20772 9936 20778 9948
rect 21266 9936 21272 9948
rect 21324 9976 21330 9988
rect 21361 9979 21419 9985
rect 21361 9976 21373 9979
rect 21324 9948 21373 9976
rect 21324 9936 21330 9948
rect 21361 9945 21373 9948
rect 21407 9945 21419 9979
rect 21361 9939 21419 9945
rect 23109 9979 23167 9985
rect 23109 9945 23121 9979
rect 23155 9976 23167 9979
rect 23750 9976 23756 9988
rect 23155 9948 23756 9976
rect 23155 9945 23167 9948
rect 23109 9939 23167 9945
rect 23750 9936 23756 9948
rect 23808 9936 23814 9988
rect 24854 9936 24860 9988
rect 24912 9976 24918 9988
rect 24912 9948 25714 9976
rect 24912 9936 24918 9948
rect 26786 9936 26792 9988
rect 26844 9976 26850 9988
rect 27982 9976 27988 9988
rect 26844 9948 27988 9976
rect 26844 9936 26850 9948
rect 27982 9936 27988 9948
rect 28040 9936 28046 9988
rect 32692 9985 32720 10084
rect 33134 10072 33140 10124
rect 33192 10072 33198 10124
rect 33152 10044 33180 10072
rect 35345 10047 35403 10053
rect 35345 10044 35357 10047
rect 33152 10016 35357 10044
rect 35345 10013 35357 10016
rect 35391 10044 35403 10047
rect 35805 10047 35863 10053
rect 35805 10044 35817 10047
rect 35391 10016 35817 10044
rect 35391 10013 35403 10016
rect 35345 10007 35403 10013
rect 35805 10013 35817 10016
rect 35851 10013 35863 10047
rect 35805 10007 35863 10013
rect 28169 9979 28227 9985
rect 28169 9945 28181 9979
rect 28215 9945 28227 9979
rect 32677 9979 32735 9985
rect 28169 9939 28227 9945
rect 28368 9948 29960 9976
rect 30866 9948 30972 9976
rect 14737 9911 14795 9917
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 15746 9908 15752 9920
rect 14783 9880 15752 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 18322 9908 18328 9920
rect 16071 9880 18328 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 18598 9868 18604 9920
rect 18656 9908 18662 9920
rect 24026 9908 24032 9920
rect 18656 9880 24032 9908
rect 18656 9868 18662 9880
rect 24026 9868 24032 9880
rect 24084 9868 24090 9920
rect 24118 9868 24124 9920
rect 24176 9908 24182 9920
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 24176 9880 24685 9908
rect 24176 9868 24182 9880
rect 24673 9877 24685 9880
rect 24719 9877 24731 9911
rect 24673 9871 24731 9877
rect 24762 9868 24768 9920
rect 24820 9908 24826 9920
rect 28074 9908 28080 9920
rect 24820 9880 28080 9908
rect 24820 9868 24826 9880
rect 28074 9868 28080 9880
rect 28132 9868 28138 9920
rect 28184 9908 28212 9939
rect 28368 9908 28396 9948
rect 28184 9880 28396 9908
rect 28442 9868 28448 9920
rect 28500 9908 28506 9920
rect 29546 9908 29552 9920
rect 28500 9880 29552 9908
rect 28500 9868 28506 9880
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 29730 9868 29736 9920
rect 29788 9908 29794 9920
rect 29825 9911 29883 9917
rect 29825 9908 29837 9911
rect 29788 9880 29837 9908
rect 29788 9868 29794 9880
rect 29825 9877 29837 9880
rect 29871 9877 29883 9911
rect 29932 9908 29960 9948
rect 30466 9908 30472 9920
rect 29932 9880 30472 9908
rect 29825 9871 29883 9877
rect 30466 9868 30472 9880
rect 30524 9868 30530 9920
rect 30944 9908 30972 9948
rect 32677 9945 32689 9979
rect 32723 9976 32735 9979
rect 33137 9979 33195 9985
rect 33137 9976 33149 9979
rect 32723 9948 33149 9976
rect 32723 9945 32735 9948
rect 32677 9939 32735 9945
rect 33137 9945 33149 9948
rect 33183 9945 33195 9979
rect 35253 9979 35311 9985
rect 35253 9976 35265 9979
rect 33137 9939 33195 9945
rect 33244 9948 35265 9976
rect 33244 9908 33272 9948
rect 35253 9945 35265 9948
rect 35299 9945 35311 9979
rect 35253 9939 35311 9945
rect 30944 9880 33272 9908
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 9214 9704 9220 9716
rect 6880 9676 9220 9704
rect 6880 9664 6886 9676
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 14734 9704 14740 9716
rect 14292 9676 14740 9704
rect 9401 9639 9459 9645
rect 9401 9605 9413 9639
rect 9447 9636 9459 9639
rect 11974 9636 11980 9648
rect 9447 9608 11980 9636
rect 9447 9605 9459 9608
rect 9401 9599 9459 9605
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 9416 9568 9444 9599
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 13173 9639 13231 9645
rect 13173 9605 13185 9639
rect 13219 9636 13231 9639
rect 14292 9636 14320 9676
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 15013 9707 15071 9713
rect 15013 9673 15025 9707
rect 15059 9704 15071 9707
rect 20806 9704 20812 9716
rect 15059 9676 20812 9704
rect 15059 9673 15071 9676
rect 15013 9667 15071 9673
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 22462 9704 22468 9716
rect 20956 9676 22468 9704
rect 20956 9664 20962 9676
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 24762 9704 24768 9716
rect 22664 9676 24768 9704
rect 13219 9608 14320 9636
rect 14369 9639 14427 9645
rect 13219 9605 13231 9608
rect 13173 9599 13231 9605
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 14415 9608 15761 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 15749 9605 15761 9608
rect 15795 9605 15807 9639
rect 15749 9599 15807 9605
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 15896 9608 17141 9636
rect 15896 9596 15902 9608
rect 17129 9605 17141 9608
rect 17175 9605 17187 9639
rect 17678 9636 17684 9648
rect 17639 9608 17684 9636
rect 17129 9599 17187 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18322 9636 18328 9648
rect 18283 9608 18328 9636
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 18874 9596 18880 9648
rect 18932 9636 18938 9648
rect 22097 9639 22155 9645
rect 18932 9608 20470 9636
rect 18932 9596 18938 9608
rect 22097 9605 22109 9639
rect 22143 9636 22155 9639
rect 22278 9636 22284 9648
rect 22143 9608 22284 9636
rect 22143 9605 22155 9608
rect 22097 9599 22155 9605
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 22664 9645 22692 9676
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 25682 9664 25688 9716
rect 25740 9704 25746 9716
rect 34790 9704 34796 9716
rect 25740 9676 34796 9704
rect 25740 9664 25746 9676
rect 34790 9664 34796 9676
rect 34848 9664 34854 9716
rect 22649 9639 22707 9645
rect 22649 9636 22661 9639
rect 22428 9608 22661 9636
rect 22428 9596 22434 9608
rect 22649 9605 22661 9608
rect 22695 9605 22707 9639
rect 22649 9599 22707 9605
rect 23201 9639 23259 9645
rect 23201 9605 23213 9639
rect 23247 9636 23259 9639
rect 24118 9636 24124 9648
rect 23247 9608 24124 9636
rect 23247 9605 23259 9608
rect 23201 9599 23259 9605
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 25590 9636 25596 9648
rect 25162 9608 25596 9636
rect 25590 9596 25596 9608
rect 25648 9596 25654 9648
rect 25958 9596 25964 9648
rect 26016 9636 26022 9648
rect 26421 9639 26479 9645
rect 26421 9636 26433 9639
rect 26016 9608 26433 9636
rect 26016 9596 26022 9608
rect 26421 9605 26433 9608
rect 26467 9605 26479 9639
rect 26421 9599 26479 9605
rect 27249 9639 27307 9645
rect 27249 9605 27261 9639
rect 27295 9636 27307 9639
rect 27522 9636 27528 9648
rect 27295 9608 27528 9636
rect 27295 9605 27307 9608
rect 27249 9599 27307 9605
rect 27522 9596 27528 9608
rect 27580 9596 27586 9648
rect 27614 9596 27620 9648
rect 27672 9636 27678 9648
rect 29638 9636 29644 9648
rect 27672 9608 28474 9636
rect 29551 9608 29644 9636
rect 27672 9596 27678 9608
rect 29638 9596 29644 9608
rect 29696 9636 29702 9648
rect 30006 9636 30012 9648
rect 29696 9608 30012 9636
rect 29696 9596 29702 9608
rect 30006 9596 30012 9608
rect 30064 9596 30070 9648
rect 30469 9639 30527 9645
rect 30469 9605 30481 9639
rect 30515 9636 30527 9639
rect 30558 9636 30564 9648
rect 30515 9608 30564 9636
rect 30515 9605 30527 9608
rect 30469 9599 30527 9605
rect 30558 9596 30564 9608
rect 30616 9596 30622 9648
rect 30650 9596 30656 9648
rect 30708 9636 30714 9648
rect 32766 9636 32772 9648
rect 30708 9608 32772 9636
rect 30708 9596 30714 9608
rect 32766 9596 32772 9608
rect 32824 9596 32830 9648
rect 8895 9540 9444 9568
rect 12621 9571 12679 9577
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 12621 9537 12633 9571
rect 12667 9568 12679 9571
rect 13630 9568 13636 9580
rect 12667 9540 13636 9568
rect 12667 9537 12679 9540
rect 12621 9531 12679 9537
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13964 9540 14289 9568
rect 13964 9528 13970 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14936 9432 14964 9531
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21784 9540 22017 9568
rect 21784 9528 21790 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 25869 9571 25927 9577
rect 25869 9537 25881 9571
rect 25915 9568 25927 9571
rect 26234 9568 26240 9580
rect 25915 9540 26240 9568
rect 25915 9537 25927 9540
rect 25869 9531 25927 9537
rect 26234 9528 26240 9540
rect 26292 9528 26298 9580
rect 26513 9571 26571 9577
rect 26513 9537 26525 9571
rect 26559 9568 26571 9571
rect 27157 9571 27215 9577
rect 26559 9540 26832 9568
rect 26559 9537 26571 9540
rect 26513 9531 26571 9537
rect 15654 9500 15660 9512
rect 15615 9472 15660 9500
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15930 9500 15936 9512
rect 15891 9472 15936 9500
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 17037 9503 17095 9509
rect 17037 9469 17049 9503
rect 17083 9500 17095 9503
rect 17126 9500 17132 9512
rect 17083 9472 17132 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 17920 9472 18245 9500
rect 17920 9460 17926 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 21453 9503 21511 9509
rect 20027 9472 21036 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 17954 9432 17960 9444
rect 14056 9404 17960 9432
rect 14056 9392 14062 9404
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 18782 9432 18788 9444
rect 18743 9404 18788 9432
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 8662 9364 8668 9376
rect 8623 9336 8668 9364
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 13722 9364 13728 9376
rect 13683 9336 13728 9364
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 17126 9324 17132 9376
rect 17184 9364 17190 9376
rect 18230 9364 18236 9376
rect 17184 9336 18236 9364
rect 17184 9324 17190 9336
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 19720 9364 19748 9463
rect 21008 9432 21036 9472
rect 21453 9469 21465 9503
rect 21499 9500 21511 9503
rect 21499 9472 23152 9500
rect 21499 9469 21511 9472
rect 21453 9463 21511 9469
rect 22554 9432 22560 9444
rect 21008 9404 22560 9432
rect 22554 9392 22560 9404
rect 22612 9392 22618 9444
rect 21358 9364 21364 9376
rect 19720 9336 21364 9364
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 23124 9364 23152 9472
rect 23198 9460 23204 9512
rect 23256 9500 23262 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 23256 9472 23305 9500
rect 23256 9460 23262 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 23566 9460 23572 9512
rect 23624 9500 23630 9512
rect 23845 9503 23903 9509
rect 23845 9500 23857 9503
rect 23624 9472 23857 9500
rect 23624 9460 23630 9472
rect 23845 9469 23857 9472
rect 23891 9500 23903 9503
rect 23934 9500 23940 9512
rect 23891 9472 23940 9500
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 23934 9460 23940 9472
rect 23992 9460 23998 9512
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 26694 9500 26700 9512
rect 25639 9472 26700 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 26694 9460 26700 9472
rect 26752 9460 26758 9512
rect 26804 9364 26832 9540
rect 27157 9537 27169 9571
rect 27203 9568 27215 9571
rect 27706 9568 27712 9580
rect 27203 9540 27712 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 27706 9528 27712 9540
rect 27764 9528 27770 9580
rect 32398 9568 32404 9580
rect 32359 9540 32404 9568
rect 32398 9528 32404 9540
rect 32456 9528 32462 9580
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9537 32551 9571
rect 33134 9568 33140 9580
rect 33095 9540 33140 9568
rect 32493 9531 32551 9537
rect 27338 9460 27344 9512
rect 27396 9500 27402 9512
rect 27893 9503 27951 9509
rect 27893 9500 27905 9503
rect 27396 9472 27905 9500
rect 27396 9460 27402 9472
rect 27893 9469 27905 9472
rect 27939 9469 27951 9503
rect 27893 9463 27951 9469
rect 28074 9460 28080 9512
rect 28132 9500 28138 9512
rect 28132 9472 29868 9500
rect 28132 9460 28138 9472
rect 29840 9432 29868 9472
rect 29914 9460 29920 9512
rect 29972 9500 29978 9512
rect 29972 9472 30017 9500
rect 29972 9460 29978 9472
rect 32508 9432 32536 9531
rect 33134 9528 33140 9540
rect 33192 9528 33198 9580
rect 34149 9435 34207 9441
rect 34149 9432 34161 9435
rect 29840 9404 34161 9432
rect 34149 9401 34161 9404
rect 34195 9432 34207 9435
rect 36078 9432 36084 9444
rect 34195 9404 36084 9432
rect 34195 9401 34207 9404
rect 34149 9395 34207 9401
rect 36078 9392 36084 9404
rect 36136 9392 36142 9444
rect 29086 9364 29092 9376
rect 23124 9336 29092 9364
rect 29086 9324 29092 9336
rect 29144 9324 29150 9376
rect 29178 9324 29184 9376
rect 29236 9364 29242 9376
rect 30650 9364 30656 9376
rect 29236 9336 30656 9364
rect 29236 9324 29242 9336
rect 30650 9324 30656 9336
rect 30708 9324 30714 9376
rect 30926 9364 30932 9376
rect 30887 9336 30932 9364
rect 30926 9324 30932 9336
rect 30984 9364 30990 9376
rect 31481 9367 31539 9373
rect 31481 9364 31493 9367
rect 30984 9336 31493 9364
rect 30984 9324 30990 9336
rect 31481 9333 31493 9336
rect 31527 9333 31539 9367
rect 33042 9364 33048 9376
rect 33003 9336 33048 9364
rect 31481 9327 31539 9333
rect 33042 9324 33048 9336
rect 33100 9324 33106 9376
rect 33594 9364 33600 9376
rect 33555 9336 33600 9364
rect 33594 9324 33600 9336
rect 33652 9324 33658 9376
rect 37550 9364 37556 9376
rect 37511 9336 37556 9364
rect 37550 9324 37556 9336
rect 37608 9324 37614 9376
rect 38286 9364 38292 9376
rect 38247 9336 38292 9364
rect 38286 9324 38292 9336
rect 38344 9324 38350 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 20622 9160 20628 9172
rect 13780 9132 20628 9160
rect 13780 9120 13786 9132
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 22094 9160 22100 9172
rect 21560 9132 22100 9160
rect 14829 9095 14887 9101
rect 14829 9061 14841 9095
rect 14875 9092 14887 9095
rect 17862 9092 17868 9104
rect 14875 9064 17868 9092
rect 14875 9061 14887 9064
rect 14829 9055 14887 9061
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 17954 9052 17960 9104
rect 18012 9092 18018 9104
rect 19702 9092 19708 9104
rect 18012 9064 19708 9092
rect 18012 9052 18018 9064
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 19978 9052 19984 9104
rect 20036 9092 20042 9104
rect 20717 9095 20775 9101
rect 20717 9092 20729 9095
rect 20036 9064 20729 9092
rect 20036 9052 20042 9064
rect 20717 9061 20729 9064
rect 20763 9061 20775 9095
rect 20717 9055 20775 9061
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 21560 9092 21588 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 22704 9132 23673 9160
rect 22704 9120 22710 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 26602 9160 26608 9172
rect 23661 9123 23719 9129
rect 25148 9132 26608 9160
rect 21048 9064 21588 9092
rect 21048 9052 21054 9064
rect 23198 9052 23204 9104
rect 23256 9092 23262 9104
rect 25148 9092 25176 9132
rect 26602 9120 26608 9132
rect 26660 9120 26666 9172
rect 26694 9120 26700 9172
rect 26752 9160 26758 9172
rect 26973 9163 27031 9169
rect 26973 9160 26985 9163
rect 26752 9132 26985 9160
rect 26752 9120 26758 9132
rect 26973 9129 26985 9132
rect 27019 9129 27031 9163
rect 26973 9123 27031 9129
rect 27356 9132 29316 9160
rect 27356 9104 27384 9132
rect 27338 9092 27344 9104
rect 23256 9064 25176 9092
rect 26344 9064 27344 9092
rect 23256 9052 23262 9064
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 4062 9024 4068 9036
rect 1903 8996 4068 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 15930 9024 15936 9036
rect 15519 8996 15936 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 9024 16175 9027
rect 17126 9024 17132 9036
rect 16163 8996 17132 9024
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 18690 9024 18696 9036
rect 18651 8996 18696 9024
rect 18690 8984 18696 8996
rect 18748 9024 18754 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 18748 8996 19809 9024
rect 18748 8984 18754 8996
rect 19797 8993 19809 8996
rect 19843 9024 19855 9027
rect 21174 9024 21180 9036
rect 19843 8996 21180 9024
rect 19843 8993 19855 8996
rect 19797 8987 19855 8993
rect 21174 8984 21180 8996
rect 21232 8984 21238 9036
rect 21358 8984 21364 9036
rect 21416 9024 21422 9036
rect 23109 9027 23167 9033
rect 23109 9024 23121 9027
rect 21416 8996 23121 9024
rect 21416 8984 21422 8996
rect 23109 8993 23121 8996
rect 23155 9024 23167 9027
rect 23474 9024 23480 9036
rect 23155 8996 23480 9024
rect 23155 8993 23167 8996
rect 23109 8987 23167 8993
rect 23474 8984 23480 8996
rect 23532 8984 23538 9036
rect 24026 8984 24032 9036
rect 24084 9024 24090 9036
rect 26145 9027 26203 9033
rect 26145 9024 26157 9027
rect 24084 8996 26157 9024
rect 24084 8984 24090 8996
rect 26145 8993 26157 8996
rect 26191 9024 26203 9027
rect 26344 9024 26372 9064
rect 27338 9052 27344 9064
rect 27396 9052 27402 9104
rect 29288 9092 29316 9132
rect 29362 9120 29368 9172
rect 29420 9160 29426 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 29420 9132 29837 9160
rect 29420 9120 29426 9132
rect 29825 9129 29837 9132
rect 29871 9129 29883 9163
rect 32033 9163 32091 9169
rect 32033 9160 32045 9163
rect 29825 9123 29883 9129
rect 29932 9132 32045 9160
rect 29932 9092 29960 9132
rect 32033 9129 32045 9132
rect 32079 9129 32091 9163
rect 32033 9123 32091 9129
rect 29288 9064 29960 9092
rect 30024 9064 30236 9092
rect 28721 9027 28779 9033
rect 28721 9024 28733 9027
rect 26191 8996 26372 9024
rect 26436 8996 28733 9024
rect 26191 8993 26203 8996
rect 26145 8987 26203 8993
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 12492 8928 12725 8956
rect 12492 8916 12498 8928
rect 12713 8925 12725 8928
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 15286 8956 15292 8968
rect 14783 8928 15292 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8956 20867 8959
rect 23753 8959 23811 8965
rect 20855 8928 21128 8956
rect 20855 8925 20867 8928
rect 20809 8919 20867 8925
rect 12805 8891 12863 8897
rect 12805 8857 12817 8891
rect 12851 8857 12863 8891
rect 12805 8851 12863 8857
rect 13725 8891 13783 8897
rect 13725 8857 13737 8891
rect 13771 8888 13783 8891
rect 13998 8888 14004 8900
rect 13771 8860 14004 8888
rect 13771 8857 13783 8860
rect 13725 8851 13783 8857
rect 12820 8820 12848 8851
rect 13998 8848 14004 8860
rect 14056 8848 14062 8900
rect 15562 8888 15568 8900
rect 15523 8860 15568 8888
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 16482 8888 16488 8900
rect 15672 8860 16488 8888
rect 15672 8820 15700 8860
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 16670 8891 16728 8897
rect 16670 8888 16682 8891
rect 16592 8860 16682 8888
rect 16592 8832 16620 8860
rect 16670 8857 16682 8860
rect 16716 8857 16728 8891
rect 16670 8851 16728 8857
rect 16761 8891 16819 8897
rect 16761 8857 16773 8891
rect 16807 8888 16819 8891
rect 16850 8888 16856 8900
rect 16807 8860 16856 8888
rect 16807 8857 16819 8860
rect 16761 8851 16819 8857
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 18230 8888 18236 8900
rect 18191 8860 18236 8888
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 18322 8848 18328 8900
rect 18380 8888 18386 8900
rect 18380 8860 18425 8888
rect 18380 8848 18386 8860
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 19521 8891 19579 8897
rect 19521 8888 19533 8891
rect 19392 8860 19533 8888
rect 19392 8848 19398 8860
rect 19521 8857 19533 8860
rect 19567 8857 19579 8891
rect 19521 8851 19579 8857
rect 19613 8891 19671 8897
rect 19613 8857 19625 8891
rect 19659 8857 19671 8891
rect 19613 8851 19671 8857
rect 12820 8792 15700 8820
rect 16574 8780 16580 8832
rect 16632 8780 16638 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 19628 8820 19656 8851
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 20990 8888 20996 8900
rect 19760 8860 20996 8888
rect 19760 8848 19766 8860
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 21100 8888 21128 8928
rect 23753 8925 23765 8959
rect 23799 8956 23811 8959
rect 24302 8956 24308 8968
rect 23799 8928 24308 8956
rect 23799 8925 23811 8928
rect 23753 8919 23811 8925
rect 24302 8916 24308 8928
rect 24360 8916 24366 8968
rect 26436 8965 26464 8996
rect 28721 8993 28733 8996
rect 28767 9024 28779 9027
rect 29914 9024 29920 9036
rect 28767 8996 29920 9024
rect 28767 8993 28779 8996
rect 28721 8987 28779 8993
rect 29914 8984 29920 8996
rect 29972 9024 29978 9036
rect 30024 9024 30052 9064
rect 29972 8996 30052 9024
rect 30208 9024 30236 9064
rect 32766 9052 32772 9104
rect 32824 9092 32830 9104
rect 33137 9095 33195 9101
rect 33137 9092 33149 9095
rect 32824 9064 33149 9092
rect 32824 9052 32830 9064
rect 33137 9061 33149 9064
rect 33183 9061 33195 9095
rect 33137 9055 33195 9061
rect 30926 9024 30932 9036
rect 30208 8996 30932 9024
rect 29972 8984 29978 8996
rect 30926 8984 30932 8996
rect 30984 9024 30990 9036
rect 31570 9024 31576 9036
rect 30984 8996 31576 9024
rect 30984 8984 30990 8996
rect 31570 8984 31576 8996
rect 31628 8984 31634 9036
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8925 26479 8959
rect 36078 8956 36084 8968
rect 36039 8928 36084 8956
rect 26421 8919 26479 8925
rect 21100 8860 21496 8888
rect 17368 8792 19656 8820
rect 17368 8780 17374 8792
rect 21082 8780 21088 8832
rect 21140 8820 21146 8832
rect 21361 8823 21419 8829
rect 21361 8820 21373 8823
rect 21140 8792 21373 8820
rect 21140 8780 21146 8792
rect 21361 8789 21373 8792
rect 21407 8789 21419 8823
rect 21468 8820 21496 8860
rect 21542 8848 21548 8900
rect 21600 8888 21606 8900
rect 21600 8860 21666 8888
rect 21600 8848 21606 8860
rect 22554 8848 22560 8900
rect 22612 8888 22618 8900
rect 22833 8891 22891 8897
rect 22833 8888 22845 8891
rect 22612 8860 22845 8888
rect 22612 8848 22618 8860
rect 22833 8857 22845 8860
rect 22879 8888 22891 8891
rect 22879 8860 24716 8888
rect 22879 8857 22891 8860
rect 22833 8851 22891 8857
rect 22922 8820 22928 8832
rect 21468 8792 22928 8820
rect 21361 8783 21419 8789
rect 22922 8780 22928 8792
rect 22980 8780 22986 8832
rect 23198 8780 23204 8832
rect 23256 8820 23262 8832
rect 24578 8820 24584 8832
rect 23256 8792 24584 8820
rect 23256 8780 23262 8792
rect 24578 8780 24584 8792
rect 24636 8780 24642 8832
rect 24688 8829 24716 8860
rect 24854 8848 24860 8900
rect 24912 8888 24918 8900
rect 24912 8860 24978 8888
rect 24912 8848 24918 8860
rect 26234 8848 26240 8900
rect 26292 8888 26298 8900
rect 26436 8888 26464 8919
rect 36078 8916 36084 8928
rect 36136 8956 36142 8968
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 36136 8928 36553 8956
rect 36136 8916 36142 8928
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 37550 8956 37556 8968
rect 37511 8928 37556 8956
rect 36541 8919 36599 8925
rect 37550 8916 37556 8928
rect 37608 8956 37614 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 37608 8928 38025 8956
rect 37608 8916 37614 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 26292 8860 26464 8888
rect 26528 8860 27278 8888
rect 26292 8848 26298 8860
rect 24673 8823 24731 8829
rect 24673 8789 24685 8823
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 25498 8780 25504 8832
rect 25556 8820 25562 8832
rect 26528 8820 26556 8860
rect 28350 8848 28356 8900
rect 28408 8888 28414 8900
rect 28445 8891 28503 8897
rect 28445 8888 28457 8891
rect 28408 8860 28457 8888
rect 28408 8848 28414 8860
rect 28445 8857 28457 8860
rect 28491 8888 28503 8891
rect 29178 8888 29184 8900
rect 28491 8860 29184 8888
rect 28491 8857 28503 8860
rect 28445 8851 28503 8857
rect 29178 8848 29184 8860
rect 29236 8888 29242 8900
rect 29638 8888 29644 8900
rect 29236 8860 29644 8888
rect 29236 8848 29242 8860
rect 29638 8848 29644 8860
rect 29696 8848 29702 8900
rect 30558 8848 30564 8900
rect 30616 8848 30622 8900
rect 31294 8888 31300 8900
rect 31207 8860 31300 8888
rect 31294 8848 31300 8860
rect 31352 8848 31358 8900
rect 32582 8888 32588 8900
rect 32543 8860 32588 8888
rect 32582 8848 32588 8860
rect 32640 8888 32646 8900
rect 33594 8888 33600 8900
rect 32640 8860 33600 8888
rect 32640 8848 32646 8860
rect 33594 8848 33600 8860
rect 33652 8888 33658 8900
rect 33781 8891 33839 8897
rect 33781 8888 33793 8891
rect 33652 8860 33793 8888
rect 33652 8848 33658 8860
rect 33781 8857 33793 8860
rect 33827 8857 33839 8891
rect 35986 8888 35992 8900
rect 35947 8860 35992 8888
rect 33781 8851 33839 8857
rect 35986 8848 35992 8860
rect 36044 8848 36050 8900
rect 25556 8792 26556 8820
rect 25556 8780 25562 8792
rect 26602 8780 26608 8832
rect 26660 8820 26666 8832
rect 30282 8820 30288 8832
rect 26660 8792 30288 8820
rect 26660 8780 26666 8792
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 30926 8780 30932 8832
rect 30984 8820 30990 8832
rect 31312 8820 31340 8848
rect 30984 8792 31340 8820
rect 30984 8780 30990 8792
rect 32122 8780 32128 8832
rect 32180 8820 32186 8832
rect 37461 8823 37519 8829
rect 37461 8820 37473 8823
rect 32180 8792 37473 8820
rect 32180 8780 32186 8792
rect 37461 8789 37473 8792
rect 37507 8789 37519 8823
rect 37461 8783 37519 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 13354 8616 13360 8628
rect 13267 8588 13360 8616
rect 13354 8576 13360 8588
rect 13412 8616 13418 8628
rect 15286 8616 15292 8628
rect 13412 8588 15292 8616
rect 13412 8576 13418 8588
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15838 8616 15844 8628
rect 15611 8588 15844 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 17218 8616 17224 8628
rect 16255 8588 17224 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 20349 8619 20407 8625
rect 17788 8588 18092 8616
rect 13906 8548 13912 8560
rect 13867 8520 13912 8548
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 14461 8551 14519 8557
rect 14461 8517 14473 8551
rect 14507 8548 14519 8551
rect 17586 8548 17592 8560
rect 14507 8520 17592 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 13924 8412 13952 8508
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 16132 8489 16160 8520
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 17788 8548 17816 8588
rect 17696 8520 17816 8548
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 14700 8452 15485 8480
rect 14700 8440 14706 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 16117 8443 16175 8449
rect 14826 8412 14832 8424
rect 13924 8384 14832 8412
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 15488 8412 15516 8443
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17696 8480 17724 8520
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 17957 8551 18015 8557
rect 17957 8548 17969 8551
rect 17920 8520 17969 8548
rect 17920 8508 17926 8520
rect 17957 8517 17969 8520
rect 18003 8517 18015 8551
rect 18064 8548 18092 8588
rect 20349 8585 20361 8619
rect 20395 8616 20407 8619
rect 20806 8616 20812 8628
rect 20395 8588 20812 8616
rect 20395 8585 20407 8588
rect 20349 8579 20407 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21634 8616 21640 8628
rect 21407 8588 21640 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 22097 8619 22155 8625
rect 22097 8585 22109 8619
rect 22143 8616 22155 8619
rect 23290 8616 23296 8628
rect 22143 8588 23296 8616
rect 22143 8585 22155 8588
rect 22097 8579 22155 8585
rect 23290 8576 23296 8588
rect 23348 8576 23354 8628
rect 25590 8576 25596 8628
rect 25648 8616 25654 8628
rect 27249 8619 27307 8625
rect 27249 8616 27261 8619
rect 25648 8588 27261 8616
rect 25648 8576 25654 8588
rect 27249 8585 27261 8588
rect 27295 8585 27307 8619
rect 27249 8579 27307 8585
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 27764 8588 29684 8616
rect 27764 8576 27770 8588
rect 19334 8548 19340 8560
rect 18064 8520 19340 8548
rect 17957 8511 18015 8517
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 19613 8551 19671 8557
rect 19613 8517 19625 8551
rect 19659 8548 19671 8551
rect 20714 8548 20720 8560
rect 19659 8520 20720 8548
rect 19659 8517 19671 8520
rect 19613 8511 19671 8517
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 21082 8508 21088 8560
rect 21140 8548 21146 8560
rect 21726 8548 21732 8560
rect 21140 8520 21732 8548
rect 21140 8508 21146 8520
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 22186 8508 22192 8560
rect 22244 8548 22250 8560
rect 23569 8551 23627 8557
rect 22244 8520 22402 8548
rect 22244 8508 22250 8520
rect 23569 8517 23581 8551
rect 23615 8548 23627 8551
rect 23658 8548 23664 8560
rect 23615 8520 23664 8548
rect 23615 8517 23627 8520
rect 23569 8511 23627 8517
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 25038 8508 25044 8560
rect 25096 8508 25102 8560
rect 27724 8548 27752 8576
rect 29546 8548 29552 8560
rect 25884 8520 27752 8548
rect 29302 8520 29552 8548
rect 17236 8452 17724 8480
rect 20257 8483 20315 8489
rect 17236 8412 17264 8452
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 20346 8480 20352 8492
rect 20303 8452 20352 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 22278 8480 22284 8492
rect 20680 8452 22284 8480
rect 20680 8440 20686 8452
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 24305 8483 24363 8489
rect 24305 8480 24317 8483
rect 23900 8452 24317 8480
rect 23900 8440 23906 8452
rect 24305 8449 24317 8452
rect 24351 8449 24363 8483
rect 24305 8443 24363 8449
rect 15488 8384 17264 8412
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 17865 8415 17923 8421
rect 17865 8412 17877 8415
rect 17736 8384 17877 8412
rect 17736 8372 17742 8384
rect 17865 8381 17877 8384
rect 17911 8381 17923 8415
rect 19610 8412 19616 8424
rect 17865 8375 17923 8381
rect 18340 8384 19616 8412
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 14090 8344 14096 8356
rect 13688 8316 14096 8344
rect 13688 8304 13694 8316
rect 14090 8304 14096 8316
rect 14148 8344 14154 8356
rect 14921 8347 14979 8353
rect 14921 8344 14933 8347
rect 14148 8316 14933 8344
rect 14148 8304 14154 8316
rect 14921 8313 14933 8316
rect 14967 8344 14979 8347
rect 17126 8344 17132 8356
rect 14967 8316 17132 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17221 8347 17279 8353
rect 17221 8313 17233 8347
rect 17267 8344 17279 8347
rect 18340 8344 18368 8384
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8412 19763 8415
rect 20162 8412 20168 8424
rect 19751 8384 20168 8412
rect 19751 8381 19763 8384
rect 19705 8375 19763 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 21450 8372 21456 8424
rect 21508 8412 21514 8424
rect 21726 8412 21732 8424
rect 21508 8384 21732 8412
rect 21508 8372 21514 8384
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 21910 8372 21916 8424
rect 21968 8412 21974 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 21968 8384 24593 8412
rect 21968 8372 21974 8384
rect 24581 8381 24593 8384
rect 24627 8381 24639 8415
rect 24581 8375 24639 8381
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 25884 8412 25912 8520
rect 29546 8508 29552 8520
rect 29604 8508 29610 8560
rect 29656 8548 29684 8588
rect 30377 8551 30435 8557
rect 29656 8520 29960 8548
rect 27338 8480 27344 8492
rect 27299 8452 27344 8480
rect 27338 8440 27344 8452
rect 27396 8440 27402 8492
rect 29362 8440 29368 8492
rect 29420 8480 29426 8492
rect 29420 8452 29868 8480
rect 29420 8440 29426 8452
rect 24728 8384 25912 8412
rect 26053 8415 26111 8421
rect 24728 8372 24734 8384
rect 26053 8381 26065 8415
rect 26099 8412 26111 8415
rect 26878 8412 26884 8424
rect 26099 8384 26884 8412
rect 26099 8381 26111 8384
rect 26053 8375 26111 8381
rect 26878 8372 26884 8384
rect 26936 8372 26942 8424
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 27801 8415 27859 8421
rect 27801 8412 27813 8415
rect 27580 8384 27813 8412
rect 27580 8372 27586 8384
rect 27801 8381 27813 8384
rect 27847 8381 27859 8415
rect 27801 8375 27859 8381
rect 28077 8415 28135 8421
rect 28077 8381 28089 8415
rect 28123 8412 28135 8415
rect 29270 8412 29276 8424
rect 28123 8384 29276 8412
rect 28123 8381 28135 8384
rect 28077 8375 28135 8381
rect 29270 8372 29276 8384
rect 29328 8372 29334 8424
rect 29840 8421 29868 8452
rect 29825 8415 29883 8421
rect 29825 8381 29837 8415
rect 29871 8381 29883 8415
rect 29932 8412 29960 8520
rect 30377 8517 30389 8551
rect 30423 8548 30435 8551
rect 30558 8548 30564 8560
rect 30423 8520 30564 8548
rect 30423 8517 30435 8520
rect 30377 8511 30435 8517
rect 30558 8508 30564 8520
rect 30616 8508 30622 8560
rect 30282 8480 30288 8492
rect 30243 8452 30288 8480
rect 30282 8440 30288 8452
rect 30340 8440 30346 8492
rect 36814 8440 36820 8492
rect 36872 8480 36878 8492
rect 37737 8483 37795 8489
rect 37737 8480 37749 8483
rect 36872 8452 37749 8480
rect 36872 8440 36878 8452
rect 37737 8449 37749 8452
rect 37783 8449 37795 8483
rect 37737 8443 37795 8449
rect 31481 8415 31539 8421
rect 31481 8412 31493 8415
rect 29932 8384 31493 8412
rect 29825 8375 29883 8381
rect 31481 8381 31493 8384
rect 31527 8381 31539 8415
rect 31481 8375 31539 8381
rect 36909 8415 36967 8421
rect 36909 8381 36921 8415
rect 36955 8412 36967 8415
rect 37182 8412 37188 8424
rect 36955 8384 37188 8412
rect 36955 8381 36967 8384
rect 36909 8375 36967 8381
rect 17267 8316 18368 8344
rect 18417 8347 18475 8353
rect 17267 8313 17279 8316
rect 17221 8307 17279 8313
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 19150 8344 19156 8356
rect 18463 8316 19156 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 6822 8276 6828 8288
rect 2096 8248 6828 8276
rect 2096 8236 2102 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 18432 8276 18460 8307
rect 19150 8304 19156 8316
rect 19208 8304 19214 8356
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 22554 8344 22560 8356
rect 19392 8316 22560 8344
rect 19392 8304 19398 8316
rect 22554 8304 22560 8316
rect 22612 8304 22618 8356
rect 29546 8344 29552 8356
rect 29196 8316 29552 8344
rect 15068 8248 18460 8276
rect 15068 8236 15074 8248
rect 19242 8236 19248 8288
rect 19300 8276 19306 8288
rect 20622 8276 20628 8288
rect 19300 8248 20628 8276
rect 19300 8236 19306 8248
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 21450 8236 21456 8288
rect 21508 8276 21514 8288
rect 25774 8276 25780 8288
rect 21508 8248 25780 8276
rect 21508 8236 21514 8248
rect 25774 8236 25780 8248
rect 25832 8236 25838 8288
rect 25866 8236 25872 8288
rect 25924 8276 25930 8288
rect 28626 8276 28632 8288
rect 25924 8248 28632 8276
rect 25924 8236 25930 8248
rect 28626 8236 28632 8248
rect 28684 8236 28690 8288
rect 28718 8236 28724 8288
rect 28776 8276 28782 8288
rect 29196 8276 29224 8316
rect 29546 8304 29552 8316
rect 29604 8304 29610 8356
rect 28776 8248 29224 8276
rect 28776 8236 28782 8248
rect 29270 8236 29276 8288
rect 29328 8276 29334 8288
rect 29730 8276 29736 8288
rect 29328 8248 29736 8276
rect 29328 8236 29334 8248
rect 29730 8236 29736 8248
rect 29788 8236 29794 8288
rect 29840 8276 29868 8375
rect 37182 8372 37188 8384
rect 37240 8412 37246 8424
rect 37461 8415 37519 8421
rect 37461 8412 37473 8415
rect 37240 8384 37473 8412
rect 37240 8372 37246 8384
rect 37461 8381 37473 8384
rect 37507 8381 37519 8415
rect 37461 8375 37519 8381
rect 30834 8304 30840 8356
rect 30892 8344 30898 8356
rect 30929 8347 30987 8353
rect 30929 8344 30941 8347
rect 30892 8316 30941 8344
rect 30892 8304 30898 8316
rect 30929 8313 30941 8316
rect 30975 8344 30987 8347
rect 31570 8344 31576 8356
rect 30975 8316 31576 8344
rect 30975 8313 30987 8316
rect 30929 8307 30987 8313
rect 31570 8304 31576 8316
rect 31628 8344 31634 8356
rect 32309 8347 32367 8353
rect 32309 8344 32321 8347
rect 31628 8316 32321 8344
rect 31628 8304 31634 8316
rect 32309 8313 32321 8316
rect 32355 8344 32367 8347
rect 32582 8344 32588 8356
rect 32355 8316 32588 8344
rect 32355 8313 32367 8316
rect 32309 8307 32367 8313
rect 32582 8304 32588 8316
rect 32640 8344 32646 8356
rect 32861 8347 32919 8353
rect 32861 8344 32873 8347
rect 32640 8316 32873 8344
rect 32640 8304 32646 8316
rect 32861 8313 32873 8316
rect 32907 8344 32919 8347
rect 33413 8347 33471 8353
rect 33413 8344 33425 8347
rect 32907 8316 33425 8344
rect 32907 8313 32919 8316
rect 32861 8307 32919 8313
rect 33413 8313 33425 8316
rect 33459 8313 33471 8347
rect 33413 8307 33471 8313
rect 34057 8347 34115 8353
rect 34057 8313 34069 8347
rect 34103 8344 34115 8347
rect 34514 8344 34520 8356
rect 34103 8316 34520 8344
rect 34103 8313 34115 8316
rect 34057 8307 34115 8313
rect 34514 8304 34520 8316
rect 34572 8304 34578 8356
rect 36354 8344 36360 8356
rect 36315 8316 36360 8344
rect 36354 8304 36360 8316
rect 36412 8304 36418 8356
rect 33594 8276 33600 8288
rect 29840 8248 33600 8276
rect 33594 8236 33600 8248
rect 33652 8236 33658 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 18138 8072 18144 8084
rect 12759 8044 18144 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 19058 8072 19064 8084
rect 18831 8044 19064 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19610 8032 19616 8084
rect 19668 8072 19674 8084
rect 20162 8072 20168 8084
rect 19668 8044 20168 8072
rect 19668 8032 19674 8044
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20714 8072 20720 8084
rect 20675 8044 20720 8072
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 21637 8075 21695 8081
rect 21637 8041 21649 8075
rect 21683 8072 21695 8075
rect 21910 8072 21916 8084
rect 21683 8044 21916 8072
rect 21683 8041 21695 8044
rect 21637 8035 21695 8041
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 22060 8044 23949 8072
rect 22060 8032 22066 8044
rect 23937 8041 23949 8044
rect 23983 8041 23995 8075
rect 23937 8035 23995 8041
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 24360 8044 25452 8072
rect 24360 8032 24366 8044
rect 13357 8007 13415 8013
rect 13357 7973 13369 8007
rect 13403 8004 13415 8007
rect 16574 8004 16580 8016
rect 13403 7976 16580 8004
rect 13403 7973 13415 7976
rect 13357 7967 13415 7973
rect 16574 7964 16580 7976
rect 16632 7964 16638 8016
rect 16868 7976 18828 8004
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 15194 7936 15200 7948
rect 14415 7908 15200 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 16390 7936 16396 7948
rect 15703 7908 16396 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16868 7945 16896 7976
rect 18800 7948 18828 7976
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 18932 7976 22140 8004
rect 18932 7964 18938 7976
rect 16853 7939 16911 7945
rect 16853 7905 16865 7939
rect 16899 7905 16911 7939
rect 17770 7936 17776 7948
rect 17731 7908 17776 7936
rect 16853 7899 16911 7905
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7936 18199 7939
rect 18414 7936 18420 7948
rect 18187 7908 18420 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 18782 7896 18788 7948
rect 18840 7896 18846 7948
rect 20073 7939 20131 7945
rect 20073 7905 20085 7939
rect 20119 7936 20131 7939
rect 21450 7936 21456 7948
rect 20119 7908 21456 7936
rect 20119 7905 20131 7908
rect 20073 7899 20131 7905
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 22112 7936 22140 7976
rect 23308 7976 25360 8004
rect 23308 7936 23336 7976
rect 22112 7908 23336 7936
rect 23385 7939 23443 7945
rect 23385 7905 23397 7939
rect 23431 7936 23443 7939
rect 23474 7936 23480 7948
rect 23431 7908 23480 7936
rect 23431 7905 23443 7908
rect 23385 7899 23443 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 12492 7840 12633 7868
rect 12492 7828 12498 7840
rect 12621 7837 12633 7840
rect 12667 7868 12679 7871
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12667 7840 13277 7868
rect 12667 7837 12679 7840
rect 12621 7831 12679 7837
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15068 7840 15113 7868
rect 15068 7828 15074 7840
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15344 7840 15577 7868
rect 15344 7828 15350 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19242 7868 19248 7880
rect 18923 7840 19248 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 21174 7868 21180 7880
rect 20855 7840 21180 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 24026 7868 24032 7880
rect 23987 7840 24032 7868
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 25332 7854 25360 7976
rect 25424 7936 25452 8044
rect 28258 8032 28264 8084
rect 28316 8072 28322 8084
rect 28917 8075 28975 8081
rect 28917 8072 28929 8075
rect 28316 8044 28929 8072
rect 28316 8032 28322 8044
rect 28917 8041 28929 8044
rect 28963 8072 28975 8075
rect 35989 8075 36047 8081
rect 28963 8044 31754 8072
rect 28963 8041 28975 8044
rect 28917 8035 28975 8041
rect 27433 8007 27491 8013
rect 27433 8004 27445 8007
rect 26620 7976 27445 8004
rect 26421 7939 26479 7945
rect 26421 7936 26433 7939
rect 25424 7908 26433 7936
rect 26421 7905 26433 7908
rect 26467 7936 26479 7939
rect 26620 7936 26648 7976
rect 27433 7973 27445 7976
rect 27479 7973 27491 8007
rect 27433 7967 27491 7973
rect 31202 7964 31208 8016
rect 31260 8004 31266 8016
rect 31481 8007 31539 8013
rect 31481 8004 31493 8007
rect 31260 7976 31493 8004
rect 31260 7964 31266 7976
rect 31481 7973 31493 7976
rect 31527 7973 31539 8007
rect 31726 8004 31754 8044
rect 35989 8041 36001 8075
rect 36035 8072 36047 8075
rect 36078 8072 36084 8084
rect 36035 8044 36084 8072
rect 36035 8041 36047 8044
rect 35989 8035 36047 8041
rect 36078 8032 36084 8044
rect 36136 8032 36142 8084
rect 33045 8007 33103 8013
rect 33045 8004 33057 8007
rect 31726 7976 33057 8004
rect 31481 7967 31539 7973
rect 33045 7973 33057 7976
rect 33091 7973 33103 8007
rect 37921 8007 37979 8013
rect 37921 8004 37933 8007
rect 33045 7967 33103 7973
rect 34808 7976 37933 8004
rect 27522 7936 27528 7948
rect 26467 7908 26648 7936
rect 26712 7908 27528 7936
rect 26467 7905 26479 7908
rect 26421 7899 26479 7905
rect 26712 7880 26740 7908
rect 27522 7896 27528 7908
rect 27580 7936 27586 7948
rect 30009 7939 30067 7945
rect 27580 7908 29224 7936
rect 27580 7896 27586 7908
rect 26694 7828 26700 7880
rect 26752 7868 26758 7880
rect 29196 7877 29224 7908
rect 30009 7905 30021 7939
rect 30055 7936 30067 7939
rect 30374 7936 30380 7948
rect 30055 7908 30380 7936
rect 30055 7905 30067 7908
rect 30009 7899 30067 7905
rect 30374 7896 30380 7908
rect 30432 7896 30438 7948
rect 34808 7936 34836 7976
rect 37921 7973 37933 7976
rect 37967 7973 37979 8007
rect 37921 7967 37979 7973
rect 36630 7936 36636 7948
rect 31128 7908 34836 7936
rect 36591 7908 36636 7936
rect 29181 7871 29239 7877
rect 26752 7840 26797 7868
rect 26752 7828 26758 7840
rect 29181 7837 29193 7871
rect 29227 7868 29239 7871
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29227 7840 29745 7868
rect 29227 7837 29239 7840
rect 29181 7831 29239 7837
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 31128 7854 31156 7908
rect 36630 7896 36636 7908
rect 36688 7896 36694 7948
rect 35437 7871 35495 7877
rect 29733 7831 29791 7837
rect 35437 7837 35449 7871
rect 35483 7868 35495 7871
rect 36078 7868 36084 7880
rect 35483 7840 36084 7868
rect 35483 7837 35495 7840
rect 35437 7831 35495 7837
rect 36078 7828 36084 7840
rect 36136 7828 36142 7880
rect 36648 7868 36676 7896
rect 37185 7871 37243 7877
rect 37185 7868 37197 7871
rect 36648 7840 37197 7868
rect 37185 7837 37197 7840
rect 37231 7837 37243 7871
rect 37826 7868 37832 7880
rect 37787 7840 37832 7868
rect 37185 7831 37243 7837
rect 37826 7828 37832 7840
rect 37884 7828 37890 7880
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 14476 7732 14504 7763
rect 14550 7760 14556 7812
rect 14608 7800 14614 7812
rect 16114 7800 16120 7812
rect 14608 7772 16120 7800
rect 14608 7760 14614 7772
rect 16114 7760 16120 7772
rect 16172 7800 16178 7812
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 16172 7772 16221 7800
rect 16172 7760 16178 7772
rect 16209 7769 16221 7772
rect 16255 7769 16267 7803
rect 16209 7763 16267 7769
rect 16390 7760 16396 7812
rect 16448 7800 16454 7812
rect 16761 7803 16819 7809
rect 16761 7800 16773 7803
rect 16448 7772 16773 7800
rect 16448 7760 16454 7772
rect 16761 7769 16773 7772
rect 16807 7769 16819 7803
rect 18049 7803 18107 7809
rect 18049 7800 18061 7803
rect 16761 7763 16819 7769
rect 16868 7772 18061 7800
rect 13504 7704 14504 7732
rect 13504 7692 13510 7704
rect 14642 7692 14648 7744
rect 14700 7732 14706 7744
rect 16868 7732 16896 7772
rect 18049 7769 18061 7772
rect 18095 7769 18107 7803
rect 18049 7763 18107 7769
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 18840 7772 19441 7800
rect 18840 7760 18846 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 19978 7800 19984 7812
rect 19939 7772 19984 7800
rect 19429 7763 19487 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 22646 7760 22652 7812
rect 22704 7760 22710 7812
rect 23014 7760 23020 7812
rect 23072 7800 23078 7812
rect 23109 7803 23167 7809
rect 23109 7800 23121 7803
rect 23072 7772 23121 7800
rect 23072 7760 23078 7772
rect 23109 7769 23121 7772
rect 23155 7769 23167 7803
rect 23109 7763 23167 7769
rect 24673 7803 24731 7809
rect 24673 7769 24685 7803
rect 24719 7800 24731 7803
rect 25038 7800 25044 7812
rect 24719 7772 25044 7800
rect 24719 7769 24731 7772
rect 24673 7763 24731 7769
rect 14700 7704 16896 7732
rect 14700 7692 14706 7704
rect 18138 7692 18144 7744
rect 18196 7732 18202 7744
rect 20806 7732 20812 7744
rect 18196 7704 20812 7732
rect 18196 7692 18202 7704
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 20898 7692 20904 7744
rect 20956 7732 20962 7744
rect 21634 7732 21640 7744
rect 20956 7704 21640 7732
rect 20956 7692 20962 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 24688 7732 24716 7763
rect 25038 7760 25044 7772
rect 25096 7760 25102 7812
rect 26326 7760 26332 7812
rect 26384 7800 26390 7812
rect 26384 7772 27738 7800
rect 26384 7760 26390 7772
rect 28626 7760 28632 7812
rect 28684 7800 28690 7812
rect 29454 7800 29460 7812
rect 28684 7772 29460 7800
rect 28684 7760 28690 7772
rect 29454 7760 29460 7772
rect 29512 7760 29518 7812
rect 31294 7760 31300 7812
rect 31352 7800 31358 7812
rect 35345 7803 35403 7809
rect 35345 7800 35357 7803
rect 31352 7772 35357 7800
rect 31352 7760 31358 7772
rect 35345 7769 35357 7772
rect 35391 7769 35403 7803
rect 35345 7763 35403 7769
rect 22796 7704 24716 7732
rect 22796 7692 22802 7704
rect 26234 7692 26240 7744
rect 26292 7732 26298 7744
rect 31478 7732 31484 7744
rect 26292 7704 31484 7732
rect 26292 7692 26298 7704
rect 31478 7692 31484 7704
rect 31536 7692 31542 7744
rect 31938 7732 31944 7744
rect 31899 7704 31944 7732
rect 31938 7692 31944 7704
rect 31996 7692 32002 7744
rect 32585 7735 32643 7741
rect 32585 7701 32597 7735
rect 32631 7732 32643 7735
rect 33410 7732 33416 7744
rect 32631 7704 33416 7732
rect 32631 7701 32643 7704
rect 32585 7695 32643 7701
rect 33410 7692 33416 7704
rect 33468 7732 33474 7744
rect 33597 7735 33655 7741
rect 33597 7732 33609 7735
rect 33468 7704 33609 7732
rect 33468 7692 33474 7704
rect 33597 7701 33609 7704
rect 33643 7701 33655 7735
rect 33597 7695 33655 7701
rect 37369 7735 37427 7741
rect 37369 7701 37381 7735
rect 37415 7732 37427 7735
rect 37458 7732 37464 7744
rect 37415 7704 37464 7732
rect 37415 7701 37427 7704
rect 37369 7695 37427 7701
rect 37458 7692 37464 7704
rect 37516 7692 37522 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 14642 7528 14648 7540
rect 13679 7500 14648 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 16390 7528 16396 7540
rect 14967 7500 16396 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 19150 7528 19156 7540
rect 16632 7500 19156 7528
rect 16632 7488 16638 7500
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19610 7488 19616 7540
rect 19668 7528 19674 7540
rect 26326 7528 26332 7540
rect 19668 7500 26332 7528
rect 19668 7488 19674 7500
rect 26326 7488 26332 7500
rect 26384 7488 26390 7540
rect 26878 7488 26884 7540
rect 26936 7528 26942 7540
rect 26936 7500 28304 7528
rect 26936 7488 26942 7500
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2038 7460 2044 7472
rect 1903 7432 2044 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2038 7420 2044 7432
rect 2096 7420 2102 7472
rect 15286 7460 15292 7472
rect 14200 7432 15292 7460
rect 14200 7404 14228 7432
rect 15286 7420 15292 7432
rect 15344 7460 15350 7472
rect 16209 7463 16267 7469
rect 15344 7432 15516 7460
rect 15344 7420 15350 7432
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 12492 7364 12633 7392
rect 12492 7352 12498 7364
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7392 13599 7395
rect 13814 7392 13820 7404
rect 13587 7364 13820 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 13556 7324 13584 7355
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 14182 7392 14188 7404
rect 14143 7364 14188 7392
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 15488 7401 15516 7432
rect 16209 7429 16221 7463
rect 16255 7460 16267 7463
rect 16666 7460 16672 7472
rect 16255 7432 16672 7460
rect 16255 7429 16267 7432
rect 16209 7423 16267 7429
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 16942 7460 16948 7472
rect 16903 7432 16948 7460
rect 16942 7420 16948 7432
rect 17000 7420 17006 7472
rect 17037 7463 17095 7469
rect 17037 7429 17049 7463
rect 17083 7460 17095 7463
rect 17126 7460 17132 7472
rect 17083 7432 17132 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 17126 7420 17132 7432
rect 17184 7420 17190 7472
rect 19334 7420 19340 7472
rect 19392 7460 19398 7472
rect 19521 7463 19579 7469
rect 19521 7460 19533 7463
rect 19392 7432 19533 7460
rect 19392 7420 19398 7432
rect 19521 7429 19533 7432
rect 19567 7429 19579 7463
rect 19521 7423 19579 7429
rect 20162 7420 20168 7472
rect 20220 7460 20226 7472
rect 20220 7432 22586 7460
rect 20220 7420 20226 7432
rect 23474 7420 23480 7472
rect 23532 7460 23538 7472
rect 23842 7460 23848 7472
rect 23532 7432 23848 7460
rect 23532 7420 23538 7432
rect 23842 7420 23848 7432
rect 23900 7460 23906 7472
rect 24486 7460 24492 7472
rect 23900 7432 24072 7460
rect 24447 7432 24492 7460
rect 23900 7420 23906 7432
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16022 7392 16028 7404
rect 15611 7364 16028 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16390 7392 16396 7404
rect 16347 7364 16396 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 17586 7352 17592 7404
rect 17644 7392 17650 7404
rect 18325 7395 18383 7401
rect 18325 7392 18337 7395
rect 17644 7364 18337 7392
rect 17644 7352 17650 7364
rect 18325 7361 18337 7364
rect 18371 7361 18383 7395
rect 18325 7355 18383 7361
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 21266 7392 21272 7404
rect 19852 7364 21272 7392
rect 19852 7352 19858 7364
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 24044 7401 24072 7432
rect 24486 7420 24492 7432
rect 24544 7420 24550 7472
rect 27246 7460 27252 7472
rect 25806 7432 27252 7460
rect 27246 7420 27252 7432
rect 27304 7420 27310 7472
rect 28276 7469 28304 7500
rect 28350 7488 28356 7540
rect 28408 7528 28414 7540
rect 29733 7531 29791 7537
rect 29733 7528 29745 7531
rect 28408 7500 29745 7528
rect 28408 7488 28414 7500
rect 29733 7497 29745 7500
rect 29779 7528 29791 7531
rect 30650 7528 30656 7540
rect 29779 7500 30656 7528
rect 29779 7497 29791 7500
rect 29733 7491 29791 7497
rect 30650 7488 30656 7500
rect 30708 7488 30714 7540
rect 34790 7488 34796 7540
rect 34848 7528 34854 7540
rect 35069 7531 35127 7537
rect 35069 7528 35081 7531
rect 34848 7500 35081 7528
rect 34848 7488 34854 7500
rect 35069 7497 35081 7500
rect 35115 7528 35127 7531
rect 35526 7528 35532 7540
rect 35115 7500 35532 7528
rect 35115 7497 35127 7500
rect 35069 7491 35127 7497
rect 35526 7488 35532 7500
rect 35584 7488 35590 7540
rect 36078 7488 36084 7540
rect 36136 7528 36142 7540
rect 36265 7531 36323 7537
rect 36265 7528 36277 7531
rect 36136 7500 36277 7528
rect 36136 7488 36142 7500
rect 36265 7497 36277 7500
rect 36311 7497 36323 7531
rect 36265 7491 36323 7497
rect 28261 7463 28319 7469
rect 28261 7429 28273 7463
rect 28307 7429 28319 7463
rect 28261 7423 28319 7429
rect 28994 7420 29000 7472
rect 29052 7420 29058 7472
rect 29546 7420 29552 7472
rect 29604 7460 29610 7472
rect 30193 7463 30251 7469
rect 30193 7460 30205 7463
rect 29604 7432 30205 7460
rect 29604 7420 29610 7432
rect 30193 7429 30205 7432
rect 30239 7429 30251 7463
rect 30193 7423 30251 7429
rect 33134 7420 33140 7472
rect 33192 7460 33198 7472
rect 36817 7463 36875 7469
rect 36817 7460 36829 7463
rect 33192 7432 36829 7460
rect 33192 7420 33198 7432
rect 36817 7429 36829 7432
rect 36863 7460 36875 7463
rect 37550 7460 37556 7472
rect 36863 7432 37556 7460
rect 36863 7429 36875 7432
rect 36817 7423 36875 7429
rect 37550 7420 37556 7432
rect 37608 7460 37614 7472
rect 37608 7432 37688 7460
rect 37608 7420 37614 7432
rect 24029 7395 24087 7401
rect 21508 7364 22600 7392
rect 21508 7352 21514 7364
rect 12207 7296 13584 7324
rect 14277 7327 14335 7333
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 19518 7324 19524 7336
rect 14323 7296 19524 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 19518 7284 19524 7296
rect 19576 7284 19582 7336
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 19886 7324 19892 7336
rect 19659 7296 19892 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 20162 7312 20168 7336
rect 19996 7284 20168 7312
rect 20220 7284 20226 7336
rect 22005 7327 22063 7333
rect 22005 7293 22017 7327
rect 22051 7324 22063 7327
rect 22094 7324 22100 7336
rect 22051 7296 22100 7324
rect 22051 7293 22063 7296
rect 22005 7287 22063 7293
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22572 7324 22600 7364
rect 24029 7361 24041 7395
rect 24075 7361 24087 7395
rect 24029 7355 24087 7361
rect 26786 7352 26792 7404
rect 26844 7392 26850 7404
rect 27154 7392 27160 7404
rect 26844 7364 27160 7392
rect 26844 7352 26850 7364
rect 27154 7352 27160 7364
rect 27212 7352 27218 7404
rect 37660 7401 37688 7432
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7392 37703 7395
rect 38105 7395 38163 7401
rect 38105 7392 38117 7395
rect 37691 7364 38117 7392
rect 37691 7361 37703 7364
rect 37645 7355 37703 7361
rect 38105 7361 38117 7364
rect 38151 7392 38163 7395
rect 38194 7392 38200 7404
rect 38151 7364 38200 7392
rect 38151 7361 38163 7364
rect 38105 7355 38163 7361
rect 38194 7352 38200 7364
rect 38252 7352 38258 7404
rect 23658 7324 23664 7336
rect 22572 7296 23664 7324
rect 23658 7284 23664 7296
rect 23716 7284 23722 7336
rect 23753 7327 23811 7333
rect 23753 7293 23765 7327
rect 23799 7324 23811 7327
rect 25866 7324 25872 7336
rect 23799 7296 25872 7324
rect 23799 7293 23811 7296
rect 23753 7287 23811 7293
rect 25866 7284 25872 7296
rect 25924 7284 25930 7336
rect 26234 7324 26240 7336
rect 26195 7296 26240 7324
rect 26234 7284 26240 7296
rect 26292 7284 26298 7336
rect 26513 7327 26571 7333
rect 26513 7293 26525 7327
rect 26559 7324 26571 7327
rect 26602 7324 26608 7336
rect 26559 7296 26608 7324
rect 26559 7293 26571 7296
rect 26513 7287 26571 7293
rect 26602 7284 26608 7296
rect 26660 7324 26666 7336
rect 27985 7327 28043 7333
rect 27985 7324 27997 7327
rect 26660 7296 27997 7324
rect 26660 7284 26666 7296
rect 27985 7293 27997 7296
rect 28031 7293 28043 7327
rect 31389 7327 31447 7333
rect 31389 7324 31401 7327
rect 27985 7287 28043 7293
rect 28092 7296 31401 7324
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 17034 7256 17040 7268
rect 16724 7228 17040 7256
rect 16724 7216 16730 7228
rect 17034 7216 17040 7228
rect 17092 7216 17098 7268
rect 17497 7259 17555 7265
rect 17497 7225 17509 7259
rect 17543 7256 17555 7259
rect 17770 7256 17776 7268
rect 17543 7228 17776 7256
rect 17543 7225 17555 7228
rect 17497 7219 17555 7225
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 18874 7256 18880 7268
rect 17880 7228 18880 7256
rect 12713 7191 12771 7197
rect 12713 7157 12725 7191
rect 12759 7188 12771 7191
rect 12802 7188 12808 7200
rect 12759 7160 12808 7188
rect 12759 7157 12771 7160
rect 12713 7151 12771 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 17880 7188 17908 7228
rect 18874 7216 18880 7228
rect 18932 7256 18938 7268
rect 19061 7259 19119 7265
rect 19061 7256 19073 7259
rect 18932 7228 19073 7256
rect 18932 7216 18938 7228
rect 19061 7225 19073 7228
rect 19107 7225 19119 7259
rect 19061 7219 19119 7225
rect 19242 7216 19248 7268
rect 19300 7256 19306 7268
rect 19996 7256 20024 7284
rect 19300 7228 20024 7256
rect 19300 7216 19306 7228
rect 21174 7216 21180 7268
rect 21232 7256 21238 7268
rect 22462 7256 22468 7268
rect 21232 7228 22468 7256
rect 21232 7216 21238 7228
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 27249 7259 27307 7265
rect 27249 7225 27261 7259
rect 27295 7256 27307 7259
rect 27430 7256 27436 7268
rect 27295 7228 27436 7256
rect 27295 7225 27307 7228
rect 27249 7219 27307 7225
rect 27430 7216 27436 7228
rect 27488 7216 27494 7268
rect 27522 7216 27528 7268
rect 27580 7256 27586 7268
rect 28092 7256 28120 7296
rect 31389 7293 31401 7296
rect 31435 7324 31447 7327
rect 31938 7324 31944 7336
rect 31435 7296 31944 7324
rect 31435 7293 31447 7296
rect 31389 7287 31447 7293
rect 31938 7284 31944 7296
rect 31996 7324 32002 7336
rect 34606 7324 34612 7336
rect 31996 7296 34612 7324
rect 31996 7284 32002 7296
rect 34606 7284 34612 7296
rect 34664 7284 34670 7336
rect 34698 7284 34704 7336
rect 34756 7324 34762 7336
rect 37553 7327 37611 7333
rect 37553 7324 37565 7327
rect 34756 7296 37565 7324
rect 34756 7284 34762 7296
rect 37553 7293 37565 7296
rect 37599 7293 37611 7327
rect 37553 7287 37611 7293
rect 30650 7256 30656 7268
rect 27580 7228 28120 7256
rect 30116 7228 30656 7256
rect 27580 7216 27586 7228
rect 16172 7160 17908 7188
rect 18417 7191 18475 7197
rect 16172 7148 16178 7160
rect 18417 7157 18429 7191
rect 18463 7188 18475 7191
rect 19610 7188 19616 7200
rect 18463 7160 19616 7188
rect 18463 7157 18475 7160
rect 18417 7151 18475 7157
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 20346 7148 20352 7200
rect 20404 7188 20410 7200
rect 20901 7191 20959 7197
rect 20404 7160 20449 7188
rect 20404 7148 20410 7160
rect 20901 7157 20913 7191
rect 20947 7188 20959 7191
rect 21082 7188 21088 7200
rect 20947 7160 21088 7188
rect 20947 7157 20959 7160
rect 20901 7151 20959 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 21358 7188 21364 7200
rect 21319 7160 21364 7188
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 28994 7148 29000 7200
rect 29052 7188 29058 7200
rect 30116 7188 30144 7228
rect 30650 7216 30656 7228
rect 30708 7256 30714 7268
rect 31570 7256 31576 7268
rect 30708 7228 31576 7256
rect 30708 7216 30714 7228
rect 31570 7216 31576 7228
rect 31628 7216 31634 7268
rect 32030 7216 32036 7268
rect 32088 7256 32094 7268
rect 32401 7259 32459 7265
rect 32401 7256 32413 7259
rect 32088 7228 32413 7256
rect 32088 7216 32094 7228
rect 32401 7225 32413 7228
rect 32447 7256 32459 7259
rect 32953 7259 33011 7265
rect 32953 7256 32965 7259
rect 32447 7228 32965 7256
rect 32447 7225 32459 7228
rect 32401 7219 32459 7225
rect 32953 7225 32965 7228
rect 32999 7256 33011 7259
rect 33410 7256 33416 7268
rect 32999 7228 33416 7256
rect 32999 7225 33011 7228
rect 32953 7219 33011 7225
rect 33410 7216 33416 7228
rect 33468 7256 33474 7268
rect 34517 7259 34575 7265
rect 34517 7256 34529 7259
rect 33468 7228 34529 7256
rect 33468 7216 33474 7228
rect 34517 7225 34529 7228
rect 34563 7225 34575 7259
rect 34517 7219 34575 7225
rect 35618 7216 35624 7268
rect 35676 7256 35682 7268
rect 38197 7259 38255 7265
rect 38197 7256 38209 7259
rect 35676 7228 38209 7256
rect 35676 7216 35682 7228
rect 38197 7225 38209 7228
rect 38243 7225 38255 7259
rect 38197 7219 38255 7225
rect 30834 7188 30840 7200
rect 29052 7160 30144 7188
rect 30747 7160 30840 7188
rect 29052 7148 29058 7160
rect 30834 7148 30840 7160
rect 30892 7188 30898 7200
rect 32048 7188 32076 7216
rect 30892 7160 32076 7188
rect 30892 7148 30898 7160
rect 32674 7148 32680 7200
rect 32732 7188 32738 7200
rect 33965 7191 34023 7197
rect 33965 7188 33977 7191
rect 32732 7160 33977 7188
rect 32732 7148 32738 7160
rect 33965 7157 33977 7160
rect 34011 7157 34023 7191
rect 35710 7188 35716 7200
rect 35671 7160 35716 7188
rect 33965 7151 34023 7157
rect 35710 7148 35716 7160
rect 35768 7148 35774 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 14274 6984 14280 6996
rect 13035 6956 14280 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 15010 6944 15016 6996
rect 15068 6984 15074 6996
rect 26234 6984 26240 6996
rect 15068 6956 26240 6984
rect 15068 6944 15074 6956
rect 26234 6944 26240 6956
rect 26292 6944 26298 6996
rect 28994 6984 29000 6996
rect 26344 6956 29000 6984
rect 12802 6876 12808 6928
rect 12860 6916 12866 6928
rect 12860 6888 19380 6916
rect 12860 6876 12866 6888
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6848 12403 6851
rect 15654 6848 15660 6860
rect 12391 6820 15660 6848
rect 12391 6817 12403 6820
rect 12345 6811 12403 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 16206 6848 16212 6860
rect 15887 6820 16212 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6848 16543 6851
rect 16850 6848 16856 6860
rect 16531 6820 16856 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6848 17831 6851
rect 17954 6848 17960 6860
rect 17819 6820 17960 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18598 6808 18604 6860
rect 18656 6848 18662 6860
rect 19242 6848 19248 6860
rect 18656 6820 19248 6848
rect 18656 6808 18662 6820
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 12250 6780 12256 6792
rect 12211 6752 12256 6780
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13354 6780 13360 6792
rect 12943 6752 13360 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13814 6780 13820 6792
rect 13587 6752 13820 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 13814 6740 13820 6752
rect 13872 6780 13878 6792
rect 14182 6780 14188 6792
rect 13872 6752 14188 6780
rect 13872 6740 13878 6752
rect 14182 6740 14188 6752
rect 14240 6780 14246 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14240 6752 14473 6780
rect 14240 6740 14246 6752
rect 14461 6749 14473 6752
rect 14507 6780 14519 6783
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 14507 6752 15117 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6780 15255 6783
rect 15378 6780 15384 6792
rect 15243 6752 15384 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6780 15807 6783
rect 16114 6780 16120 6792
rect 15795 6752 16120 6780
rect 15795 6749 15807 6752
rect 15749 6743 15807 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6780 16635 6783
rect 16942 6780 16948 6792
rect 16623 6752 16948 6780
rect 16623 6749 16635 6752
rect 16577 6743 16635 6749
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17218 6780 17224 6792
rect 17179 6752 17224 6780
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 18104 6752 18337 6780
rect 18104 6740 18110 6752
rect 18325 6749 18337 6752
rect 18371 6780 18383 6783
rect 18966 6780 18972 6792
rect 18371 6752 18972 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19352 6780 19380 6888
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 21177 6919 21235 6925
rect 21177 6916 21189 6919
rect 20772 6888 21189 6916
rect 20772 6876 20778 6888
rect 21177 6885 21189 6888
rect 21223 6916 21235 6919
rect 23382 6916 23388 6928
rect 21223 6888 21772 6916
rect 23343 6888 23388 6916
rect 21223 6885 21235 6888
rect 21177 6879 21235 6885
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 20898 6848 20904 6860
rect 19475 6820 20904 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 20898 6808 20904 6820
rect 20956 6848 20962 6860
rect 21358 6848 21364 6860
rect 20956 6820 21364 6848
rect 20956 6808 20962 6820
rect 21358 6808 21364 6820
rect 21416 6848 21422 6860
rect 21637 6851 21695 6857
rect 21637 6848 21649 6851
rect 21416 6820 21649 6848
rect 21416 6808 21422 6820
rect 21637 6817 21649 6820
rect 21683 6817 21695 6851
rect 21744 6848 21772 6888
rect 23382 6876 23388 6888
rect 23440 6876 23446 6928
rect 23658 6876 23664 6928
rect 23716 6916 23722 6928
rect 26344 6916 26372 6956
rect 28994 6944 29000 6956
rect 29052 6944 29058 6996
rect 29086 6944 29092 6996
rect 29144 6984 29150 6996
rect 29990 6987 30048 6993
rect 29990 6984 30002 6987
rect 29144 6956 30002 6984
rect 29144 6944 29150 6956
rect 29990 6953 30002 6956
rect 30036 6953 30048 6987
rect 31478 6984 31484 6996
rect 31439 6956 31484 6984
rect 29990 6947 30048 6953
rect 31478 6944 31484 6956
rect 31536 6944 31542 6996
rect 32030 6984 32036 6996
rect 31991 6956 32036 6984
rect 32030 6944 32036 6956
rect 32088 6944 32094 6996
rect 36078 6944 36084 6996
rect 36136 6984 36142 6996
rect 37093 6987 37151 6993
rect 37093 6984 37105 6987
rect 36136 6956 37105 6984
rect 36136 6944 36142 6956
rect 37093 6953 37105 6956
rect 37139 6984 37151 6987
rect 37645 6987 37703 6993
rect 37645 6984 37657 6987
rect 37139 6956 37657 6984
rect 37139 6953 37151 6956
rect 37093 6947 37151 6953
rect 37645 6953 37657 6956
rect 37691 6984 37703 6987
rect 37826 6984 37832 6996
rect 37691 6956 37832 6984
rect 37691 6953 37703 6956
rect 37645 6947 37703 6953
rect 37826 6944 37832 6956
rect 37884 6944 37890 6996
rect 38194 6984 38200 6996
rect 38155 6956 38200 6984
rect 38194 6944 38200 6956
rect 38252 6944 38258 6996
rect 23716 6888 26372 6916
rect 23716 6876 23722 6888
rect 24946 6848 24952 6860
rect 21744 6820 24952 6848
rect 21637 6811 21695 6817
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 25498 6848 25504 6860
rect 25459 6820 25504 6848
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 24026 6780 24032 6792
rect 19352 6752 19472 6780
rect 23939 6752 24032 6780
rect 13630 6712 13636 6724
rect 13591 6684 13636 6712
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 14553 6715 14611 6721
rect 14553 6681 14565 6715
rect 14599 6712 14611 6715
rect 17034 6712 17040 6724
rect 14599 6684 17040 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 17034 6672 17040 6684
rect 17092 6672 17098 6724
rect 17129 6715 17187 6721
rect 17129 6681 17141 6715
rect 17175 6712 17187 6715
rect 19334 6712 19340 6724
rect 17175 6684 19340 6712
rect 17175 6681 17187 6684
rect 17129 6675 17187 6681
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 18506 6644 18512 6656
rect 18467 6616 18512 6644
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 19444 6644 19472 6752
rect 24026 6740 24032 6752
rect 24084 6780 24090 6792
rect 24765 6783 24823 6789
rect 24765 6780 24777 6783
rect 24084 6752 24777 6780
rect 24084 6740 24090 6752
rect 24765 6749 24777 6752
rect 24811 6780 24823 6783
rect 24811 6752 24900 6780
rect 24811 6749 24823 6752
rect 24765 6743 24823 6749
rect 19705 6715 19763 6721
rect 19705 6681 19717 6715
rect 19751 6712 19763 6715
rect 19794 6712 19800 6724
rect 19751 6684 19800 6712
rect 19751 6681 19763 6684
rect 19705 6675 19763 6681
rect 19794 6672 19800 6684
rect 19852 6672 19858 6724
rect 21542 6712 21548 6724
rect 20930 6684 21548 6712
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 21634 6672 21640 6724
rect 21692 6712 21698 6724
rect 21913 6715 21971 6721
rect 21913 6712 21925 6715
rect 21692 6684 21925 6712
rect 21692 6672 21698 6684
rect 21913 6681 21925 6684
rect 21959 6681 21971 6715
rect 23934 6712 23940 6724
rect 21913 6675 21971 6681
rect 22020 6684 22402 6712
rect 23895 6684 23940 6712
rect 20714 6644 20720 6656
rect 19444 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 20990 6604 20996 6656
rect 21048 6644 21054 6656
rect 22020 6644 22048 6684
rect 23934 6672 23940 6684
rect 23992 6672 23998 6724
rect 24872 6712 24900 6752
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25409 6783 25467 6789
rect 25409 6780 25421 6783
rect 25188 6752 25421 6780
rect 25188 6740 25194 6752
rect 25409 6749 25421 6752
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 26050 6712 26056 6724
rect 24872 6684 26056 6712
rect 26050 6672 26056 6684
rect 26108 6672 26114 6724
rect 26160 6712 26188 6888
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26602 6848 26608 6860
rect 26283 6820 26608 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 27154 6808 27160 6860
rect 27212 6848 27218 6860
rect 27212 6820 28764 6848
rect 27212 6808 27218 6820
rect 28736 6789 28764 6820
rect 31570 6808 31576 6860
rect 31628 6848 31634 6860
rect 32493 6851 32551 6857
rect 32493 6848 32505 6851
rect 31628 6820 32505 6848
rect 31628 6808 31634 6820
rect 32493 6817 32505 6820
rect 32539 6817 32551 6851
rect 32493 6811 32551 6817
rect 34606 6808 34612 6860
rect 34664 6848 34670 6860
rect 35434 6848 35440 6860
rect 34664 6820 35440 6848
rect 34664 6808 34670 6820
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 28721 6783 28779 6789
rect 28721 6749 28733 6783
rect 28767 6749 28779 6783
rect 29730 6780 29736 6792
rect 29691 6752 29736 6780
rect 28721 6743 28779 6749
rect 26513 6715 26571 6721
rect 26513 6712 26525 6715
rect 26160 6684 26525 6712
rect 26513 6681 26525 6684
rect 26559 6681 26571 6715
rect 28629 6715 28687 6721
rect 28629 6712 28641 6715
rect 27738 6684 28641 6712
rect 26513 6675 26571 6681
rect 28629 6681 28641 6684
rect 28675 6681 28687 6715
rect 28736 6712 28764 6743
rect 29730 6740 29736 6752
rect 29788 6740 29794 6792
rect 30282 6712 30288 6724
rect 28736 6684 30288 6712
rect 28629 6675 28687 6681
rect 30282 6672 30288 6684
rect 30340 6672 30346 6724
rect 30466 6672 30472 6724
rect 30524 6672 30530 6724
rect 34149 6715 34207 6721
rect 34149 6712 34161 6715
rect 33612 6684 34161 6712
rect 21048 6616 22048 6644
rect 21048 6604 21054 6616
rect 24486 6604 24492 6656
rect 24544 6644 24550 6656
rect 24673 6647 24731 6653
rect 24673 6644 24685 6647
rect 24544 6616 24685 6644
rect 24544 6604 24550 6616
rect 24673 6613 24685 6616
rect 24719 6613 24731 6647
rect 27982 6644 27988 6656
rect 27943 6616 27988 6644
rect 24673 6607 24731 6613
rect 27982 6604 27988 6616
rect 28040 6604 28046 6656
rect 30300 6644 30328 6672
rect 32490 6644 32496 6656
rect 30300 6616 32496 6644
rect 32490 6604 32496 6616
rect 32548 6644 32554 6656
rect 33137 6647 33195 6653
rect 33137 6644 33149 6647
rect 32548 6616 33149 6644
rect 32548 6604 32554 6616
rect 33137 6613 33149 6616
rect 33183 6613 33195 6647
rect 33137 6607 33195 6613
rect 33410 6604 33416 6656
rect 33468 6644 33474 6656
rect 33612 6653 33640 6684
rect 34149 6681 34161 6684
rect 34195 6681 34207 6715
rect 34149 6675 34207 6681
rect 33597 6647 33655 6653
rect 33597 6644 33609 6647
rect 33468 6616 33609 6644
rect 33468 6604 33474 6616
rect 33597 6613 33609 6616
rect 33643 6613 33655 6647
rect 33597 6607 33655 6613
rect 33686 6604 33692 6656
rect 33744 6644 33750 6656
rect 34885 6647 34943 6653
rect 34885 6644 34897 6647
rect 33744 6616 34897 6644
rect 33744 6604 33750 6616
rect 34885 6613 34897 6616
rect 34931 6613 34943 6647
rect 34885 6607 34943 6613
rect 35802 6604 35808 6656
rect 35860 6644 35866 6656
rect 35989 6647 36047 6653
rect 35989 6644 36001 6647
rect 35860 6616 36001 6644
rect 35860 6604 35866 6616
rect 35989 6613 36001 6616
rect 36035 6613 36047 6647
rect 36630 6644 36636 6656
rect 36591 6616 36636 6644
rect 35989 6607 36047 6613
rect 36630 6604 36636 6616
rect 36688 6604 36694 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 12526 6440 12532 6452
rect 12483 6412 12532 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 13081 6443 13139 6449
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 13446 6440 13452 6452
rect 13127 6412 13452 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 13906 6440 13912 6452
rect 13771 6412 13912 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 15013 6443 15071 6449
rect 15013 6409 15025 6443
rect 15059 6440 15071 6443
rect 16574 6440 16580 6452
rect 15059 6412 16580 6440
rect 15059 6409 15071 6412
rect 15013 6403 15071 6409
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 19334 6440 19340 6452
rect 17000 6412 19340 6440
rect 17000 6400 17006 6412
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20257 6443 20315 6449
rect 20257 6440 20269 6443
rect 20036 6412 20269 6440
rect 20036 6400 20042 6412
rect 20257 6409 20269 6412
rect 20303 6409 20315 6443
rect 20257 6403 20315 6409
rect 22278 6400 22284 6452
rect 22336 6440 22342 6452
rect 22336 6412 26004 6440
rect 22336 6400 22342 6412
rect 15746 6332 15752 6384
rect 15804 6372 15810 6384
rect 18322 6372 18328 6384
rect 15804 6344 15849 6372
rect 18283 6344 18328 6372
rect 15804 6332 15810 6344
rect 18322 6332 18328 6344
rect 18380 6332 18386 6384
rect 18414 6332 18420 6384
rect 18472 6372 18478 6384
rect 19521 6375 19579 6381
rect 19521 6372 19533 6375
rect 18472 6344 19533 6372
rect 18472 6332 18478 6344
rect 19521 6341 19533 6344
rect 19567 6341 19579 6375
rect 19521 6335 19579 6341
rect 19613 6375 19671 6381
rect 19613 6341 19625 6375
rect 19659 6372 19671 6375
rect 20070 6372 20076 6384
rect 19659 6344 20076 6372
rect 19659 6341 19671 6344
rect 19613 6335 19671 6341
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 22094 6372 22100 6384
rect 20180 6344 22100 6372
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6273 12587 6307
rect 13170 6304 13176 6316
rect 13131 6276 13176 6304
rect 12529 6267 12587 6273
rect 12544 6236 12572 6267
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13633 6307 13691 6313
rect 13633 6304 13645 6307
rect 13412 6276 13645 6304
rect 13412 6264 13418 6276
rect 13633 6273 13645 6276
rect 13679 6304 13691 6307
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13679 6276 14289 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 14277 6273 14289 6276
rect 14323 6304 14335 6307
rect 14458 6304 14464 6316
rect 14323 6276 14464 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 14458 6264 14464 6276
rect 14516 6304 14522 6316
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14516 6276 14933 6304
rect 14516 6264 14522 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16356 6276 16401 6304
rect 16356 6264 16362 6276
rect 13372 6236 13400 6264
rect 12544 6208 13400 6236
rect 15378 6196 15384 6248
rect 15436 6236 15442 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15436 6208 15669 6236
rect 15436 6196 15442 6208
rect 15657 6205 15669 6208
rect 15703 6236 15715 6239
rect 16666 6236 16672 6248
rect 15703 6208 16672 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 17678 6236 17684 6248
rect 17359 6208 17684 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6236 18475 6239
rect 19426 6236 19432 6248
rect 18463 6208 19432 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 14369 6171 14427 6177
rect 14369 6137 14381 6171
rect 14415 6168 14427 6171
rect 16022 6168 16028 6180
rect 14415 6140 16028 6168
rect 14415 6137 14427 6140
rect 14369 6131 14427 6137
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 17865 6171 17923 6177
rect 17865 6168 17877 6171
rect 16500 6140 17877 6168
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 16500 6100 16528 6140
rect 17865 6137 17877 6140
rect 17911 6168 17923 6171
rect 18782 6168 18788 6180
rect 17911 6140 18788 6168
rect 17911 6137 17923 6140
rect 17865 6131 17923 6137
rect 18782 6128 18788 6140
rect 18840 6168 18846 6180
rect 19061 6171 19119 6177
rect 19061 6168 19073 6171
rect 18840 6140 19073 6168
rect 18840 6128 18846 6140
rect 19061 6137 19073 6140
rect 19107 6137 19119 6171
rect 19061 6131 19119 6137
rect 14332 6072 16528 6100
rect 14332 6060 14338 6072
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 20180 6100 20208 6344
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 23658 6332 23664 6384
rect 23716 6372 23722 6384
rect 23716 6344 24808 6372
rect 23716 6332 23722 6344
rect 20346 6304 20352 6316
rect 20307 6276 20352 6304
rect 20346 6264 20352 6276
rect 20404 6264 20410 6316
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 20496 6276 22494 6304
rect 20496 6264 20502 6276
rect 23842 6264 23848 6316
rect 23900 6304 23906 6316
rect 24670 6304 24676 6316
rect 23900 6276 23945 6304
rect 24136 6276 24676 6304
rect 23900 6264 23906 6276
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 22097 6239 22155 6245
rect 22097 6236 22109 6239
rect 20864 6208 22109 6236
rect 20864 6196 20870 6208
rect 22097 6205 22109 6208
rect 22143 6236 22155 6239
rect 23014 6236 23020 6248
rect 22143 6208 23020 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 23474 6196 23480 6248
rect 23532 6236 23538 6248
rect 23569 6239 23627 6245
rect 23569 6236 23581 6239
rect 23532 6208 23581 6236
rect 23532 6196 23538 6208
rect 23569 6205 23581 6208
rect 23615 6236 23627 6239
rect 24136 6236 24164 6276
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 24578 6236 24584 6248
rect 23615 6208 24164 6236
rect 24539 6208 24584 6236
rect 23615 6205 23627 6208
rect 23569 6199 23627 6205
rect 24578 6196 24584 6208
rect 24636 6196 24642 6248
rect 24780 6236 24808 6344
rect 24854 6332 24860 6384
rect 24912 6372 24918 6384
rect 25976 6372 26004 6412
rect 26050 6400 26056 6452
rect 26108 6440 26114 6452
rect 26510 6440 26516 6452
rect 26108 6412 26516 6440
rect 26108 6400 26114 6412
rect 26510 6400 26516 6412
rect 26568 6400 26574 6452
rect 27246 6440 27252 6452
rect 27207 6412 27252 6440
rect 27246 6400 27252 6412
rect 27304 6400 27310 6452
rect 27985 6443 28043 6449
rect 27985 6409 27997 6443
rect 28031 6440 28043 6443
rect 28442 6440 28448 6452
rect 28031 6412 28448 6440
rect 28031 6409 28043 6412
rect 27985 6403 28043 6409
rect 28442 6400 28448 6412
rect 28500 6400 28506 6452
rect 28810 6400 28816 6452
rect 28868 6440 28874 6452
rect 28868 6412 31754 6440
rect 28868 6400 28874 6412
rect 24912 6344 25162 6372
rect 25976 6344 28290 6372
rect 24912 6332 24918 6344
rect 29362 6332 29368 6384
rect 29420 6372 29426 6384
rect 29457 6375 29515 6381
rect 29457 6372 29469 6375
rect 29420 6344 29469 6372
rect 29420 6332 29426 6344
rect 29457 6341 29469 6344
rect 29503 6372 29515 6375
rect 29822 6372 29828 6384
rect 29503 6344 29828 6372
rect 29503 6341 29515 6344
rect 29457 6335 29515 6341
rect 29822 6332 29828 6344
rect 29880 6332 29886 6384
rect 30006 6332 30012 6384
rect 30064 6372 30070 6384
rect 31570 6372 31576 6384
rect 30064 6344 31576 6372
rect 30064 6332 30070 6344
rect 31570 6332 31576 6344
rect 31628 6332 31634 6384
rect 31726 6372 31754 6412
rect 33594 6400 33600 6452
rect 33652 6440 33658 6452
rect 33965 6443 34023 6449
rect 33965 6440 33977 6443
rect 33652 6412 33977 6440
rect 33652 6400 33658 6412
rect 33965 6409 33977 6412
rect 34011 6409 34023 6443
rect 33965 6403 34023 6409
rect 35989 6375 36047 6381
rect 35989 6372 36001 6375
rect 31726 6344 36001 6372
rect 35989 6341 36001 6344
rect 36035 6341 36047 6375
rect 38010 6372 38016 6384
rect 37971 6344 38016 6372
rect 35989 6335 36047 6341
rect 38010 6332 38016 6344
rect 38068 6332 38074 6384
rect 27157 6307 27215 6313
rect 27157 6273 27169 6307
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 26234 6236 26240 6248
rect 24780 6208 26240 6236
rect 26234 6196 26240 6208
rect 26292 6236 26298 6248
rect 26329 6239 26387 6245
rect 26329 6236 26341 6239
rect 26292 6208 26341 6236
rect 26292 6196 26298 6208
rect 26329 6205 26341 6208
rect 26375 6205 26387 6239
rect 26602 6236 26608 6248
rect 26563 6208 26608 6236
rect 26329 6199 26387 6205
rect 26602 6196 26608 6208
rect 26660 6196 26666 6248
rect 23934 6128 23940 6180
rect 23992 6168 23998 6180
rect 23992 6140 24992 6168
rect 23992 6128 23998 6140
rect 20898 6100 20904 6112
rect 16908 6072 20208 6100
rect 20859 6072 20904 6100
rect 16908 6060 16914 6072
rect 20898 6060 20904 6072
rect 20956 6100 20962 6112
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 20956 6072 21373 6100
rect 20956 6060 20962 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 21361 6063 21419 6069
rect 21726 6060 21732 6112
rect 21784 6100 21790 6112
rect 24854 6100 24860 6112
rect 21784 6072 24860 6100
rect 21784 6060 21790 6072
rect 24854 6060 24860 6072
rect 24912 6060 24918 6112
rect 24964 6100 24992 6140
rect 27172 6100 27200 6267
rect 30282 6264 30288 6316
rect 30340 6304 30346 6316
rect 30377 6307 30435 6313
rect 30377 6304 30389 6307
rect 30340 6276 30389 6304
rect 30340 6264 30346 6276
rect 30377 6273 30389 6276
rect 30423 6273 30435 6307
rect 30377 6267 30435 6273
rect 30558 6264 30564 6316
rect 30616 6304 30622 6316
rect 34054 6304 34060 6316
rect 30616 6276 34060 6304
rect 30616 6264 30622 6276
rect 34054 6264 34060 6276
rect 34112 6264 34118 6316
rect 35434 6304 35440 6316
rect 35395 6276 35440 6304
rect 35434 6264 35440 6276
rect 35492 6304 35498 6316
rect 36081 6307 36139 6313
rect 36081 6304 36093 6307
rect 35492 6276 36093 6304
rect 35492 6264 35498 6276
rect 36081 6273 36093 6276
rect 36127 6304 36139 6307
rect 36541 6307 36599 6313
rect 36541 6304 36553 6307
rect 36127 6276 36553 6304
rect 36127 6273 36139 6276
rect 36081 6267 36139 6273
rect 36541 6273 36553 6276
rect 36587 6273 36599 6307
rect 36541 6267 36599 6273
rect 37553 6307 37611 6313
rect 37553 6273 37565 6307
rect 37599 6304 37611 6307
rect 38194 6304 38200 6316
rect 37599 6276 38200 6304
rect 37599 6273 37611 6276
rect 37553 6267 37611 6273
rect 38194 6264 38200 6276
rect 38252 6264 38258 6316
rect 29730 6236 29736 6248
rect 29691 6208 29736 6236
rect 29730 6196 29736 6208
rect 29788 6196 29794 6248
rect 30929 6239 30987 6245
rect 30929 6205 30941 6239
rect 30975 6236 30987 6239
rect 31938 6236 31944 6248
rect 30975 6208 31944 6236
rect 30975 6205 30987 6208
rect 30929 6199 30987 6205
rect 31938 6196 31944 6208
rect 31996 6236 32002 6248
rect 32401 6239 32459 6245
rect 32401 6236 32413 6239
rect 31996 6208 32413 6236
rect 31996 6196 32002 6208
rect 32401 6205 32413 6208
rect 32447 6236 32459 6239
rect 32953 6239 33011 6245
rect 32953 6236 32965 6239
rect 32447 6208 32965 6236
rect 32447 6205 32459 6208
rect 32401 6199 32459 6205
rect 32953 6205 32965 6208
rect 32999 6236 33011 6239
rect 32999 6208 33456 6236
rect 32999 6205 33011 6208
rect 32953 6199 33011 6205
rect 33428 6180 33456 6208
rect 31570 6128 31576 6180
rect 31628 6168 31634 6180
rect 33134 6168 33140 6180
rect 31628 6140 33140 6168
rect 31628 6128 31634 6140
rect 33134 6128 33140 6140
rect 33192 6128 33198 6180
rect 33410 6168 33416 6180
rect 33371 6140 33416 6168
rect 33410 6128 33416 6140
rect 33468 6128 33474 6180
rect 24964 6072 27200 6100
rect 29270 6060 29276 6112
rect 29328 6100 29334 6112
rect 30285 6103 30343 6109
rect 30285 6100 30297 6103
rect 29328 6072 30297 6100
rect 29328 6060 29334 6072
rect 30285 6069 30297 6072
rect 30331 6069 30343 6103
rect 30285 6063 30343 6069
rect 30374 6060 30380 6112
rect 30432 6100 30438 6112
rect 31389 6103 31447 6109
rect 31389 6100 31401 6103
rect 30432 6072 31401 6100
rect 30432 6060 30438 6072
rect 31389 6069 31401 6072
rect 31435 6069 31447 6103
rect 31389 6063 31447 6069
rect 32490 6060 32496 6112
rect 32548 6100 32554 6112
rect 34514 6100 34520 6112
rect 32548 6072 34520 6100
rect 32548 6060 32554 6072
rect 34514 6060 34520 6072
rect 34572 6060 34578 6112
rect 35342 6100 35348 6112
rect 35303 6072 35348 6100
rect 35342 6060 35348 6072
rect 35400 6060 35406 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 13262 5896 13268 5908
rect 12299 5868 13268 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 12268 5692 12296 5859
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 13633 5899 13691 5905
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 13722 5896 13728 5908
rect 13679 5868 13728 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 15378 5896 15384 5908
rect 14415 5868 15384 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 15562 5896 15568 5908
rect 15523 5868 15568 5896
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 16850 5896 16856 5908
rect 16080 5868 16856 5896
rect 16080 5856 16086 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 20162 5896 20168 5908
rect 17083 5868 20168 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20404 5868 23980 5896
rect 20404 5856 20410 5868
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 15930 5828 15936 5840
rect 14792 5800 15936 5828
rect 14792 5788 14798 5800
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 16666 5788 16672 5840
rect 16724 5828 16730 5840
rect 17586 5828 17592 5840
rect 16724 5800 17592 5828
rect 16724 5788 16730 5800
rect 17586 5788 17592 5800
rect 17644 5788 17650 5840
rect 17678 5788 17684 5840
rect 17736 5828 17742 5840
rect 17736 5800 18092 5828
rect 17736 5788 17742 5800
rect 17954 5760 17960 5772
rect 15672 5732 17960 5760
rect 11747 5664 12296 5692
rect 13541 5695 13599 5701
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13630 5692 13636 5704
rect 13587 5664 13636 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 15672 5701 15700 5732
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18064 5760 18092 5800
rect 18138 5788 18144 5840
rect 18196 5828 18202 5840
rect 20622 5828 20628 5840
rect 18196 5800 20628 5828
rect 18196 5788 18202 5800
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 20806 5828 20812 5840
rect 20767 5800 20812 5828
rect 20806 5788 20812 5800
rect 20864 5788 20870 5840
rect 20990 5788 20996 5840
rect 21048 5828 21054 5840
rect 21358 5828 21364 5840
rect 21048 5800 21364 5828
rect 21048 5788 21054 5800
rect 21358 5788 21364 5800
rect 21416 5788 21422 5840
rect 23952 5828 23980 5868
rect 24026 5856 24032 5908
rect 24084 5896 24090 5908
rect 31570 5896 31576 5908
rect 24084 5868 31576 5896
rect 24084 5856 24090 5868
rect 31570 5856 31576 5868
rect 31628 5856 31634 5908
rect 31662 5856 31668 5908
rect 31720 5896 31726 5908
rect 33689 5899 33747 5905
rect 33689 5896 33701 5899
rect 31720 5868 33701 5896
rect 31720 5856 31726 5868
rect 33689 5865 33701 5868
rect 33735 5865 33747 5899
rect 35618 5896 35624 5908
rect 33689 5859 33747 5865
rect 33980 5868 35624 5896
rect 24394 5828 24400 5840
rect 23952 5800 24400 5828
rect 24394 5788 24400 5800
rect 24452 5788 24458 5840
rect 26326 5828 26332 5840
rect 26287 5800 26332 5828
rect 26326 5788 26332 5800
rect 26384 5788 26390 5840
rect 28902 5828 28908 5840
rect 28863 5800 28908 5828
rect 28902 5788 28908 5800
rect 28960 5788 28966 5840
rect 31386 5788 31392 5840
rect 31444 5828 31450 5840
rect 31481 5831 31539 5837
rect 31481 5828 31493 5831
rect 31444 5800 31493 5828
rect 31444 5788 31450 5800
rect 31481 5797 31493 5800
rect 31527 5828 31539 5831
rect 31527 5800 31754 5828
rect 31527 5797 31539 5800
rect 31481 5791 31539 5797
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 18064 5732 18245 5760
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 23658 5760 23664 5772
rect 19208 5732 23664 5760
rect 19208 5720 19214 5732
rect 23658 5720 23664 5732
rect 23716 5720 23722 5772
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 24581 5763 24639 5769
rect 24581 5760 24593 5763
rect 23900 5732 24593 5760
rect 23900 5720 23906 5732
rect 24581 5729 24593 5732
rect 24627 5729 24639 5763
rect 24854 5760 24860 5772
rect 24815 5732 24860 5760
rect 24581 5723 24639 5729
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 24946 5720 24952 5772
rect 25004 5760 25010 5772
rect 27433 5763 27491 5769
rect 27433 5760 27445 5763
rect 25004 5732 27445 5760
rect 25004 5720 25010 5732
rect 27433 5729 27445 5732
rect 27479 5729 27491 5763
rect 29730 5760 29736 5772
rect 29691 5732 29736 5760
rect 27433 5723 27491 5729
rect 29730 5720 29736 5732
rect 29788 5720 29794 5772
rect 30006 5760 30012 5772
rect 29919 5732 30012 5760
rect 30006 5720 30012 5732
rect 30064 5760 30070 5772
rect 31018 5760 31024 5772
rect 30064 5732 31024 5760
rect 30064 5720 30070 5732
rect 31018 5720 31024 5732
rect 31076 5720 31082 5772
rect 14829 5695 14887 5701
rect 14829 5692 14841 5695
rect 14516 5664 14841 5692
rect 14516 5652 14522 5664
rect 14829 5661 14841 5664
rect 14875 5692 14887 5695
rect 15657 5695 15715 5701
rect 14875 5664 15240 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15212 5624 15240 5664
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 16114 5692 16120 5704
rect 15657 5655 15715 5661
rect 15764 5664 16120 5692
rect 15764 5624 15792 5664
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16937 5697 16995 5703
rect 16937 5694 16949 5697
rect 16868 5666 16949 5694
rect 16206 5624 16212 5636
rect 15212 5596 15792 5624
rect 16167 5596 16212 5624
rect 16206 5584 16212 5596
rect 16264 5584 16270 5636
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 16868 5624 16896 5666
rect 16937 5663 16949 5666
rect 16983 5663 16995 5697
rect 16937 5657 16995 5663
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 21361 5695 21419 5701
rect 18932 5664 18977 5692
rect 18932 5652 18938 5664
rect 21361 5661 21373 5695
rect 21407 5661 21419 5695
rect 24026 5692 24032 5704
rect 23987 5664 24032 5692
rect 21361 5655 21419 5661
rect 16632 5596 16896 5624
rect 18318 5627 18376 5633
rect 16632 5584 16638 5596
rect 18318 5593 18330 5627
rect 18364 5624 18376 5627
rect 19150 5624 19156 5636
rect 18364 5596 19156 5624
rect 18364 5593 18376 5596
rect 18318 5587 18376 5593
rect 19150 5584 19156 5596
rect 19208 5584 19214 5636
rect 19797 5627 19855 5633
rect 19797 5593 19809 5627
rect 19843 5624 19855 5627
rect 20257 5627 20315 5633
rect 20257 5624 20269 5627
rect 19843 5596 20269 5624
rect 19843 5593 19855 5596
rect 19797 5587 19855 5593
rect 20257 5593 20269 5596
rect 20303 5624 20315 5627
rect 20898 5624 20904 5636
rect 20303 5596 20904 5624
rect 20303 5593 20315 5596
rect 20257 5587 20315 5593
rect 20898 5584 20904 5596
rect 20956 5624 20962 5636
rect 21266 5624 21272 5636
rect 20956 5596 21272 5624
rect 20956 5584 20962 5596
rect 21266 5584 21272 5596
rect 21324 5624 21330 5636
rect 21376 5624 21404 5655
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 26326 5652 26332 5704
rect 26384 5692 26390 5704
rect 26602 5692 26608 5704
rect 26384 5664 26608 5692
rect 26384 5652 26390 5664
rect 26602 5652 26608 5664
rect 26660 5692 26666 5704
rect 27157 5695 27215 5701
rect 27157 5692 27169 5695
rect 26660 5664 27169 5692
rect 26660 5652 26666 5664
rect 27157 5661 27169 5664
rect 27203 5661 27215 5695
rect 27157 5655 27215 5661
rect 21324 5596 21404 5624
rect 21324 5584 21330 5596
rect 21542 5584 21548 5636
rect 21600 5624 21606 5636
rect 21637 5627 21695 5633
rect 21637 5624 21649 5627
rect 21600 5596 21649 5624
rect 21600 5584 21606 5596
rect 21637 5593 21649 5596
rect 21683 5624 21695 5627
rect 21910 5624 21916 5636
rect 21683 5596 21916 5624
rect 21683 5593 21695 5596
rect 21637 5587 21695 5593
rect 21910 5584 21916 5596
rect 21968 5584 21974 5636
rect 22370 5584 22376 5636
rect 22428 5584 22434 5636
rect 23198 5584 23204 5636
rect 23256 5624 23262 5636
rect 23385 5627 23443 5633
rect 23385 5624 23397 5627
rect 23256 5596 23397 5624
rect 23256 5584 23262 5596
rect 23385 5593 23397 5596
rect 23431 5593 23443 5627
rect 23385 5587 23443 5593
rect 25314 5584 25320 5636
rect 25372 5584 25378 5636
rect 28718 5624 28724 5636
rect 28658 5596 28724 5624
rect 28718 5584 28724 5596
rect 28776 5584 28782 5636
rect 31726 5624 31754 5800
rect 31938 5760 31944 5772
rect 31899 5732 31944 5760
rect 31938 5720 31944 5732
rect 31996 5720 32002 5772
rect 33980 5692 34008 5868
rect 35618 5856 35624 5868
rect 35676 5856 35682 5908
rect 37090 5896 37096 5908
rect 37051 5868 37096 5896
rect 37090 5856 37096 5868
rect 37148 5856 37154 5908
rect 38102 5856 38108 5908
rect 38160 5896 38166 5908
rect 38197 5899 38255 5905
rect 38197 5896 38209 5899
rect 38160 5868 38209 5896
rect 38160 5856 38166 5868
rect 38197 5865 38209 5868
rect 38243 5865 38255 5899
rect 38197 5859 38255 5865
rect 34514 5788 34520 5840
rect 34572 5828 34578 5840
rect 35802 5828 35808 5840
rect 34572 5800 35808 5828
rect 34572 5788 34578 5800
rect 35802 5788 35808 5800
rect 35860 5828 35866 5840
rect 35989 5831 36047 5837
rect 35989 5828 36001 5831
rect 35860 5800 36001 5828
rect 35860 5788 35866 5800
rect 35989 5797 36001 5800
rect 36035 5828 36047 5831
rect 37645 5831 37703 5837
rect 37645 5828 37657 5831
rect 36035 5800 37657 5828
rect 36035 5797 36047 5800
rect 35989 5791 36047 5797
rect 37645 5797 37657 5800
rect 37691 5797 37703 5831
rect 37645 5791 37703 5797
rect 34054 5720 34060 5772
rect 34112 5760 34118 5772
rect 35437 5763 35495 5769
rect 35437 5760 35449 5763
rect 34112 5732 35449 5760
rect 34112 5720 34118 5732
rect 35437 5729 35449 5732
rect 35483 5729 35495 5763
rect 35437 5723 35495 5729
rect 33350 5664 34008 5692
rect 32217 5627 32275 5633
rect 32217 5624 32229 5627
rect 31234 5596 31616 5624
rect 31726 5596 32229 5624
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 9272 5528 11529 5556
rect 9272 5516 9278 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 14918 5556 14924 5568
rect 14879 5528 14924 5556
rect 11517 5519 11575 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 18782 5516 18788 5568
rect 18840 5556 18846 5568
rect 20438 5556 20444 5568
rect 18840 5528 20444 5556
rect 18840 5516 18846 5528
rect 20438 5516 20444 5528
rect 20496 5516 20502 5568
rect 20530 5516 20536 5568
rect 20588 5556 20594 5568
rect 22646 5556 22652 5568
rect 20588 5528 22652 5556
rect 20588 5516 20594 5528
rect 22646 5516 22652 5528
rect 22704 5516 22710 5568
rect 23290 5516 23296 5568
rect 23348 5556 23354 5568
rect 23937 5559 23995 5565
rect 23937 5556 23949 5559
rect 23348 5528 23949 5556
rect 23348 5516 23354 5528
rect 23937 5525 23949 5528
rect 23983 5525 23995 5559
rect 23937 5519 23995 5525
rect 24394 5516 24400 5568
rect 24452 5556 24458 5568
rect 31018 5556 31024 5568
rect 24452 5528 31024 5556
rect 24452 5516 24458 5528
rect 31018 5516 31024 5528
rect 31076 5516 31082 5568
rect 31588 5556 31616 5596
rect 32217 5593 32229 5596
rect 32263 5593 32275 5627
rect 34698 5624 34704 5636
rect 32217 5587 32275 5593
rect 34164 5596 34704 5624
rect 34164 5556 34192 5596
rect 34698 5584 34704 5596
rect 34756 5584 34762 5636
rect 31588 5528 34192 5556
rect 34241 5559 34299 5565
rect 34241 5525 34253 5559
rect 34287 5556 34299 5559
rect 34790 5556 34796 5568
rect 34287 5528 34796 5556
rect 34287 5525 34299 5528
rect 34241 5519 34299 5525
rect 34790 5516 34796 5528
rect 34848 5556 34854 5568
rect 34885 5559 34943 5565
rect 34885 5556 34897 5559
rect 34848 5528 34897 5556
rect 34848 5516 34854 5528
rect 34885 5525 34897 5528
rect 34931 5556 34943 5559
rect 36541 5559 36599 5565
rect 36541 5556 36553 5559
rect 34931 5528 36553 5556
rect 34931 5525 34943 5528
rect 34885 5519 34943 5525
rect 36541 5525 36553 5528
rect 36587 5525 36599 5559
rect 36541 5519 36599 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 14090 5352 14096 5364
rect 14047 5324 14096 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 15197 5355 15255 5361
rect 15197 5321 15209 5355
rect 15243 5352 15255 5355
rect 15746 5352 15752 5364
rect 15243 5324 15752 5352
rect 15243 5321 15255 5324
rect 15197 5315 15255 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16942 5352 16948 5364
rect 16903 5324 16948 5352
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 23750 5352 23756 5364
rect 18196 5324 23612 5352
rect 23711 5324 23756 5352
rect 18196 5312 18202 5324
rect 13449 5287 13507 5293
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 16117 5287 16175 5293
rect 13495 5256 16068 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 16040 5228 16068 5256
rect 16117 5253 16129 5287
rect 16163 5284 16175 5287
rect 17126 5284 17132 5296
rect 16163 5256 17132 5284
rect 16163 5253 16175 5256
rect 16117 5247 16175 5253
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 18046 5244 18052 5296
rect 18104 5284 18110 5296
rect 18417 5287 18475 5293
rect 18417 5284 18429 5287
rect 18104 5256 18429 5284
rect 18104 5244 18110 5256
rect 18417 5253 18429 5256
rect 18463 5253 18475 5287
rect 18417 5247 18475 5253
rect 18509 5287 18567 5293
rect 18509 5253 18521 5287
rect 18555 5284 18567 5287
rect 18690 5284 18696 5296
rect 18555 5256 18696 5284
rect 18555 5253 18567 5256
rect 18509 5247 18567 5253
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 18966 5244 18972 5296
rect 19024 5284 19030 5296
rect 19061 5287 19119 5293
rect 19061 5284 19073 5287
rect 19024 5256 19073 5284
rect 19024 5244 19030 5256
rect 19061 5253 19073 5256
rect 19107 5253 19119 5287
rect 19061 5247 19119 5253
rect 20717 5287 20775 5293
rect 20717 5253 20729 5287
rect 20763 5284 20775 5287
rect 20806 5284 20812 5296
rect 20763 5256 20812 5284
rect 20763 5253 20775 5256
rect 20717 5247 20775 5253
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 20898 5244 20904 5296
rect 20956 5284 20962 5296
rect 23584 5284 23612 5324
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 23842 5312 23848 5364
rect 23900 5352 23906 5364
rect 24946 5352 24952 5364
rect 23900 5324 24952 5352
rect 23900 5312 23906 5324
rect 24946 5312 24952 5324
rect 25004 5312 25010 5364
rect 25038 5312 25044 5364
rect 25096 5352 25102 5364
rect 30006 5352 30012 5364
rect 25096 5324 29868 5352
rect 29967 5324 30012 5352
rect 25096 5312 25102 5324
rect 25792 5293 25820 5324
rect 25777 5287 25835 5293
rect 20956 5256 21312 5284
rect 23584 5256 24610 5284
rect 20956 5244 20962 5256
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 10318 5216 10324 5228
rect 1903 5188 10324 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12434 5216 12440 5228
rect 12299 5188 12440 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 14458 5216 14464 5228
rect 14419 5188 14464 5216
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5185 15347 5219
rect 16022 5216 16028 5228
rect 15983 5188 16028 5216
rect 15289 5179 15347 5185
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 15194 5148 15200 5160
rect 12391 5120 15200 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15304 5080 15332 5179
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 17034 5216 17040 5228
rect 16995 5188 17040 5216
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 19242 5176 19248 5228
rect 19300 5216 19306 5228
rect 20625 5219 20683 5225
rect 19300 5188 20576 5216
rect 19300 5176 19306 5188
rect 18230 5108 18236 5160
rect 18288 5148 18294 5160
rect 20438 5148 20444 5160
rect 18288 5120 20444 5148
rect 18288 5108 18294 5120
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 17678 5080 17684 5092
rect 15304 5052 17684 5080
rect 17678 5040 17684 5052
rect 17736 5040 17742 5092
rect 17954 5080 17960 5092
rect 17915 5052 17960 5080
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 18782 5040 18788 5092
rect 18840 5080 18846 5092
rect 19978 5080 19984 5092
rect 18840 5052 19984 5080
rect 18840 5040 18846 5052
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 20548 5080 20576 5188
rect 20625 5185 20637 5219
rect 20671 5216 20683 5219
rect 21174 5216 21180 5228
rect 20671 5188 21180 5216
rect 20671 5185 20683 5188
rect 20625 5179 20683 5185
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 21284 5225 21312 5256
rect 25777 5253 25789 5287
rect 25823 5253 25835 5287
rect 26326 5284 26332 5296
rect 25777 5247 25835 5253
rect 26068 5256 26332 5284
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 21358 5216 21364 5228
rect 21315 5188 21364 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 24486 5216 24492 5228
rect 23414 5188 24492 5216
rect 24486 5176 24492 5188
rect 24544 5176 24550 5228
rect 26068 5225 26096 5256
rect 26326 5244 26332 5256
rect 26384 5244 26390 5296
rect 26602 5284 26608 5296
rect 26515 5256 26608 5284
rect 26602 5244 26608 5256
rect 26660 5284 26666 5296
rect 28074 5284 28080 5296
rect 26660 5256 28080 5284
rect 26660 5244 26666 5256
rect 28074 5244 28080 5256
rect 28132 5244 28138 5296
rect 29840 5284 29868 5324
rect 30006 5312 30012 5324
rect 30064 5312 30070 5364
rect 34517 5355 34575 5361
rect 34517 5321 34529 5355
rect 34563 5352 34575 5355
rect 34606 5352 34612 5364
rect 34563 5324 34612 5352
rect 34563 5321 34575 5324
rect 34517 5315 34575 5321
rect 34606 5312 34612 5324
rect 34664 5312 34670 5364
rect 35802 5312 35808 5364
rect 35860 5352 35866 5364
rect 36081 5355 36139 5361
rect 36081 5352 36093 5355
rect 35860 5324 36093 5352
rect 35860 5312 35866 5324
rect 36081 5321 36093 5324
rect 36127 5352 36139 5355
rect 37461 5355 37519 5361
rect 37461 5352 37473 5355
rect 36127 5324 37473 5352
rect 36127 5321 36139 5324
rect 36081 5315 36139 5321
rect 37461 5321 37473 5324
rect 37507 5321 37519 5355
rect 37461 5315 37519 5321
rect 33873 5287 33931 5293
rect 33873 5284 33885 5287
rect 29840 5256 33885 5284
rect 33873 5253 33885 5256
rect 33919 5253 33931 5287
rect 33873 5247 33931 5253
rect 37918 5244 37924 5296
rect 37976 5284 37982 5296
rect 38013 5287 38071 5293
rect 38013 5284 38025 5287
rect 37976 5256 38025 5284
rect 37976 5244 37982 5256
rect 38013 5253 38025 5256
rect 38059 5253 38071 5287
rect 38013 5247 38071 5253
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5185 26111 5219
rect 27338 5216 27344 5228
rect 26053 5179 26111 5185
rect 26252 5188 27344 5216
rect 22002 5148 22008 5160
rect 21963 5120 22008 5148
rect 22002 5108 22008 5120
rect 22060 5108 22066 5160
rect 22281 5151 22339 5157
rect 22281 5148 22293 5151
rect 22112 5120 22293 5148
rect 22112 5080 22140 5120
rect 22281 5117 22293 5120
rect 22327 5148 22339 5151
rect 24578 5148 24584 5160
rect 22327 5120 24584 5148
rect 22327 5117 22339 5120
rect 22281 5111 22339 5117
rect 24578 5108 24584 5120
rect 24636 5108 24642 5160
rect 25130 5108 25136 5160
rect 25188 5148 25194 5160
rect 25188 5120 26004 5148
rect 25188 5108 25194 5120
rect 20548 5052 22140 5080
rect 23750 5040 23756 5092
rect 23808 5080 23814 5092
rect 25976 5080 26004 5120
rect 26252 5080 26280 5188
rect 27338 5176 27344 5188
rect 27396 5176 27402 5228
rect 26326 5108 26332 5160
rect 26384 5148 26390 5160
rect 28261 5151 28319 5157
rect 28261 5148 28273 5151
rect 26384 5120 28273 5148
rect 26384 5108 26390 5120
rect 28261 5117 28273 5120
rect 28307 5117 28319 5151
rect 28261 5111 28319 5117
rect 28537 5151 28595 5157
rect 28537 5117 28549 5151
rect 28583 5148 28595 5151
rect 29178 5148 29184 5160
rect 28583 5120 29184 5148
rect 28583 5117 28595 5120
rect 28537 5111 28595 5117
rect 29178 5108 29184 5120
rect 29236 5108 29242 5160
rect 23808 5052 24440 5080
rect 25976 5052 26280 5080
rect 23808 5040 23814 5052
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 14553 5015 14611 5021
rect 14553 4981 14565 5015
rect 14599 5012 14611 5015
rect 18230 5012 18236 5024
rect 14599 4984 18236 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 18690 4972 18696 5024
rect 18748 5012 18754 5024
rect 20165 5015 20223 5021
rect 20165 5012 20177 5015
rect 18748 4984 20177 5012
rect 18748 4972 18754 4984
rect 20165 4981 20177 4984
rect 20211 5012 20223 5015
rect 21174 5012 21180 5024
rect 20211 4984 21180 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 21361 5015 21419 5021
rect 21361 4981 21373 5015
rect 21407 5012 21419 5015
rect 22738 5012 22744 5024
rect 21407 4984 22744 5012
rect 21407 4981 21419 4984
rect 21361 4975 21419 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 22830 4972 22836 5024
rect 22888 5012 22894 5024
rect 24305 5015 24363 5021
rect 24305 5012 24317 5015
rect 22888 4984 24317 5012
rect 22888 4972 22894 4984
rect 24305 4981 24317 4984
rect 24351 4981 24363 5015
rect 24412 5012 24440 5052
rect 27249 5015 27307 5021
rect 27249 5012 27261 5015
rect 24412 4984 27261 5012
rect 24305 4975 24363 4981
rect 27249 4981 27261 4984
rect 27295 4981 27307 5015
rect 29656 5012 29684 5202
rect 30098 5176 30104 5228
rect 30156 5216 30162 5228
rect 30745 5219 30803 5225
rect 30745 5216 30757 5219
rect 30156 5188 30757 5216
rect 30156 5176 30162 5188
rect 30745 5185 30757 5188
rect 30791 5216 30803 5219
rect 31478 5216 31484 5228
rect 30791 5188 31484 5216
rect 30791 5185 30803 5188
rect 30745 5179 30803 5185
rect 31478 5176 31484 5188
rect 31536 5176 31542 5228
rect 32490 5216 32496 5228
rect 32451 5188 32496 5216
rect 32490 5176 32496 5188
rect 32548 5216 32554 5228
rect 33413 5219 33471 5225
rect 33413 5216 33425 5219
rect 32548 5188 33425 5216
rect 32548 5176 32554 5188
rect 33413 5185 33425 5188
rect 33459 5185 33471 5219
rect 33413 5179 33471 5185
rect 36630 5176 36636 5228
rect 36688 5216 36694 5228
rect 38194 5216 38200 5228
rect 36688 5188 38200 5216
rect 36688 5176 36694 5188
rect 38194 5176 38200 5188
rect 38252 5176 38258 5228
rect 30374 5108 30380 5160
rect 30432 5148 30438 5160
rect 30469 5151 30527 5157
rect 30469 5148 30481 5151
rect 30432 5120 30481 5148
rect 30432 5108 30438 5120
rect 30469 5117 30481 5120
rect 30515 5148 30527 5151
rect 30558 5148 30564 5160
rect 30515 5120 30564 5148
rect 30515 5117 30527 5120
rect 30469 5111 30527 5117
rect 30558 5108 30564 5120
rect 30616 5108 30622 5160
rect 32306 5040 32312 5092
rect 32364 5080 32370 5092
rect 36633 5083 36691 5089
rect 36633 5080 36645 5083
rect 32364 5052 36645 5080
rect 32364 5040 32370 5052
rect 36633 5049 36645 5052
rect 36679 5049 36691 5083
rect 36633 5043 36691 5049
rect 32122 5012 32128 5024
rect 29656 4984 32128 5012
rect 27249 4975 27307 4981
rect 32122 4972 32128 4984
rect 32180 4972 32186 5024
rect 32585 5015 32643 5021
rect 32585 4981 32597 5015
rect 32631 5012 32643 5015
rect 32766 5012 32772 5024
rect 32631 4984 32772 5012
rect 32631 4981 32643 4984
rect 32585 4975 32643 4981
rect 32766 4972 32772 4984
rect 32824 4972 32830 5024
rect 32858 4972 32864 5024
rect 32916 5012 32922 5024
rect 33321 5015 33379 5021
rect 33321 5012 33333 5015
rect 32916 4984 33333 5012
rect 32916 4972 32922 4984
rect 33321 4981 33333 4984
rect 33367 4981 33379 5015
rect 33321 4975 33379 4981
rect 34790 4972 34796 5024
rect 34848 5012 34854 5024
rect 34977 5015 35035 5021
rect 34977 5012 34989 5015
rect 34848 4984 34989 5012
rect 34848 4972 34854 4984
rect 34977 4981 34989 4984
rect 35023 5012 35035 5015
rect 35529 5015 35587 5021
rect 35529 5012 35541 5015
rect 35023 4984 35541 5012
rect 35023 4981 35035 4984
rect 34977 4975 35035 4981
rect 35529 4981 35541 4984
rect 35575 4981 35587 5015
rect 35529 4975 35587 4981
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 10318 4808 10324 4820
rect 10279 4780 10324 4808
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 14553 4811 14611 4817
rect 14553 4777 14565 4811
rect 14599 4808 14611 4811
rect 18138 4808 18144 4820
rect 14599 4780 18144 4808
rect 14599 4777 14611 4780
rect 14553 4771 14611 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 18414 4808 18420 4820
rect 18279 4780 18420 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 21910 4808 21916 4820
rect 18748 4780 21916 4808
rect 18748 4768 18754 4780
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 23934 4808 23940 4820
rect 22152 4780 23940 4808
rect 22152 4768 22158 4780
rect 23934 4768 23940 4780
rect 23992 4768 23998 4820
rect 24762 4768 24768 4820
rect 24820 4808 24826 4820
rect 24820 4780 26280 4808
rect 24820 4768 24826 4780
rect 13725 4743 13783 4749
rect 13725 4709 13737 4743
rect 13771 4740 13783 4743
rect 17494 4740 17500 4752
rect 13771 4712 17500 4740
rect 13771 4709 13783 4712
rect 13725 4703 13783 4709
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15804 4644 15849 4672
rect 15804 4632 15810 4644
rect 15930 4632 15936 4684
rect 15988 4672 15994 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 15988 4644 16405 4672
rect 15988 4632 15994 4644
rect 16393 4641 16405 4644
rect 16439 4672 16451 4675
rect 16850 4672 16856 4684
rect 16439 4644 16856 4672
rect 16439 4641 16451 4644
rect 16393 4635 16451 4641
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 17052 4681 17080 4712
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 17586 4700 17592 4752
rect 17644 4740 17650 4752
rect 20165 4743 20223 4749
rect 20165 4740 20177 4743
rect 17644 4712 20177 4740
rect 17644 4700 17650 4712
rect 20165 4709 20177 4712
rect 20211 4740 20223 4743
rect 20717 4743 20775 4749
rect 20717 4740 20729 4743
rect 20211 4712 20729 4740
rect 20211 4709 20223 4712
rect 20165 4703 20223 4709
rect 20717 4709 20729 4712
rect 20763 4740 20775 4743
rect 20898 4740 20904 4752
rect 20763 4712 20904 4740
rect 20763 4709 20775 4712
rect 20717 4703 20775 4709
rect 20898 4700 20904 4712
rect 20956 4700 20962 4752
rect 21177 4743 21235 4749
rect 21177 4709 21189 4743
rect 21223 4740 21235 4743
rect 21634 4740 21640 4752
rect 21223 4712 21640 4740
rect 21223 4709 21235 4712
rect 21177 4703 21235 4709
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 26252 4740 26280 4780
rect 30650 4768 30656 4820
rect 30708 4808 30714 4820
rect 31481 4811 31539 4817
rect 31481 4808 31493 4811
rect 30708 4780 31493 4808
rect 30708 4768 30714 4780
rect 31481 4777 31493 4780
rect 31527 4777 31539 4811
rect 31481 4771 31539 4777
rect 32493 4811 32551 4817
rect 32493 4777 32505 4811
rect 32539 4808 32551 4811
rect 33226 4808 33232 4820
rect 32539 4780 33232 4808
rect 32539 4777 32551 4780
rect 32493 4771 32551 4777
rect 33226 4768 33232 4780
rect 33284 4768 33290 4820
rect 26252 4712 27384 4740
rect 17037 4675 17095 4681
rect 17037 4641 17049 4675
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 17310 4632 17316 4684
rect 17368 4672 17374 4684
rect 18966 4672 18972 4684
rect 17368 4644 18972 4672
rect 17368 4632 17374 4644
rect 18966 4632 18972 4644
rect 19024 4672 19030 4684
rect 20254 4672 20260 4684
rect 19024 4644 20260 4672
rect 19024 4632 19030 4644
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 22002 4672 22008 4684
rect 21324 4644 22008 4672
rect 21324 4632 21330 4644
rect 22002 4632 22008 4644
rect 22060 4672 22066 4684
rect 22925 4675 22983 4681
rect 22925 4672 22937 4675
rect 22060 4644 22937 4672
rect 22060 4632 22066 4644
rect 22925 4641 22937 4644
rect 22971 4641 22983 4675
rect 25958 4672 25964 4684
rect 22925 4635 22983 4641
rect 23768 4644 25964 4672
rect 10410 4604 10416 4616
rect 10371 4576 10416 4604
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13688 4576 14473 4604
rect 13688 4564 13694 4576
rect 14461 4573 14473 4576
rect 14507 4604 14519 4607
rect 14507 4598 15608 4604
rect 15654 4598 15660 4616
rect 15712 4607 15718 4616
rect 18325 4607 18383 4613
rect 14507 4576 15660 4598
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 15580 4570 15660 4576
rect 15654 4564 15660 4570
rect 15712 4564 15723 4607
rect 18325 4573 18337 4607
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19242 4604 19248 4616
rect 18923 4576 19248 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 15665 4561 15723 4564
rect 17106 4539 17164 4545
rect 17106 4505 17118 4539
rect 17152 4536 17164 4539
rect 17681 4539 17739 4545
rect 17152 4505 17172 4536
rect 17106 4499 17172 4505
rect 17681 4505 17693 4539
rect 17727 4536 17739 4539
rect 17954 4536 17960 4548
rect 17727 4508 17960 4536
rect 17727 4505 17739 4508
rect 17681 4499 17739 4505
rect 14090 4428 14096 4480
rect 14148 4468 14154 4480
rect 14642 4468 14648 4480
rect 14148 4440 14648 4468
rect 14148 4428 14154 4440
rect 14642 4428 14648 4440
rect 14700 4468 14706 4480
rect 15197 4471 15255 4477
rect 15197 4468 15209 4471
rect 14700 4440 15209 4468
rect 14700 4428 14706 4440
rect 15197 4437 15209 4440
rect 15243 4468 15255 4471
rect 16574 4468 16580 4480
rect 15243 4440 16580 4468
rect 15243 4437 15255 4440
rect 15197 4431 15255 4437
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 17144 4468 17172 4499
rect 17218 4468 17224 4480
rect 17144 4440 17224 4468
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 17696 4468 17724 4499
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 18340 4536 18368 4567
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 20772 4576 21574 4604
rect 20772 4564 20778 4576
rect 18340 4508 21312 4536
rect 17368 4440 17724 4468
rect 17368 4428 17374 4440
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18874 4468 18880 4480
rect 17828 4440 18880 4468
rect 17828 4428 17834 4440
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19521 4471 19579 4477
rect 19521 4468 19533 4471
rect 19484 4440 19533 4468
rect 19484 4428 19490 4440
rect 19521 4437 19533 4440
rect 19567 4437 19579 4471
rect 21284 4468 21312 4508
rect 22554 4496 22560 4548
rect 22612 4536 22618 4548
rect 22649 4539 22707 4545
rect 22649 4536 22661 4539
rect 22612 4508 22661 4536
rect 22612 4496 22618 4508
rect 22649 4505 22661 4508
rect 22695 4505 22707 4539
rect 22649 4499 22707 4505
rect 23768 4468 23796 4644
rect 25958 4632 25964 4644
rect 26016 4632 26022 4684
rect 26053 4675 26111 4681
rect 26053 4641 26065 4675
rect 26099 4672 26111 4675
rect 26418 4672 26424 4684
rect 26099 4644 26424 4672
rect 26099 4641 26111 4644
rect 26053 4635 26111 4641
rect 26418 4632 26424 4644
rect 26476 4632 26482 4684
rect 27356 4672 27384 4712
rect 32674 4700 32680 4752
rect 32732 4740 32738 4752
rect 36173 4743 36231 4749
rect 36173 4740 36185 4743
rect 32732 4712 36185 4740
rect 32732 4700 32738 4712
rect 36173 4709 36185 4712
rect 36219 4709 36231 4743
rect 36173 4703 36231 4709
rect 28537 4675 28595 4681
rect 28537 4672 28549 4675
rect 27356 4644 28549 4672
rect 28537 4641 28549 4644
rect 28583 4672 28595 4675
rect 31386 4672 31392 4684
rect 28583 4644 31392 4672
rect 28583 4641 28595 4644
rect 28537 4635 28595 4641
rect 31386 4632 31392 4644
rect 31444 4632 31450 4684
rect 31726 4644 33272 4672
rect 23842 4564 23848 4616
rect 23900 4604 23906 4616
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 23900 4576 24041 4604
rect 23900 4564 23906 4576
rect 24029 4573 24041 4576
rect 24075 4573 24087 4607
rect 24029 4567 24087 4573
rect 24946 4564 24952 4616
rect 25004 4564 25010 4616
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 28813 4607 28871 4613
rect 26384 4576 26429 4604
rect 26384 4564 26390 4576
rect 28813 4573 28825 4607
rect 28859 4604 28871 4607
rect 28994 4604 29000 4616
rect 28859 4576 29000 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 28994 4564 29000 4576
rect 29052 4604 29058 4616
rect 29730 4604 29736 4616
rect 29052 4576 29736 4604
rect 29052 4564 29058 4576
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 31294 4604 31300 4616
rect 31142 4576 31300 4604
rect 31294 4564 31300 4576
rect 31352 4564 31358 4616
rect 28106 4508 28488 4536
rect 23934 4468 23940 4480
rect 21284 4440 23796 4468
rect 23895 4440 23940 4468
rect 19521 4431 19579 4437
rect 23934 4428 23940 4440
rect 23992 4428 23998 4480
rect 24581 4471 24639 4477
rect 24581 4437 24593 4471
rect 24627 4468 24639 4471
rect 25038 4468 25044 4480
rect 24627 4440 25044 4468
rect 24627 4437 24639 4440
rect 24581 4431 24639 4437
rect 25038 4428 25044 4440
rect 25096 4428 25102 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 27065 4471 27123 4477
rect 27065 4468 27077 4471
rect 26292 4440 27077 4468
rect 26292 4428 26298 4440
rect 27065 4437 27077 4440
rect 27111 4437 27123 4471
rect 28460 4468 28488 4508
rect 28902 4496 28908 4548
rect 28960 4536 28966 4548
rect 30009 4539 30067 4545
rect 30009 4536 30021 4539
rect 28960 4508 30021 4536
rect 28960 4496 28966 4508
rect 30009 4505 30021 4508
rect 30055 4505 30067 4539
rect 31726 4536 31754 4644
rect 32306 4604 32312 4616
rect 32267 4576 32312 4604
rect 32306 4564 32312 4576
rect 32364 4564 32370 4616
rect 33244 4604 33272 4644
rect 33318 4632 33324 4684
rect 33376 4672 33382 4684
rect 35529 4675 35587 4681
rect 35529 4672 35541 4675
rect 33376 4644 35541 4672
rect 33376 4632 33382 4644
rect 35529 4641 35541 4644
rect 35575 4641 35587 4675
rect 35529 4635 35587 4641
rect 34054 4604 34060 4616
rect 33244 4576 34060 4604
rect 34054 4564 34060 4576
rect 34112 4564 34118 4616
rect 34241 4607 34299 4613
rect 34241 4573 34253 4607
rect 34287 4604 34299 4607
rect 34514 4604 34520 4616
rect 34287 4576 34520 4604
rect 34287 4573 34299 4576
rect 34241 4567 34299 4573
rect 34514 4564 34520 4576
rect 34572 4604 34578 4616
rect 35621 4607 35679 4613
rect 35621 4604 35633 4607
rect 34572 4576 35633 4604
rect 34572 4564 34578 4576
rect 35621 4573 35633 4576
rect 35667 4604 35679 4607
rect 36265 4607 36323 4613
rect 36265 4604 36277 4607
rect 35667 4576 36277 4604
rect 35667 4573 35679 4576
rect 35621 4567 35679 4573
rect 36265 4573 36277 4576
rect 36311 4573 36323 4607
rect 37826 4604 37832 4616
rect 37787 4576 37832 4604
rect 36265 4567 36323 4573
rect 37826 4564 37832 4576
rect 37884 4564 37890 4616
rect 30009 4499 30067 4505
rect 31312 4508 31754 4536
rect 33045 4539 33103 4545
rect 31312 4468 31340 4508
rect 33045 4505 33057 4539
rect 33091 4536 33103 4539
rect 33410 4536 33416 4548
rect 33091 4508 33416 4536
rect 33091 4505 33103 4508
rect 33045 4499 33103 4505
rect 33410 4496 33416 4508
rect 33468 4536 33474 4548
rect 33597 4539 33655 4545
rect 33597 4536 33609 4539
rect 33468 4508 33609 4536
rect 33468 4496 33474 4508
rect 33597 4505 33609 4508
rect 33643 4536 33655 4539
rect 33643 4508 34928 4536
rect 33643 4505 33655 4508
rect 33597 4499 33655 4505
rect 34900 4480 34928 4508
rect 36078 4496 36084 4548
rect 36136 4536 36142 4548
rect 36725 4539 36783 4545
rect 36725 4536 36737 4539
rect 36136 4508 36737 4536
rect 36136 4496 36142 4508
rect 36725 4505 36737 4508
rect 36771 4505 36783 4539
rect 36725 4499 36783 4505
rect 28460 4440 31340 4468
rect 27065 4431 27123 4437
rect 31570 4428 31576 4480
rect 31628 4468 31634 4480
rect 33502 4468 33508 4480
rect 31628 4440 33508 4468
rect 31628 4428 31634 4440
rect 33502 4428 33508 4440
rect 33560 4428 33566 4480
rect 34146 4468 34152 4480
rect 34107 4440 34152 4468
rect 34146 4428 34152 4440
rect 34204 4428 34210 4480
rect 34882 4468 34888 4480
rect 34843 4440 34888 4468
rect 34882 4428 34888 4440
rect 34940 4428 34946 4480
rect 36262 4428 36268 4480
rect 36320 4468 36326 4480
rect 37737 4471 37795 4477
rect 37737 4468 37749 4471
rect 36320 4440 37749 4468
rect 36320 4428 36326 4440
rect 37737 4437 37749 4440
rect 37783 4437 37795 4471
rect 37737 4431 37795 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 15396 4236 16620 4264
rect 14642 4196 14648 4208
rect 14603 4168 14648 4196
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 10008 4100 13461 4128
rect 10008 4088 10014 4100
rect 13449 4097 13461 4100
rect 13495 4128 13507 4131
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13495 4100 14013 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 14001 4097 14013 4100
rect 14047 4128 14059 4131
rect 14090 4128 14096 4140
rect 14047 4100 14096 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14921 4131 14979 4137
rect 14921 4128 14933 4131
rect 14516 4100 14933 4128
rect 14516 4088 14522 4100
rect 14921 4097 14933 4100
rect 14967 4128 14979 4131
rect 15396 4128 15424 4236
rect 15654 4196 15660 4208
rect 15488 4168 15660 4196
rect 15488 4137 15516 4168
rect 15654 4156 15660 4168
rect 15712 4196 15718 4208
rect 16482 4196 16488 4208
rect 15712 4168 16488 4196
rect 15712 4156 15718 4168
rect 16482 4156 16488 4168
rect 16540 4156 16546 4208
rect 14967 4100 15424 4128
rect 15473 4131 15531 4137
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15473 4097 15485 4131
rect 15519 4097 15531 4131
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 15473 4091 15531 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16592 4128 16620 4236
rect 17034 4224 17040 4276
rect 17092 4264 17098 4276
rect 17092 4236 19564 4264
rect 17092 4224 17098 4236
rect 17589 4199 17647 4205
rect 17589 4165 17601 4199
rect 17635 4196 17647 4199
rect 17954 4196 17960 4208
rect 17635 4168 17960 4196
rect 17635 4165 17647 4168
rect 17589 4159 17647 4165
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 19536 4196 19564 4236
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 22094 4264 22100 4276
rect 20036 4236 22100 4264
rect 20036 4224 20042 4236
rect 22094 4224 22100 4236
rect 22152 4224 22158 4276
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 25038 4264 25044 4276
rect 22244 4236 22289 4264
rect 23124 4236 25044 4264
rect 22244 4224 22250 4236
rect 23124 4196 23152 4236
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 25130 4224 25136 4276
rect 25188 4264 25194 4276
rect 28718 4264 28724 4276
rect 25188 4236 28724 4264
rect 25188 4224 25194 4236
rect 28718 4224 28724 4236
rect 28776 4224 28782 4276
rect 32858 4264 32864 4276
rect 29564 4236 32864 4264
rect 19536 4168 23152 4196
rect 23934 4156 23940 4208
rect 23992 4156 23998 4208
rect 24394 4196 24400 4208
rect 24355 4168 24400 4196
rect 24394 4156 24400 4168
rect 24452 4156 24458 4208
rect 26326 4196 26332 4208
rect 24688 4168 26332 4196
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 16592 4100 17233 4128
rect 17221 4097 17233 4100
rect 17267 4097 17279 4131
rect 18230 4128 18236 4140
rect 18191 4100 18236 4128
rect 17221 4091 17279 4097
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4097 18383 4131
rect 18966 4128 18972 4140
rect 18927 4100 18972 4128
rect 18325 4091 18383 4097
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 18138 4060 18144 4072
rect 15611 4032 18144 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 18340 4060 18368 4091
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19610 4088 19616 4140
rect 19668 4128 19674 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 19668 4100 22017 4128
rect 19668 4088 19674 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 23106 4128 23112 4140
rect 22005 4091 22063 4097
rect 22112 4100 23112 4128
rect 22112 4060 22140 4100
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 24688 4072 24716 4168
rect 26326 4156 26332 4168
rect 26384 4156 26390 4208
rect 26602 4196 26608 4208
rect 26563 4168 26608 4196
rect 26602 4156 26608 4168
rect 26660 4156 26666 4208
rect 29564 4196 29592 4236
rect 32858 4224 32864 4236
rect 32916 4224 32922 4276
rect 33410 4264 33416 4276
rect 33371 4236 33416 4264
rect 33410 4224 33416 4236
rect 33468 4224 33474 4276
rect 34054 4224 34060 4276
rect 34112 4264 34118 4276
rect 37366 4264 37372 4276
rect 34112 4236 37372 4264
rect 34112 4224 34118 4236
rect 37366 4224 37372 4236
rect 37424 4224 37430 4276
rect 36262 4196 36268 4208
rect 28198 4168 29592 4196
rect 30406 4168 36268 4196
rect 36262 4156 36268 4168
rect 36320 4156 36326 4208
rect 25777 4131 25835 4137
rect 25777 4097 25789 4131
rect 25823 4128 25835 4131
rect 25866 4128 25872 4140
rect 25823 4100 25872 4128
rect 25823 4097 25835 4100
rect 25777 4091 25835 4097
rect 25866 4088 25872 4100
rect 25924 4088 25930 4140
rect 28905 4131 28963 4137
rect 26068 4100 27476 4128
rect 24670 4060 24676 4072
rect 18340 4032 22140 4060
rect 24631 4032 24676 4060
rect 24670 4020 24676 4032
rect 24728 4020 24734 4072
rect 25130 4020 25136 4072
rect 25188 4060 25194 4072
rect 26068 4069 26096 4100
rect 26053 4063 26111 4069
rect 26053 4060 26065 4063
rect 25188 4032 26065 4060
rect 25188 4020 25194 4032
rect 26053 4029 26065 4032
rect 26099 4029 26111 4063
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 26053 4023 26111 4029
rect 26160 4032 27169 4060
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 19426 3992 19432 4004
rect 13964 3964 19432 3992
rect 13964 3952 13970 3964
rect 19426 3952 19432 3964
rect 19484 3992 19490 4004
rect 19705 3995 19763 4001
rect 19705 3992 19717 3995
rect 19484 3964 19717 3992
rect 19484 3952 19490 3964
rect 19705 3961 19717 3964
rect 19751 3992 19763 3995
rect 20257 3995 20315 4001
rect 20257 3992 20269 3995
rect 19751 3964 20269 3992
rect 19751 3961 19763 3964
rect 19705 3955 19763 3961
rect 20257 3961 20269 3964
rect 20303 3992 20315 3995
rect 21266 3992 21272 4004
rect 20303 3964 21272 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 22094 3992 22100 4004
rect 21376 3964 22100 3992
rect 16209 3927 16267 3933
rect 16209 3893 16221 3927
rect 16255 3924 16267 3927
rect 18046 3924 18052 3936
rect 16255 3896 18052 3924
rect 16255 3893 16267 3896
rect 16209 3887 16267 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 18877 3927 18935 3933
rect 18877 3924 18889 3927
rect 18288 3896 18889 3924
rect 18288 3884 18294 3896
rect 18877 3893 18889 3896
rect 18923 3893 18935 3927
rect 18877 3887 18935 3893
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 20588 3896 20821 3924
rect 20588 3884 20594 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 20898 3884 20904 3936
rect 20956 3924 20962 3936
rect 21376 3924 21404 3964
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 22278 3952 22284 4004
rect 22336 3992 22342 4004
rect 22925 3995 22983 4001
rect 22925 3992 22937 3995
rect 22336 3964 22937 3992
rect 22336 3952 22342 3964
rect 22925 3961 22937 3964
rect 22971 3961 22983 3995
rect 22925 3955 22983 3961
rect 24762 3952 24768 4004
rect 24820 3992 24826 4004
rect 25866 3992 25872 4004
rect 24820 3964 25872 3992
rect 24820 3952 24826 3964
rect 25866 3952 25872 3964
rect 25924 3952 25930 4004
rect 25958 3952 25964 4004
rect 26016 3992 26022 4004
rect 26160 3992 26188 4032
rect 27157 4029 27169 4032
rect 27203 4060 27215 4063
rect 27338 4060 27344 4072
rect 27203 4032 27344 4060
rect 27203 4029 27215 4032
rect 27157 4023 27215 4029
rect 27338 4020 27344 4032
rect 27396 4020 27402 4072
rect 27448 4060 27476 4100
rect 28905 4097 28917 4131
rect 28951 4128 28963 4131
rect 28994 4128 29000 4140
rect 28951 4100 29000 4128
rect 28951 4097 28963 4100
rect 28905 4091 28963 4097
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 31573 4131 31631 4137
rect 31573 4128 31585 4131
rect 31536 4100 31585 4128
rect 31536 4088 31542 4100
rect 31573 4097 31585 4100
rect 31619 4097 31631 4131
rect 31573 4091 31631 4097
rect 32677 4131 32735 4137
rect 32677 4097 32689 4131
rect 32723 4128 32735 4131
rect 33226 4128 33232 4140
rect 32723 4100 33232 4128
rect 32723 4097 32735 4100
rect 32677 4091 32735 4097
rect 33226 4088 33232 4100
rect 33284 4088 33290 4140
rect 36909 4131 36967 4137
rect 36909 4097 36921 4131
rect 36955 4097 36967 4131
rect 36909 4091 36967 4097
rect 37737 4131 37795 4137
rect 37737 4097 37749 4131
rect 37783 4128 37795 4131
rect 37826 4128 37832 4140
rect 37783 4100 37832 4128
rect 37783 4097 37795 4100
rect 37737 4091 37795 4097
rect 29362 4060 29368 4072
rect 27448 4032 28856 4060
rect 29323 4032 29368 4060
rect 28828 3992 28856 4032
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 31113 4063 31171 4069
rect 29472 4032 31064 4060
rect 29472 3992 29500 4032
rect 26016 3964 26188 3992
rect 26436 3964 27660 3992
rect 28828 3964 29500 3992
rect 31036 3992 31064 4032
rect 31113 4029 31125 4063
rect 31159 4060 31171 4063
rect 31202 4060 31208 4072
rect 31159 4032 31208 4060
rect 31159 4029 31171 4032
rect 31113 4023 31171 4029
rect 31202 4020 31208 4032
rect 31260 4060 31266 4072
rect 32122 4060 32128 4072
rect 31260 4032 32128 4060
rect 31260 4020 31266 4032
rect 32122 4020 32128 4032
rect 32180 4020 32186 4072
rect 36817 4063 36875 4069
rect 36817 4060 36829 4063
rect 32324 4032 36829 4060
rect 31662 3992 31668 4004
rect 31036 3964 31668 3992
rect 26016 3952 26022 3964
rect 20956 3896 21404 3924
rect 20956 3884 20962 3896
rect 21450 3884 21456 3936
rect 21508 3924 21514 3936
rect 21508 3896 21553 3924
rect 21508 3884 21514 3896
rect 24026 3884 24032 3936
rect 24084 3924 24090 3936
rect 26436 3924 26464 3964
rect 24084 3896 26464 3924
rect 27632 3924 27660 3964
rect 31662 3952 31668 3964
rect 31720 3952 31726 4004
rect 31938 3952 31944 4004
rect 31996 3992 32002 4004
rect 32324 3992 32352 4032
rect 36817 4029 36829 4032
rect 36863 4029 36875 4063
rect 36924 4060 36952 4091
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 37550 4060 37556 4072
rect 36924 4032 37556 4060
rect 36817 4023 36875 4029
rect 37550 4020 37556 4032
rect 37608 4060 37614 4072
rect 38102 4060 38108 4072
rect 37608 4032 38108 4060
rect 37608 4020 37614 4032
rect 38102 4020 38108 4032
rect 38160 4020 38166 4072
rect 31996 3964 32352 3992
rect 32861 3995 32919 4001
rect 31996 3952 32002 3964
rect 32861 3961 32873 3995
rect 32907 3992 32919 3995
rect 34330 3992 34336 4004
rect 32907 3964 34336 3992
rect 32907 3961 32919 3964
rect 32861 3955 32919 3961
rect 34330 3952 34336 3964
rect 34388 3952 34394 4004
rect 36630 3952 36636 4004
rect 36688 3992 36694 4004
rect 37645 3995 37703 4001
rect 37645 3992 37657 3995
rect 36688 3964 37657 3992
rect 36688 3952 36694 3964
rect 37645 3961 37657 3964
rect 37691 3961 37703 3995
rect 37645 3955 37703 3961
rect 28442 3924 28448 3936
rect 27632 3896 28448 3924
rect 24084 3884 24090 3896
rect 28442 3884 28448 3896
rect 28500 3884 28506 3936
rect 28626 3884 28632 3936
rect 28684 3933 28690 3936
rect 28684 3927 28699 3933
rect 28687 3893 28699 3927
rect 28684 3887 28699 3893
rect 30855 3927 30913 3933
rect 30855 3893 30867 3927
rect 30901 3924 30913 3927
rect 31110 3924 31116 3936
rect 30901 3896 31116 3924
rect 30901 3893 30913 3896
rect 30855 3887 30913 3893
rect 28684 3884 28690 3887
rect 31110 3884 31116 3896
rect 31168 3924 31174 3936
rect 31478 3924 31484 3936
rect 31168 3896 31484 3924
rect 31168 3884 31174 3896
rect 31478 3884 31484 3896
rect 31536 3884 31542 3936
rect 31757 3927 31815 3933
rect 31757 3893 31769 3927
rect 31803 3924 31815 3927
rect 33502 3924 33508 3936
rect 31803 3896 33508 3924
rect 31803 3893 31815 3896
rect 31757 3887 31815 3893
rect 33502 3884 33508 3896
rect 33560 3884 33566 3936
rect 33870 3924 33876 3936
rect 33831 3896 33876 3924
rect 33870 3884 33876 3896
rect 33928 3884 33934 3936
rect 34517 3927 34575 3933
rect 34517 3893 34529 3927
rect 34563 3924 34575 3927
rect 34882 3924 34888 3936
rect 34563 3896 34888 3924
rect 34563 3893 34575 3896
rect 34517 3887 34575 3893
rect 34882 3884 34888 3896
rect 34940 3924 34946 3936
rect 35069 3927 35127 3933
rect 35069 3924 35081 3927
rect 34940 3896 35081 3924
rect 34940 3884 34946 3896
rect 35069 3893 35081 3896
rect 35115 3924 35127 3927
rect 35621 3927 35679 3933
rect 35621 3924 35633 3927
rect 35115 3896 35633 3924
rect 35115 3893 35127 3896
rect 35069 3887 35127 3893
rect 35621 3893 35633 3896
rect 35667 3924 35679 3927
rect 36078 3924 36084 3936
rect 35667 3896 36084 3924
rect 35667 3893 35679 3896
rect 35621 3887 35679 3893
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 38194 3924 38200 3936
rect 38155 3896 38200 3924
rect 38194 3884 38200 3896
rect 38252 3884 38258 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 12069 3723 12127 3729
rect 12069 3689 12081 3723
rect 12115 3720 12127 3723
rect 13173 3723 13231 3729
rect 12115 3692 12434 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 12406 3652 12434 3692
rect 13173 3689 13185 3723
rect 13219 3720 13231 3723
rect 14090 3720 14096 3732
rect 13219 3692 14096 3720
rect 13219 3689 13231 3692
rect 13173 3683 13231 3689
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 17218 3720 17224 3732
rect 16163 3692 17224 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 19426 3720 19432 3732
rect 17736 3692 19432 3720
rect 17736 3680 17742 3692
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 19610 3720 19616 3732
rect 19571 3692 19616 3720
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 21526 3723 21584 3729
rect 21526 3720 21538 3723
rect 19944 3692 21538 3720
rect 19944 3680 19950 3692
rect 21526 3689 21538 3692
rect 21572 3720 21584 3723
rect 21910 3720 21916 3732
rect 21572 3692 21916 3720
rect 21572 3689 21584 3692
rect 21526 3683 21584 3689
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22186 3680 22192 3732
rect 22244 3720 22250 3732
rect 28273 3723 28331 3729
rect 28273 3720 28285 3723
rect 22244 3692 28285 3720
rect 22244 3680 22250 3692
rect 28273 3689 28285 3692
rect 28319 3689 28331 3723
rect 28273 3683 28331 3689
rect 28442 3680 28448 3732
rect 28500 3720 28506 3732
rect 31570 3720 31576 3732
rect 28500 3692 31576 3720
rect 28500 3680 28506 3692
rect 31570 3680 31576 3692
rect 31628 3680 31634 3732
rect 31662 3680 31668 3732
rect 31720 3720 31726 3732
rect 33870 3720 33876 3732
rect 31720 3692 33876 3720
rect 31720 3680 31726 3692
rect 33870 3680 33876 3692
rect 33928 3680 33934 3732
rect 15930 3652 15936 3664
rect 12406 3624 15936 3652
rect 15930 3612 15936 3624
rect 15988 3612 15994 3664
rect 16224 3624 21404 3652
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3516 1642 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1636 3488 2237 3516
rect 1636 3476 1642 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12434 3516 12440 3528
rect 12207 3488 12440 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 12434 3476 12440 3488
rect 12492 3516 12498 3528
rect 14458 3516 14464 3528
rect 12492 3488 14464 3516
rect 12492 3476 12498 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 16224 3525 16252 3624
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 16540 3556 17693 3584
rect 16540 3544 16546 3556
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 18138 3544 18144 3596
rect 18196 3584 18202 3596
rect 20990 3584 20996 3596
rect 18196 3556 20996 3584
rect 18196 3544 18202 3556
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 21376 3584 21404 3624
rect 22922 3612 22928 3664
rect 22980 3652 22986 3664
rect 23017 3655 23075 3661
rect 23017 3652 23029 3655
rect 22980 3624 23029 3652
rect 22980 3612 22986 3624
rect 23017 3621 23029 3624
rect 23063 3621 23075 3655
rect 23017 3615 23075 3621
rect 23106 3612 23112 3664
rect 23164 3652 23170 3664
rect 24946 3652 24952 3664
rect 23164 3624 24952 3652
rect 23164 3612 23170 3624
rect 24946 3612 24952 3624
rect 25004 3612 25010 3664
rect 31110 3612 31116 3664
rect 31168 3652 31174 3664
rect 31754 3652 31760 3664
rect 31168 3624 31760 3652
rect 31168 3612 31174 3624
rect 31754 3612 31760 3624
rect 31812 3612 31818 3664
rect 33226 3612 33232 3664
rect 33284 3652 33290 3664
rect 33686 3652 33692 3664
rect 33284 3624 33692 3652
rect 33284 3612 33290 3624
rect 33686 3612 33692 3624
rect 33744 3612 33750 3664
rect 33962 3612 33968 3664
rect 34020 3652 34026 3664
rect 34020 3624 36952 3652
rect 34020 3612 34026 3624
rect 21634 3584 21640 3596
rect 21376 3556 21640 3584
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 26053 3587 26111 3593
rect 26053 3584 26065 3587
rect 21968 3556 26065 3584
rect 21968 3544 21974 3556
rect 26053 3553 26065 3556
rect 26099 3553 26111 3587
rect 26326 3584 26332 3596
rect 26287 3556 26332 3584
rect 26053 3547 26111 3553
rect 26326 3544 26332 3556
rect 26384 3584 26390 3596
rect 28537 3587 28595 3593
rect 28537 3584 28549 3587
rect 26384 3556 28549 3584
rect 26384 3544 26390 3556
rect 28537 3553 28549 3556
rect 28583 3584 28595 3587
rect 29089 3587 29147 3593
rect 29089 3584 29101 3587
rect 28583 3556 29101 3584
rect 28583 3553 28595 3556
rect 28537 3547 28595 3553
rect 29089 3553 29101 3556
rect 29135 3584 29147 3587
rect 29730 3584 29736 3596
rect 29135 3556 29736 3584
rect 29135 3553 29147 3556
rect 29089 3547 29147 3553
rect 29730 3544 29736 3556
rect 29788 3584 29794 3596
rect 31202 3584 31208 3596
rect 29788 3556 31208 3584
rect 29788 3544 29794 3556
rect 31202 3544 31208 3556
rect 31260 3584 31266 3596
rect 31930 3587 31988 3593
rect 31930 3584 31942 3587
rect 31260 3556 31942 3584
rect 31260 3544 31266 3556
rect 31930 3553 31942 3556
rect 31976 3553 31988 3587
rect 36924 3584 36952 3624
rect 37366 3612 37372 3664
rect 37424 3652 37430 3664
rect 37461 3655 37519 3661
rect 37461 3652 37473 3655
rect 37424 3624 37473 3652
rect 37424 3612 37430 3624
rect 37461 3621 37473 3624
rect 37507 3621 37519 3655
rect 37461 3615 37519 3621
rect 38013 3587 38071 3593
rect 38013 3584 38025 3587
rect 36924 3556 38025 3584
rect 31930 3547 31988 3553
rect 38013 3553 38025 3556
rect 38059 3553 38071 3587
rect 38013 3547 38071 3553
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3485 16267 3519
rect 16850 3516 16856 3528
rect 16763 3488 16856 3516
rect 16209 3479 16267 3485
rect 16850 3476 16856 3488
rect 16908 3516 16914 3528
rect 16908 3488 17816 3516
rect 16908 3476 16914 3488
rect 15289 3451 15347 3457
rect 15289 3417 15301 3451
rect 15335 3448 15347 3451
rect 16666 3448 16672 3460
rect 15335 3420 16672 3448
rect 15335 3417 15347 3420
rect 15289 3411 15347 3417
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 17788 3448 17816 3488
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18012 3488 18429 3516
rect 18012 3476 18018 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18417 3479 18475 3485
rect 18524 3488 19441 3516
rect 18524 3448 18552 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3485 20131 3519
rect 23750 3516 23756 3528
rect 22678 3488 23756 3516
rect 20073 3479 20131 3485
rect 18690 3448 18696 3460
rect 16776 3420 17632 3448
rect 17788 3420 18552 3448
rect 18651 3420 18696 3448
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 16776 3380 16804 3420
rect 13771 3352 16804 3380
rect 16853 3383 16911 3389
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 16853 3349 16865 3383
rect 16899 3380 16911 3383
rect 17126 3380 17132 3392
rect 16899 3352 17132 3380
rect 16899 3349 16911 3352
rect 16853 3343 16911 3349
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 17604 3380 17632 3420
rect 18690 3408 18696 3420
rect 18748 3408 18754 3460
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 20088 3448 20116 3479
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 24026 3516 24032 3528
rect 23987 3488 24032 3516
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 37550 3516 37556 3528
rect 37511 3488 37556 3516
rect 37550 3476 37556 3488
rect 37608 3476 37614 3528
rect 38197 3519 38255 3525
rect 38197 3485 38209 3519
rect 38243 3516 38255 3519
rect 38286 3516 38292 3528
rect 38243 3488 38292 3516
rect 38243 3485 38255 3488
rect 38197 3479 38255 3485
rect 38286 3476 38292 3488
rect 38344 3516 38350 3528
rect 39298 3516 39304 3528
rect 38344 3488 39304 3516
rect 38344 3476 38350 3488
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 19392 3420 20116 3448
rect 19392 3408 19398 3420
rect 22922 3408 22928 3460
rect 22980 3448 22986 3460
rect 23474 3448 23480 3460
rect 22980 3420 23480 3448
rect 22980 3408 22986 3420
rect 23474 3408 23480 3420
rect 23532 3408 23538 3460
rect 25314 3408 25320 3460
rect 25372 3408 25378 3460
rect 25774 3408 25780 3460
rect 25832 3448 25838 3460
rect 30009 3451 30067 3457
rect 25832 3420 27094 3448
rect 25832 3408 25838 3420
rect 30009 3417 30021 3451
rect 30055 3417 30067 3451
rect 31938 3448 31944 3460
rect 31234 3420 31944 3448
rect 30009 3411 30067 3417
rect 19886 3380 19892 3392
rect 17604 3352 19892 3380
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 19978 3340 19984 3392
rect 20036 3380 20042 3392
rect 20257 3383 20315 3389
rect 20257 3380 20269 3383
rect 20036 3352 20269 3380
rect 20036 3340 20042 3352
rect 20257 3349 20269 3352
rect 20303 3349 20315 3383
rect 23842 3380 23848 3392
rect 23803 3352 23848 3380
rect 20257 3343 20315 3349
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 24394 3340 24400 3392
rect 24452 3380 24458 3392
rect 24581 3383 24639 3389
rect 24581 3380 24593 3383
rect 24452 3352 24593 3380
rect 24452 3340 24458 3352
rect 24581 3349 24593 3352
rect 24627 3349 24639 3383
rect 24581 3343 24639 3349
rect 26142 3340 26148 3392
rect 26200 3380 26206 3392
rect 26789 3383 26847 3389
rect 26789 3380 26801 3383
rect 26200 3352 26801 3380
rect 26200 3340 26206 3352
rect 26789 3349 26801 3352
rect 26835 3349 26847 3383
rect 26789 3343 26847 3349
rect 26878 3340 26884 3392
rect 26936 3380 26942 3392
rect 30024 3380 30052 3411
rect 31938 3408 31944 3420
rect 31996 3408 32002 3460
rect 32214 3448 32220 3460
rect 32175 3420 32220 3448
rect 32214 3408 32220 3420
rect 32272 3408 32278 3460
rect 34146 3448 34152 3460
rect 33442 3420 34152 3448
rect 34146 3408 34152 3420
rect 34204 3408 34210 3460
rect 34238 3408 34244 3460
rect 34296 3448 34302 3460
rect 34977 3451 35035 3457
rect 34977 3448 34989 3451
rect 34296 3420 34989 3448
rect 34296 3408 34302 3420
rect 34977 3417 34989 3420
rect 35023 3448 35035 3451
rect 35529 3451 35587 3457
rect 35529 3448 35541 3451
rect 35023 3420 35541 3448
rect 35023 3417 35035 3420
rect 34977 3411 35035 3417
rect 35529 3417 35541 3420
rect 35575 3448 35587 3451
rect 36078 3448 36084 3460
rect 35575 3420 36084 3448
rect 35575 3417 35587 3420
rect 35529 3411 35587 3417
rect 36078 3408 36084 3420
rect 36136 3448 36142 3460
rect 36136 3420 36676 3448
rect 36136 3408 36142 3420
rect 26936 3352 30052 3380
rect 26936 3340 26942 3352
rect 31386 3340 31392 3392
rect 31444 3380 31450 3392
rect 31481 3383 31539 3389
rect 31481 3380 31493 3383
rect 31444 3352 31493 3380
rect 31444 3340 31450 3352
rect 31481 3349 31493 3352
rect 31527 3349 31539 3383
rect 31481 3343 31539 3349
rect 31570 3340 31576 3392
rect 31628 3380 31634 3392
rect 33594 3380 33600 3392
rect 31628 3352 33600 3380
rect 31628 3340 31634 3352
rect 33594 3340 33600 3352
rect 33652 3340 33658 3392
rect 33686 3340 33692 3392
rect 33744 3380 33750 3392
rect 36354 3380 36360 3392
rect 33744 3352 36360 3380
rect 33744 3340 33750 3352
rect 36354 3340 36360 3352
rect 36412 3340 36418 3392
rect 36648 3389 36676 3420
rect 36633 3383 36691 3389
rect 36633 3349 36645 3383
rect 36679 3380 36691 3383
rect 37550 3380 37556 3392
rect 36679 3352 37556 3380
rect 36679 3349 36691 3352
rect 36633 3343 36691 3349
rect 37550 3340 37556 3352
rect 37608 3340 37614 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3145 4767 3179
rect 10042 3176 10048 3188
rect 4709 3139 4767 3145
rect 6886 3148 10048 3176
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 4724 3040 4752 3139
rect 1903 3012 4752 3040
rect 4893 3043 4951 3049
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 6886 3040 6914 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 13044 3148 13369 3176
rect 13044 3136 13050 3148
rect 13357 3145 13369 3148
rect 13403 3176 13415 3179
rect 31754 3176 31760 3188
rect 13403 3148 31760 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 14274 3108 14280 3120
rect 8404 3080 14280 3108
rect 8404 3049 8432 3080
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 14458 3068 14464 3120
rect 14516 3108 14522 3120
rect 17126 3108 17132 3120
rect 14516 3080 14872 3108
rect 17087 3080 17132 3108
rect 14516 3068 14522 3080
rect 14844 3049 14872 3080
rect 17126 3068 17132 3080
rect 17184 3068 17190 3120
rect 17221 3111 17279 3117
rect 17221 3077 17233 3111
rect 17267 3108 17279 3111
rect 18230 3108 18236 3120
rect 17267 3080 18236 3108
rect 17267 3077 17279 3080
rect 17221 3071 17279 3077
rect 18230 3068 18236 3080
rect 18288 3068 18294 3120
rect 18417 3111 18475 3117
rect 18417 3077 18429 3111
rect 18463 3108 18475 3111
rect 18598 3108 18604 3120
rect 18463 3080 18604 3108
rect 18463 3077 18475 3080
rect 18417 3071 18475 3077
rect 18598 3068 18604 3080
rect 18656 3068 18662 3120
rect 4939 3012 6914 3040
rect 8389 3043 8447 3049
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 14829 3043 14887 3049
rect 8389 3003 8447 3009
rect 12406 3012 14780 3040
rect 2406 2972 2412 2984
rect 2319 2944 2412 2972
rect 2406 2932 2412 2944
rect 2464 2972 2470 2984
rect 12253 2975 12311 2981
rect 2464 2944 6914 2972
rect 2464 2932 2470 2944
rect 6886 2904 6914 2944
rect 12253 2941 12265 2975
rect 12299 2972 12311 2975
rect 12406 2972 12434 3012
rect 12299 2944 12434 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 13998 2932 14004 2984
rect 14056 2972 14062 2984
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14056 2944 14565 2972
rect 14056 2932 14062 2944
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14752 2972 14780 3012
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 14875 3012 15761 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 18708 3040 18736 3148
rect 31754 3136 31760 3148
rect 31812 3136 31818 3188
rect 31938 3136 31944 3188
rect 31996 3176 32002 3188
rect 33226 3176 33232 3188
rect 31996 3148 33232 3176
rect 31996 3136 32002 3148
rect 33226 3136 33232 3148
rect 33284 3136 33290 3188
rect 33594 3136 33600 3188
rect 33652 3176 33658 3188
rect 34057 3179 34115 3185
rect 34057 3176 34069 3179
rect 33652 3148 34069 3176
rect 33652 3136 33658 3148
rect 34057 3145 34069 3148
rect 34103 3145 34115 3179
rect 34057 3139 34115 3145
rect 35897 3179 35955 3185
rect 35897 3145 35909 3179
rect 35943 3176 35955 3179
rect 36078 3176 36084 3188
rect 35943 3148 36084 3176
rect 35943 3145 35955 3148
rect 35897 3139 35955 3145
rect 36078 3136 36084 3148
rect 36136 3136 36142 3188
rect 36909 3179 36967 3185
rect 36909 3145 36921 3179
rect 36955 3145 36967 3179
rect 36909 3139 36967 3145
rect 18782 3068 18788 3120
rect 18840 3108 18846 3120
rect 18840 3080 20010 3108
rect 18840 3068 18846 3080
rect 21266 3068 21272 3120
rect 21324 3108 21330 3120
rect 21324 3080 21496 3108
rect 21324 3068 21330 3080
rect 21468 3052 21496 3080
rect 23290 3068 23296 3120
rect 23348 3068 23354 3120
rect 24029 3111 24087 3117
rect 24029 3077 24041 3111
rect 24075 3108 24087 3111
rect 24302 3108 24308 3120
rect 24075 3080 24308 3108
rect 24075 3077 24087 3080
rect 24029 3071 24087 3077
rect 24302 3068 24308 3080
rect 24360 3068 24366 3120
rect 24578 3108 24584 3120
rect 24539 3080 24584 3108
rect 24578 3068 24584 3080
rect 24636 3068 24642 3120
rect 24854 3068 24860 3120
rect 24912 3108 24918 3120
rect 24912 3080 25162 3108
rect 24912 3068 24918 3080
rect 26326 3068 26332 3120
rect 26384 3108 26390 3120
rect 26384 3080 26648 3108
rect 26384 3068 26390 3080
rect 18555 3012 18736 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 18932 3012 19165 3040
rect 18932 3000 18938 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 21450 3000 21456 3052
rect 21508 3040 21514 3052
rect 26620 3049 26648 3080
rect 27338 3068 27344 3120
rect 27396 3108 27402 3120
rect 27433 3111 27491 3117
rect 27433 3108 27445 3111
rect 27396 3080 27445 3108
rect 27396 3068 27402 3080
rect 27433 3077 27445 3080
rect 27479 3077 27491 3111
rect 28810 3108 28816 3120
rect 28658 3080 28816 3108
rect 27433 3071 27491 3077
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 29546 3068 29552 3120
rect 29604 3108 29610 3120
rect 29641 3111 29699 3117
rect 29641 3108 29653 3111
rect 29604 3080 29653 3108
rect 29604 3068 29610 3080
rect 29641 3077 29653 3080
rect 29687 3077 29699 3111
rect 31110 3108 31116 3120
rect 30958 3080 31116 3108
rect 29641 3071 29699 3077
rect 31110 3068 31116 3080
rect 31168 3068 31174 3120
rect 31294 3068 31300 3120
rect 31352 3108 31358 3120
rect 32585 3111 32643 3117
rect 32585 3108 32597 3111
rect 31352 3080 32597 3108
rect 31352 3068 31358 3080
rect 32585 3077 32597 3080
rect 32631 3077 32643 3111
rect 36630 3108 36636 3120
rect 33810 3080 36636 3108
rect 32585 3071 32643 3077
rect 36630 3068 36636 3080
rect 36688 3068 36694 3120
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21508 3012 22017 3040
rect 21508 3000 21514 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 26605 3043 26663 3049
rect 26605 3009 26617 3043
rect 26651 3040 26663 3043
rect 27062 3040 27068 3052
rect 26651 3012 27068 3040
rect 26651 3009 26663 3012
rect 26605 3003 26663 3009
rect 27062 3000 27068 3012
rect 27120 3040 27126 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 27120 3012 27169 3040
rect 27120 3000 27126 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 28718 3000 28724 3052
rect 28776 3040 28782 3052
rect 34793 3043 34851 3049
rect 28776 3012 29776 3040
rect 28776 3000 28782 3012
rect 15194 2972 15200 2984
rect 14752 2944 15200 2972
rect 14553 2935 14611 2941
rect 15194 2932 15200 2944
rect 15252 2972 15258 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15252 2944 15577 2972
rect 15252 2932 15258 2944
rect 15565 2941 15577 2944
rect 15611 2972 15623 2975
rect 15611 2944 16252 2972
rect 15611 2941 15623 2944
rect 15565 2935 15623 2941
rect 12710 2904 12716 2916
rect 6886 2876 12716 2904
rect 12710 2864 12716 2876
rect 12768 2864 12774 2916
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 16114 2904 16120 2916
rect 12851 2876 16120 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 16224 2904 16252 2944
rect 16298 2932 16304 2984
rect 16356 2972 16362 2984
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 16356 2944 21189 2972
rect 16356 2932 16362 2944
rect 21177 2941 21189 2944
rect 21223 2972 21235 2975
rect 22830 2972 22836 2984
rect 21223 2944 22836 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 22830 2932 22836 2944
rect 22888 2932 22894 2984
rect 26234 2932 26240 2984
rect 26292 2972 26298 2984
rect 26329 2975 26387 2981
rect 26329 2972 26341 2975
rect 26292 2944 26341 2972
rect 26292 2932 26298 2944
rect 26329 2941 26341 2944
rect 26375 2972 26387 2975
rect 26694 2972 26700 2984
rect 26375 2944 26700 2972
rect 26375 2941 26387 2944
rect 26329 2935 26387 2941
rect 26694 2932 26700 2944
rect 26752 2932 26758 2984
rect 28626 2972 28632 2984
rect 27264 2944 28632 2972
rect 16224 2876 16344 2904
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 7558 2796 7564 2848
rect 7616 2836 7622 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 7616 2808 8309 2836
rect 7616 2796 7622 2808
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 8297 2799 8355 2805
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 12434 2836 12440 2848
rect 11195 2808 12440 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 13906 2836 13912 2848
rect 13867 2808 13912 2836
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 16206 2836 16212 2848
rect 15528 2808 16212 2836
rect 15528 2796 15534 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 16316 2836 16344 2876
rect 17494 2864 17500 2916
rect 17552 2904 17558 2916
rect 17681 2907 17739 2913
rect 17681 2904 17693 2907
rect 17552 2876 17693 2904
rect 17552 2864 17558 2876
rect 17681 2873 17693 2876
rect 17727 2873 17739 2907
rect 17681 2867 17739 2873
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 17828 2876 19073 2904
rect 17828 2864 17834 2876
rect 19061 2873 19073 2876
rect 19107 2873 19119 2907
rect 19061 2867 19119 2873
rect 19260 2876 20208 2904
rect 19260 2836 19288 2876
rect 16316 2808 19288 2836
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 19705 2839 19763 2845
rect 19705 2836 19717 2839
rect 19484 2808 19717 2836
rect 19484 2796 19490 2808
rect 19705 2805 19717 2808
rect 19751 2805 19763 2839
rect 20180 2836 20208 2876
rect 24946 2864 24952 2916
rect 25004 2864 25010 2916
rect 27264 2904 27292 2944
rect 28626 2932 28632 2944
rect 28684 2972 28690 2984
rect 28902 2972 28908 2984
rect 28684 2944 28908 2972
rect 28684 2932 28690 2944
rect 28902 2932 28908 2944
rect 28960 2932 28966 2984
rect 29181 2975 29239 2981
rect 29181 2941 29193 2975
rect 29227 2972 29239 2975
rect 29638 2972 29644 2984
rect 29227 2944 29644 2972
rect 29227 2941 29239 2944
rect 29181 2935 29239 2941
rect 29638 2932 29644 2944
rect 29696 2932 29702 2984
rect 29748 2972 29776 3012
rect 34793 3009 34805 3043
rect 34839 3040 34851 3043
rect 35526 3040 35532 3052
rect 34839 3012 35532 3040
rect 34839 3009 34851 3012
rect 34793 3003 34851 3009
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 36354 3000 36360 3052
rect 36412 3040 36418 3052
rect 36725 3043 36783 3049
rect 36725 3040 36737 3043
rect 36412 3012 36737 3040
rect 36412 3000 36418 3012
rect 36725 3009 36737 3012
rect 36771 3009 36783 3043
rect 36924 3040 36952 3139
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 36924 3012 38025 3040
rect 36725 3003 36783 3009
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 31294 2972 31300 2984
rect 29748 2944 31300 2972
rect 31294 2932 31300 2944
rect 31352 2932 31358 2984
rect 31389 2975 31447 2981
rect 31389 2941 31401 2975
rect 31435 2972 31447 2975
rect 31665 2975 31723 2981
rect 31435 2944 31616 2972
rect 31435 2941 31447 2944
rect 31389 2935 31447 2941
rect 26620 2876 27292 2904
rect 21358 2836 21364 2848
rect 20180 2808 21364 2836
rect 19705 2799 19763 2805
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 22278 2845 22284 2848
rect 22268 2839 22284 2845
rect 22268 2805 22280 2839
rect 22268 2799 22284 2805
rect 22278 2796 22284 2799
rect 22336 2796 22342 2848
rect 24964 2836 24992 2864
rect 26620 2836 26648 2876
rect 28994 2864 29000 2916
rect 29052 2904 29058 2916
rect 30374 2904 30380 2916
rect 29052 2876 30380 2904
rect 29052 2864 29058 2876
rect 30374 2864 30380 2876
rect 30432 2864 30438 2916
rect 31588 2904 31616 2944
rect 31665 2941 31677 2975
rect 31711 2972 31723 2975
rect 32122 2972 32128 2984
rect 31711 2944 32128 2972
rect 31711 2941 31723 2944
rect 31665 2935 31723 2941
rect 32122 2932 32128 2944
rect 32180 2972 32186 2984
rect 32309 2975 32367 2981
rect 32309 2972 32321 2975
rect 32180 2944 32321 2972
rect 32180 2932 32186 2944
rect 32309 2941 32321 2944
rect 32355 2941 32367 2975
rect 35342 2972 35348 2984
rect 32309 2935 32367 2941
rect 32416 2944 35348 2972
rect 31754 2904 31760 2916
rect 31588 2876 31760 2904
rect 31754 2864 31760 2876
rect 31812 2864 31818 2916
rect 31846 2864 31852 2916
rect 31904 2904 31910 2916
rect 32416 2904 32444 2944
rect 35342 2932 35348 2944
rect 35400 2932 35406 2984
rect 35253 2907 35311 2913
rect 35253 2904 35265 2907
rect 31904 2876 32444 2904
rect 33612 2876 35265 2904
rect 31904 2864 31910 2876
rect 24964 2808 26648 2836
rect 26694 2796 26700 2848
rect 26752 2836 26758 2848
rect 33612 2836 33640 2876
rect 35253 2873 35265 2876
rect 35299 2873 35311 2907
rect 35253 2867 35311 2873
rect 26752 2808 33640 2836
rect 26752 2796 26758 2808
rect 34146 2796 34152 2848
rect 34204 2836 34210 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 34204 2808 34621 2836
rect 34204 2796 34210 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 37550 2836 37556 2848
rect 37511 2808 37556 2836
rect 34609 2799 34667 2805
rect 37550 2796 37556 2808
rect 37608 2796 37614 2848
rect 38197 2839 38255 2845
rect 38197 2805 38209 2839
rect 38243 2836 38255 2839
rect 38286 2836 38292 2848
rect 38243 2808 38292 2836
rect 38243 2805 38255 2808
rect 38197 2799 38255 2805
rect 38286 2796 38292 2808
rect 38344 2796 38350 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 10042 2632 10048 2644
rect 9955 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2632 10106 2644
rect 12250 2632 12256 2644
rect 10100 2604 12256 2632
rect 10100 2592 10106 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12529 2635 12587 2641
rect 12529 2601 12541 2635
rect 12575 2632 12587 2635
rect 13906 2632 13912 2644
rect 12575 2604 13912 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 17770 2632 17776 2644
rect 14384 2604 17776 2632
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 72 2536 2421 2564
rect 72 2524 78 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 8662 2564 8668 2576
rect 2409 2527 2467 2533
rect 2608 2536 8668 2564
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2406 2428 2412 2440
rect 1903 2400 2412 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 2608 2437 2636 2536
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 12986 2564 12992 2576
rect 9447 2536 12992 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 14277 2567 14335 2573
rect 14277 2564 14289 2567
rect 13688 2536 14289 2564
rect 13688 2524 13694 2536
rect 14277 2533 14289 2536
rect 14323 2533 14335 2567
rect 14277 2527 14335 2533
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4614 2496 4620 2508
rect 4295 2468 4620 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 9214 2496 9220 2508
rect 5552 2468 9220 2496
rect 5552 2437 5580 2468
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 14384 2496 14412 2604
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18049 2635 18107 2641
rect 18049 2601 18061 2635
rect 18095 2632 18107 2635
rect 19334 2632 19340 2644
rect 18095 2604 19340 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 28534 2632 28540 2644
rect 19484 2604 28540 2632
rect 19484 2592 19490 2604
rect 28534 2592 28540 2604
rect 28592 2592 28598 2644
rect 28626 2592 28632 2644
rect 28684 2632 28690 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 28684 2604 28917 2632
rect 28684 2592 28690 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 33410 2632 33416 2644
rect 28905 2595 28963 2601
rect 30024 2604 33416 2632
rect 16850 2524 16856 2576
rect 16908 2524 16914 2576
rect 23382 2524 23388 2576
rect 23440 2564 23446 2576
rect 23440 2536 24808 2564
rect 23440 2524 23446 2536
rect 16868 2496 16896 2524
rect 18874 2496 18880 2508
rect 11992 2468 14412 2496
rect 15304 2468 16896 2496
rect 17972 2468 18880 2496
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 2593 2391 2651 2397
rect 3344 2400 3985 2428
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3344 2301 3372 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 7558 2428 7564 2440
rect 6871 2400 7564 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 11992 2437 12020 2468
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2428 9919 2431
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 9907 2400 10517 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 12492 2400 13553 2428
rect 12492 2388 12498 2400
rect 13541 2397 13553 2400
rect 13587 2428 13599 2431
rect 14826 2428 14832 2440
rect 13587 2400 14832 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 11149 2363 11207 2369
rect 11149 2329 11161 2363
rect 11195 2360 11207 2363
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 11195 2332 14473 2360
rect 11195 2329 11207 2332
rect 11149 2323 11207 2329
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 4580 2264 5365 2292
rect 4580 2252 4586 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2292 8539 2295
rect 9232 2292 9260 2323
rect 13556 2304 13584 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 15304 2360 15332 2468
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 17972 2437 18000 2468
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 21450 2496 21456 2508
rect 21411 2468 21456 2496
rect 21450 2456 21456 2468
rect 21508 2496 21514 2508
rect 22005 2499 22063 2505
rect 22005 2496 22017 2499
rect 21508 2468 22017 2496
rect 21508 2456 21514 2468
rect 22005 2465 22017 2468
rect 22051 2496 22063 2499
rect 24670 2496 24676 2508
rect 22051 2468 24676 2496
rect 22051 2465 22063 2468
rect 22005 2459 22063 2465
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 24780 2496 24808 2536
rect 25958 2524 25964 2576
rect 26016 2564 26022 2576
rect 26878 2564 26884 2576
rect 26016 2536 26884 2564
rect 26016 2524 26022 2536
rect 26878 2524 26884 2536
rect 26936 2524 26942 2576
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 24780 2468 27445 2496
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 28902 2456 28908 2508
rect 28960 2496 28966 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 28960 2468 29745 2496
rect 28960 2456 28966 2468
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 29733 2459 29791 2465
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16316 2400 16865 2428
rect 14461 2323 14519 2329
rect 15120 2332 15332 2360
rect 8527 2264 9260 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 13078 2292 13084 2304
rect 13039 2264 13084 2292
rect 11793 2255 11851 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 13538 2252 13544 2304
rect 13596 2252 13602 2304
rect 13725 2295 13783 2301
rect 13725 2261 13737 2295
rect 13771 2292 13783 2295
rect 15120 2292 15148 2332
rect 15286 2292 15292 2304
rect 13771 2264 15148 2292
rect 15247 2264 15292 2292
rect 13771 2261 13783 2264
rect 13725 2255 13783 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 16316 2301 16344 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17957 2431 18015 2437
rect 17957 2397 17969 2431
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18564 2400 18613 2428
rect 18564 2388 18570 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 30024 2428 30052 2604
rect 33410 2592 33416 2604
rect 33468 2592 33474 2644
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 34422 2632 34428 2644
rect 33744 2604 34428 2632
rect 33744 2592 33750 2604
rect 34422 2592 34428 2604
rect 34480 2592 34486 2644
rect 37550 2592 37556 2644
rect 37608 2632 37614 2644
rect 38194 2632 38200 2644
rect 37608 2604 38200 2632
rect 37608 2592 37614 2604
rect 38194 2592 38200 2604
rect 38252 2592 38258 2644
rect 32674 2564 32680 2576
rect 31404 2536 32680 2564
rect 31404 2496 31432 2536
rect 32674 2524 32680 2536
rect 32732 2524 32738 2576
rect 34238 2564 34244 2576
rect 34072 2536 34244 2564
rect 28566 2400 30052 2428
rect 30116 2468 31432 2496
rect 31481 2499 31539 2505
rect 30116 2414 30144 2468
rect 31481 2465 31493 2499
rect 31527 2496 31539 2499
rect 32122 2496 32128 2508
rect 31527 2468 32128 2496
rect 31527 2465 31539 2468
rect 31481 2459 31539 2465
rect 32122 2456 32128 2468
rect 32180 2496 32186 2508
rect 34072 2505 34100 2536
rect 34238 2524 34244 2536
rect 34296 2524 34302 2576
rect 37090 2564 37096 2576
rect 35866 2536 37096 2564
rect 34057 2499 34115 2505
rect 34057 2496 34069 2499
rect 32180 2468 34069 2496
rect 32180 2456 32186 2468
rect 34057 2465 34069 2468
rect 34103 2465 34115 2499
rect 35866 2496 35894 2536
rect 37090 2524 37096 2536
rect 37148 2524 37154 2576
rect 34057 2459 34115 2465
rect 34256 2468 35894 2496
rect 27157 2391 27215 2397
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 16448 2332 19334 2360
rect 16448 2320 16454 2332
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18748 2264 18797 2292
rect 18748 2252 18754 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 19306 2292 19334 2332
rect 20162 2320 20168 2372
rect 20220 2320 20226 2372
rect 21174 2360 21180 2372
rect 21135 2332 21180 2360
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 21266 2320 21272 2372
rect 21324 2360 21330 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21324 2332 22293 2360
rect 21324 2320 21330 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 22738 2320 22744 2372
rect 22796 2320 22802 2372
rect 24946 2360 24952 2372
rect 24907 2332 24952 2360
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 26174 2332 27844 2360
rect 19705 2295 19763 2301
rect 19705 2292 19717 2295
rect 19306 2264 19717 2292
rect 18785 2255 18843 2261
rect 19705 2261 19717 2264
rect 19751 2292 19763 2295
rect 21910 2292 21916 2304
rect 19751 2264 21916 2292
rect 19751 2261 19763 2264
rect 19705 2255 19763 2261
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 22462 2252 22468 2304
rect 22520 2292 22526 2304
rect 23753 2295 23811 2301
rect 23753 2292 23765 2295
rect 22520 2264 23765 2292
rect 22520 2252 22526 2264
rect 23753 2261 23765 2264
rect 23799 2292 23811 2295
rect 25958 2292 25964 2304
rect 23799 2264 25964 2292
rect 23799 2261 23811 2264
rect 23753 2255 23811 2261
rect 25958 2252 25964 2264
rect 26016 2252 26022 2304
rect 26421 2295 26479 2301
rect 26421 2261 26433 2295
rect 26467 2292 26479 2295
rect 27614 2292 27620 2304
rect 26467 2264 27620 2292
rect 26467 2261 26479 2264
rect 26421 2255 26479 2261
rect 27614 2252 27620 2264
rect 27672 2252 27678 2304
rect 27816 2292 27844 2332
rect 31110 2320 31116 2372
rect 31168 2360 31174 2372
rect 31205 2363 31263 2369
rect 31205 2360 31217 2363
rect 31168 2332 31217 2360
rect 31168 2320 31174 2332
rect 31205 2329 31217 2332
rect 31251 2329 31263 2363
rect 31205 2323 31263 2329
rect 31312 2332 32444 2360
rect 29270 2292 29276 2304
rect 27816 2264 29276 2292
rect 29270 2252 29276 2264
rect 29328 2252 29334 2304
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 31312 2292 31340 2332
rect 30340 2264 31340 2292
rect 30340 2252 30346 2264
rect 31386 2252 31392 2304
rect 31444 2292 31450 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 31444 2264 32321 2292
rect 31444 2252 31450 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32416 2292 32444 2332
rect 32766 2320 32772 2372
rect 32824 2320 32830 2372
rect 33781 2363 33839 2369
rect 33781 2329 33793 2363
rect 33827 2360 33839 2363
rect 34256 2360 34284 2468
rect 34330 2388 34336 2440
rect 34388 2428 34394 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34388 2400 34897 2428
rect 34388 2388 34394 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35710 2428 35716 2440
rect 35492 2400 35716 2428
rect 35492 2388 35498 2400
rect 35710 2388 35716 2400
rect 35768 2428 35774 2440
rect 35805 2431 35863 2437
rect 35805 2428 35817 2431
rect 35768 2400 35817 2428
rect 35768 2388 35774 2400
rect 35805 2397 35817 2400
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 36633 2431 36691 2437
rect 36633 2397 36645 2431
rect 36679 2397 36691 2431
rect 37458 2428 37464 2440
rect 37419 2400 37464 2428
rect 36633 2391 36691 2397
rect 33827 2332 34284 2360
rect 33827 2329 33839 2332
rect 33781 2323 33839 2329
rect 34422 2320 34428 2372
rect 34480 2360 34486 2372
rect 36648 2360 36676 2391
rect 37458 2388 37464 2400
rect 37516 2388 37522 2440
rect 34480 2332 36676 2360
rect 34480 2320 34486 2332
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 32416 2264 35081 2292
rect 32309 2255 32367 2261
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35710 2292 35716 2304
rect 35671 2264 35716 2292
rect 35069 2255 35127 2261
rect 35710 2252 35716 2264
rect 35768 2252 35774 2304
rect 36817 2295 36875 2301
rect 36817 2261 36829 2295
rect 36863 2292 36875 2295
rect 37182 2292 37188 2304
rect 36863 2264 37188 2292
rect 36863 2261 36875 2264
rect 36817 2255 36875 2261
rect 37182 2252 37188 2264
rect 37240 2252 37246 2304
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37424 2264 37657 2292
rect 37424 2252 37430 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 15286 2048 15292 2100
rect 15344 2088 15350 2100
rect 24854 2088 24860 2100
rect 15344 2060 24860 2088
rect 15344 2048 15350 2060
rect 24854 2048 24860 2060
rect 24912 2048 24918 2100
rect 25866 2048 25872 2100
rect 25924 2088 25930 2100
rect 35710 2088 35716 2100
rect 25924 2060 35716 2088
rect 25924 2048 25930 2060
rect 35710 2048 35716 2060
rect 35768 2048 35774 2100
rect 16114 1980 16120 2032
rect 16172 2020 16178 2032
rect 19426 2020 19432 2032
rect 16172 1992 19432 2020
rect 16172 1980 16178 1992
rect 19426 1980 19432 1992
rect 19484 1980 19490 2032
rect 27614 1980 27620 2032
rect 27672 2020 27678 2032
rect 30926 2020 30932 2032
rect 27672 1992 30932 2020
rect 27672 1980 27678 1992
rect 30926 1980 30932 1992
rect 30984 1980 30990 2032
rect 16206 1912 16212 1964
rect 16264 1952 16270 1964
rect 21174 1952 21180 1964
rect 16264 1924 21180 1952
rect 16264 1912 16270 1924
rect 21174 1912 21180 1924
rect 21232 1952 21238 1964
rect 21232 1924 22094 1952
rect 21232 1912 21238 1924
rect 13078 1844 13084 1896
rect 13136 1884 13142 1896
rect 21082 1884 21088 1896
rect 13136 1856 21088 1884
rect 13136 1844 13142 1856
rect 21082 1844 21088 1856
rect 21140 1844 21146 1896
rect 22066 1884 22094 1924
rect 28534 1912 28540 1964
rect 28592 1952 28598 1964
rect 38010 1952 38016 1964
rect 28592 1924 38016 1952
rect 28592 1912 28598 1924
rect 38010 1912 38016 1924
rect 38068 1912 38074 1964
rect 23198 1884 23204 1896
rect 22066 1856 23204 1884
rect 23198 1844 23204 1856
rect 23256 1844 23262 1896
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 18052 37408 18104 37460
rect 14556 37340 14608 37392
rect 1768 37204 1820 37256
rect 4068 37204 4120 37256
rect 7288 37204 7340 37256
rect 7748 37204 7800 37256
rect 9680 37204 9732 37256
rect 11980 37247 12032 37256
rect 11980 37213 11989 37247
rect 11989 37213 12023 37247
rect 12023 37213 12032 37247
rect 14832 37272 14884 37324
rect 16672 37272 16724 37324
rect 16764 37272 16816 37324
rect 13268 37247 13320 37256
rect 11980 37204 12032 37213
rect 13268 37213 13277 37247
rect 13277 37213 13311 37247
rect 13311 37213 13320 37247
rect 13268 37204 13320 37213
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 18052 37204 18104 37256
rect 20352 37247 20404 37256
rect 20352 37213 20361 37247
rect 20361 37213 20395 37247
rect 20395 37213 20404 37247
rect 21916 37272 21968 37324
rect 35440 37272 35492 37324
rect 38292 37315 38344 37324
rect 38292 37281 38301 37315
rect 38301 37281 38335 37315
rect 38335 37281 38344 37315
rect 38292 37272 38344 37281
rect 22284 37247 22336 37256
rect 20352 37204 20404 37213
rect 22284 37213 22293 37247
rect 22293 37213 22327 37247
rect 22327 37213 22336 37247
rect 22284 37204 22336 37213
rect 22560 37204 22612 37256
rect 23388 37204 23440 37256
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 28448 37247 28500 37256
rect 28448 37213 28457 37247
rect 28457 37213 28491 37247
rect 28491 37213 28500 37247
rect 28448 37204 28500 37213
rect 30472 37204 30524 37256
rect 32588 37247 32640 37256
rect 32588 37213 32597 37247
rect 32597 37213 32631 37247
rect 32631 37213 32640 37247
rect 32588 37204 32640 37213
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 35808 37247 35860 37256
rect 35808 37213 35817 37247
rect 35817 37213 35851 37247
rect 35851 37213 35860 37247
rect 35808 37204 35860 37213
rect 37832 37204 37884 37256
rect 1308 37068 1360 37120
rect 2780 37111 2832 37120
rect 2780 37077 2789 37111
rect 2789 37077 2823 37111
rect 2823 37077 2832 37111
rect 2780 37068 2832 37077
rect 4620 37068 4672 37120
rect 5448 37111 5500 37120
rect 5448 37077 5457 37111
rect 5457 37077 5491 37111
rect 5491 37077 5500 37111
rect 5448 37068 5500 37077
rect 6460 37068 6512 37120
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 9956 37111 10008 37120
rect 9956 37077 9965 37111
rect 9965 37077 9999 37111
rect 9999 37077 10008 37111
rect 9956 37068 10008 37077
rect 11612 37068 11664 37120
rect 12900 37068 12952 37120
rect 19984 37068 20036 37120
rect 23204 37068 23256 37120
rect 25136 37068 25188 37120
rect 27068 37068 27120 37120
rect 28356 37068 28408 37120
rect 30380 37068 30432 37120
rect 32220 37068 32272 37120
rect 33508 37068 33560 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 5448 36864 5500 36916
rect 21180 36864 21232 36916
rect 22560 36907 22612 36916
rect 22560 36873 22569 36907
rect 22569 36873 22603 36907
rect 22603 36873 22612 36907
rect 22560 36864 22612 36873
rect 33600 36864 33652 36916
rect 37372 36864 37424 36916
rect 38292 36907 38344 36916
rect 38292 36873 38301 36907
rect 38301 36873 38335 36907
rect 38335 36873 38344 36907
rect 38292 36864 38344 36873
rect 2872 36796 2924 36848
rect 22284 36796 22336 36848
rect 2964 36728 3016 36780
rect 15200 36728 15252 36780
rect 15936 36728 15988 36780
rect 23112 36728 23164 36780
rect 36820 36728 36872 36780
rect 2044 36592 2096 36644
rect 17500 36592 17552 36644
rect 7288 36524 7340 36576
rect 13268 36524 13320 36576
rect 23112 36567 23164 36576
rect 23112 36533 23121 36567
rect 23121 36533 23155 36567
rect 23155 36533 23164 36567
rect 23112 36524 23164 36533
rect 36820 36567 36872 36576
rect 36820 36533 36829 36567
rect 36829 36533 36863 36567
rect 36863 36533 36872 36567
rect 36820 36524 36872 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2872 36320 2924 36372
rect 23112 36320 23164 36372
rect 35808 36320 35860 36372
rect 37188 36320 37240 36372
rect 38660 36320 38712 36372
rect 1860 36159 1912 36168
rect 1860 36125 1869 36159
rect 1869 36125 1903 36159
rect 1903 36125 1912 36159
rect 1860 36116 1912 36125
rect 38016 36159 38068 36168
rect 38016 36125 38025 36159
rect 38025 36125 38059 36159
rect 38059 36125 38068 36159
rect 38016 36116 38068 36125
rect 1676 36023 1728 36032
rect 1676 35989 1685 36023
rect 1685 35989 1719 36023
rect 1719 35989 1728 36023
rect 1676 35980 1728 35989
rect 36728 36023 36780 36032
rect 36728 35989 36737 36023
rect 36737 35989 36771 36023
rect 36771 35989 36780 36023
rect 36728 35980 36780 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 37464 35615 37516 35624
rect 37464 35581 37473 35615
rect 37473 35581 37507 35615
rect 37507 35581 37516 35615
rect 37464 35572 37516 35581
rect 37740 35615 37792 35624
rect 37740 35581 37749 35615
rect 37749 35581 37783 35615
rect 37783 35581 37792 35615
rect 37740 35572 37792 35581
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 23388 35232 23440 35284
rect 30472 35232 30524 35284
rect 38016 35275 38068 35284
rect 38016 35241 38025 35275
rect 38025 35241 38059 35275
rect 38059 35241 38068 35275
rect 38016 35232 38068 35241
rect 21088 35028 21140 35080
rect 29644 35028 29696 35080
rect 30748 35028 30800 35080
rect 37740 35028 37792 35080
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1860 34688 1912 34740
rect 2136 34552 2188 34604
rect 18144 34484 18196 34536
rect 1676 34391 1728 34400
rect 1676 34357 1685 34391
rect 1685 34357 1719 34391
rect 1719 34357 1728 34391
rect 1676 34348 1728 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2136 33804 2188 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 15844 33260 15896 33312
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 32588 32555 32640 32564
rect 32588 32521 32597 32555
rect 32597 32521 32631 32555
rect 32631 32521 32640 32555
rect 32588 32512 32640 32521
rect 1584 32376 1636 32428
rect 27988 32376 28040 32428
rect 29644 32308 29696 32360
rect 38292 32351 38344 32360
rect 38292 32317 38301 32351
rect 38301 32317 38335 32351
rect 38335 32317 38344 32351
rect 38292 32308 38344 32317
rect 21088 32172 21140 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 38292 32011 38344 32020
rect 38292 31977 38301 32011
rect 38301 31977 38335 32011
rect 38335 31977 38344 32011
rect 38292 31968 38344 31977
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 1860 30651 1912 30660
rect 1860 30617 1869 30651
rect 1869 30617 1903 30651
rect 1903 30617 1912 30651
rect 1860 30608 1912 30617
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 1676 30379 1728 30388
rect 1676 30345 1685 30379
rect 1685 30345 1719 30379
rect 1719 30345 1728 30379
rect 1676 30336 1728 30345
rect 38016 30243 38068 30252
rect 4068 30064 4120 30116
rect 38016 30209 38025 30243
rect 38025 30209 38059 30243
rect 38059 30209 38068 30243
rect 38016 30200 38068 30209
rect 12440 30039 12492 30048
rect 12440 30005 12449 30039
rect 12449 30005 12483 30039
rect 12483 30005 12492 30039
rect 12440 29996 12492 30005
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 22192 29792 22244 29844
rect 23112 29792 23164 29844
rect 38016 29835 38068 29844
rect 38016 29801 38025 29835
rect 38025 29801 38059 29835
rect 38059 29801 38068 29835
rect 38016 29792 38068 29801
rect 37832 29631 37884 29640
rect 37832 29597 37841 29631
rect 37841 29597 37875 29631
rect 37875 29597 37884 29631
rect 37832 29588 37884 29597
rect 20720 29520 20772 29572
rect 36728 29452 36780 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1584 29112 1636 29164
rect 22192 29155 22244 29164
rect 22192 29121 22201 29155
rect 22201 29121 22235 29155
rect 22235 29121 22244 29155
rect 22192 29112 22244 29121
rect 22284 29112 22336 29164
rect 12440 29044 12492 29096
rect 23756 29044 23808 29096
rect 20720 28976 20772 29028
rect 22192 28976 22244 29028
rect 23572 28976 23624 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 21180 28747 21232 28756
rect 21180 28713 21189 28747
rect 21189 28713 21223 28747
rect 21223 28713 21232 28747
rect 21180 28704 21232 28713
rect 1584 28679 1636 28688
rect 1584 28645 1593 28679
rect 1593 28645 1627 28679
rect 1627 28645 1636 28679
rect 1584 28636 1636 28645
rect 23388 28364 23440 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 15936 28067 15988 28076
rect 15936 28033 15945 28067
rect 15945 28033 15979 28067
rect 15979 28033 15988 28067
rect 15936 28024 15988 28033
rect 16120 27820 16172 27872
rect 20628 27820 20680 27872
rect 38200 27931 38252 27940
rect 38200 27897 38209 27931
rect 38209 27897 38243 27931
rect 38243 27897 38252 27931
rect 38200 27888 38252 27897
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 23388 27616 23440 27668
rect 38016 27616 38068 27668
rect 30748 27455 30800 27464
rect 30748 27421 30757 27455
rect 30757 27421 30791 27455
rect 30791 27421 30800 27455
rect 30748 27412 30800 27421
rect 27804 27276 27856 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 20628 27072 20680 27124
rect 38016 27047 38068 27056
rect 38016 27013 38025 27047
rect 38025 27013 38059 27047
rect 38059 27013 38068 27047
rect 38016 27004 38068 27013
rect 6828 26936 6880 26988
rect 2044 26868 2096 26920
rect 20076 26979 20128 26988
rect 20076 26945 20085 26979
rect 20085 26945 20119 26979
rect 20119 26945 20128 26979
rect 20076 26936 20128 26945
rect 38200 26979 38252 26988
rect 38200 26945 38209 26979
rect 38209 26945 38243 26979
rect 38243 26945 38252 26979
rect 38200 26936 38252 26945
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 1768 26027 1820 26036
rect 1768 25993 1777 26027
rect 1777 25993 1811 26027
rect 1811 25993 1820 26027
rect 1768 25984 1820 25993
rect 2044 25848 2096 25900
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 21088 25440 21140 25492
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 1952 25236 2004 25288
rect 21088 25236 21140 25288
rect 29644 25440 29696 25492
rect 37832 25236 37884 25288
rect 20536 25100 20588 25152
rect 26700 25100 26752 25152
rect 32036 25143 32088 25152
rect 32036 25109 32045 25143
rect 32045 25109 32079 25143
rect 32079 25109 32088 25143
rect 32036 25100 32088 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 38016 24803 38068 24812
rect 38016 24769 38025 24803
rect 38025 24769 38059 24803
rect 38059 24769 38068 24803
rect 38016 24760 38068 24769
rect 27160 24624 27212 24676
rect 29920 24556 29972 24608
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 11980 24080 12032 24132
rect 21272 24080 21324 24132
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 2872 23672 2924 23724
rect 1676 23511 1728 23520
rect 1676 23477 1685 23511
rect 1685 23477 1719 23511
rect 1719 23477 1728 23511
rect 1676 23468 1728 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 20076 22720 20128 22772
rect 34060 22584 34112 22636
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 20904 22380 20956 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 20812 21632 20864 21684
rect 1768 21496 1820 21548
rect 37464 21496 37516 21548
rect 13268 21360 13320 21412
rect 25136 21360 25188 21412
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 22836 21292 22888 21344
rect 37464 21335 37516 21344
rect 37464 21301 37473 21335
rect 37473 21301 37507 21335
rect 37507 21301 37516 21335
rect 37464 21292 37516 21301
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1768 21131 1820 21140
rect 1768 21097 1777 21131
rect 1777 21097 1811 21131
rect 1811 21097 1820 21131
rect 1768 21088 1820 21097
rect 6828 21088 6880 21140
rect 1952 20927 2004 20936
rect 1952 20893 1961 20927
rect 1961 20893 1995 20927
rect 1995 20893 2004 20927
rect 1952 20884 2004 20893
rect 8944 20748 8996 20800
rect 13452 20748 13504 20800
rect 14464 20748 14516 20800
rect 25320 20748 25372 20800
rect 38016 20748 38068 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 23388 20544 23440 20596
rect 21088 20408 21140 20460
rect 23204 20340 23256 20392
rect 25044 20272 25096 20324
rect 27528 20272 27580 20324
rect 1860 20204 1912 20256
rect 19984 20204 20036 20256
rect 22468 20204 22520 20256
rect 24400 20204 24452 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 28448 20000 28500 20052
rect 20904 19864 20956 19916
rect 26884 19864 26936 19916
rect 37464 19864 37516 19916
rect 4712 19796 4764 19848
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 22100 19771 22152 19780
rect 22100 19737 22109 19771
rect 22109 19737 22143 19771
rect 22143 19737 22152 19771
rect 22652 19771 22704 19780
rect 22100 19728 22152 19737
rect 22652 19737 22661 19771
rect 22661 19737 22695 19771
rect 22695 19737 22704 19771
rect 22652 19728 22704 19737
rect 26148 19796 26200 19848
rect 26792 19728 26844 19780
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 19340 19660 19392 19712
rect 20260 19703 20312 19712
rect 20260 19669 20269 19703
rect 20269 19669 20303 19703
rect 20303 19669 20312 19703
rect 20260 19660 20312 19669
rect 20720 19660 20772 19712
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 24124 19660 24176 19712
rect 25596 19660 25648 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 26884 19456 26936 19508
rect 34060 19499 34112 19508
rect 34060 19465 34069 19499
rect 34069 19465 34103 19499
rect 34103 19465 34112 19499
rect 34060 19456 34112 19465
rect 18696 19388 18748 19440
rect 20536 19388 20588 19440
rect 20812 19431 20864 19440
rect 20812 19397 20821 19431
rect 20821 19397 20855 19431
rect 20855 19397 20864 19431
rect 20812 19388 20864 19397
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 21732 19320 21784 19372
rect 22468 19431 22520 19440
rect 22468 19397 22477 19431
rect 22477 19397 22511 19431
rect 22511 19397 22520 19431
rect 22468 19388 22520 19397
rect 23756 19388 23808 19440
rect 25872 19388 25924 19440
rect 26056 19431 26108 19440
rect 26056 19397 26065 19431
rect 26065 19397 26099 19431
rect 26099 19397 26108 19431
rect 26056 19388 26108 19397
rect 26700 19388 26752 19440
rect 29184 19320 29236 19372
rect 38016 19363 38068 19372
rect 38016 19329 38025 19363
rect 38025 19329 38059 19363
rect 38059 19329 38068 19363
rect 38016 19320 38068 19329
rect 20904 19252 20956 19304
rect 24768 19252 24820 19304
rect 25412 19252 25464 19304
rect 20904 19116 20956 19168
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4712 18955 4764 18964
rect 4712 18921 4721 18955
rect 4721 18921 4755 18955
rect 4755 18921 4764 18955
rect 4712 18912 4764 18921
rect 20812 18912 20864 18964
rect 22100 18912 22152 18964
rect 25504 18912 25556 18964
rect 30932 18912 30984 18964
rect 18972 18708 19024 18760
rect 20260 18819 20312 18828
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 22192 18776 22244 18828
rect 22376 18819 22428 18828
rect 22376 18785 22385 18819
rect 22385 18785 22419 18819
rect 22419 18785 22428 18819
rect 22376 18776 22428 18785
rect 21088 18708 21140 18760
rect 20720 18640 20772 18692
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 8024 18572 8076 18624
rect 12900 18572 12952 18624
rect 19432 18572 19484 18624
rect 23664 18708 23716 18760
rect 24032 18844 24084 18896
rect 27160 18844 27212 18896
rect 24124 18708 24176 18760
rect 22192 18683 22244 18692
rect 22192 18649 22201 18683
rect 22201 18649 22235 18683
rect 22235 18649 22244 18683
rect 22192 18640 22244 18649
rect 22560 18572 22612 18624
rect 22652 18572 22704 18624
rect 23388 18572 23440 18624
rect 23756 18640 23808 18692
rect 25504 18683 25556 18692
rect 25504 18649 25513 18683
rect 25513 18649 25547 18683
rect 25547 18649 25556 18683
rect 25504 18640 25556 18649
rect 26700 18776 26752 18828
rect 25688 18572 25740 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 15844 18411 15896 18420
rect 15844 18377 15853 18411
rect 15853 18377 15887 18411
rect 15887 18377 15896 18411
rect 15844 18368 15896 18377
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 1584 18232 1636 18284
rect 1952 18232 2004 18284
rect 17684 18300 17736 18352
rect 19708 18368 19760 18420
rect 20536 18368 20588 18420
rect 22192 18368 22244 18420
rect 19524 18300 19576 18352
rect 25780 18368 25832 18420
rect 38016 18368 38068 18420
rect 15476 18232 15528 18284
rect 21364 18232 21416 18284
rect 22192 18232 22244 18284
rect 16488 18096 16540 18148
rect 19340 18164 19392 18216
rect 19708 18164 19760 18216
rect 22376 18164 22428 18216
rect 19984 18096 20036 18148
rect 21548 18096 21600 18148
rect 23756 18343 23808 18352
rect 23756 18309 23765 18343
rect 23765 18309 23799 18343
rect 23799 18309 23808 18343
rect 23756 18300 23808 18309
rect 25596 18343 25648 18352
rect 25596 18309 25605 18343
rect 25605 18309 25639 18343
rect 25639 18309 25648 18343
rect 25596 18300 25648 18309
rect 25688 18343 25740 18352
rect 25688 18309 25697 18343
rect 25697 18309 25731 18343
rect 25731 18309 25740 18343
rect 27160 18343 27212 18352
rect 25688 18300 25740 18309
rect 27160 18309 27169 18343
rect 27169 18309 27203 18343
rect 27203 18309 27212 18343
rect 27160 18300 27212 18309
rect 27528 18300 27580 18352
rect 27804 18343 27856 18352
rect 27804 18309 27813 18343
rect 27813 18309 27847 18343
rect 27847 18309 27856 18343
rect 27804 18300 27856 18309
rect 24400 18275 24452 18284
rect 24400 18241 24409 18275
rect 24409 18241 24443 18275
rect 24443 18241 24452 18275
rect 24400 18232 24452 18241
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 24860 18164 24912 18216
rect 23204 18096 23256 18148
rect 23664 18096 23716 18148
rect 28908 18232 28960 18284
rect 22468 18028 22520 18080
rect 23756 18028 23808 18080
rect 24400 18028 24452 18080
rect 26608 18096 26660 18148
rect 26332 18071 26384 18080
rect 26332 18037 26341 18071
rect 26341 18037 26375 18071
rect 26375 18037 26384 18071
rect 26332 18028 26384 18037
rect 29000 18028 29052 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 20904 17824 20956 17876
rect 23296 17824 23348 17876
rect 25964 17824 26016 17876
rect 26056 17824 26108 17876
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 19156 17756 19208 17808
rect 21732 17756 21784 17808
rect 22192 17756 22244 17808
rect 22744 17756 22796 17808
rect 24768 17756 24820 17808
rect 21364 17688 21416 17740
rect 27804 17756 27856 17808
rect 26516 17688 26568 17740
rect 19156 17620 19208 17672
rect 19984 17620 20036 17672
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 23664 17663 23716 17672
rect 23664 17629 23673 17663
rect 23673 17629 23707 17663
rect 23707 17629 23716 17663
rect 23664 17620 23716 17629
rect 23940 17620 23992 17672
rect 24308 17620 24360 17672
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 26884 17620 26936 17672
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 19432 17552 19484 17604
rect 20996 17552 21048 17604
rect 22376 17595 22428 17604
rect 22376 17561 22385 17595
rect 22385 17561 22419 17595
rect 22419 17561 22428 17595
rect 22376 17552 22428 17561
rect 18512 17484 18564 17536
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 24952 17484 25004 17536
rect 26240 17552 26292 17604
rect 26332 17484 26384 17536
rect 27620 17484 27672 17536
rect 28448 17527 28500 17536
rect 28448 17493 28457 17527
rect 28457 17493 28491 17527
rect 28491 17493 28500 17527
rect 28448 17484 28500 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 17408 17255 17460 17264
rect 17408 17221 17417 17255
rect 17417 17221 17451 17255
rect 17451 17221 17460 17255
rect 17408 17212 17460 17221
rect 18696 17280 18748 17332
rect 18512 17255 18564 17264
rect 18512 17221 18521 17255
rect 18521 17221 18555 17255
rect 18555 17221 18564 17255
rect 18512 17212 18564 17221
rect 20904 17212 20956 17264
rect 20260 17187 20312 17196
rect 20260 17153 20269 17187
rect 20269 17153 20303 17187
rect 20303 17153 20312 17187
rect 23296 17280 23348 17332
rect 23480 17280 23532 17332
rect 21180 17212 21232 17264
rect 23756 17255 23808 17264
rect 23756 17221 23765 17255
rect 23765 17221 23799 17255
rect 23799 17221 23808 17255
rect 23756 17212 23808 17221
rect 24952 17255 25004 17264
rect 24952 17221 24961 17255
rect 24961 17221 24995 17255
rect 24995 17221 25004 17255
rect 24952 17212 25004 17221
rect 25044 17255 25096 17264
rect 25044 17221 25053 17255
rect 25053 17221 25087 17255
rect 25087 17221 25096 17255
rect 25044 17212 25096 17221
rect 25688 17212 25740 17264
rect 26056 17212 26108 17264
rect 20260 17144 20312 17153
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 25596 17187 25648 17196
rect 21088 17144 21140 17153
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 25964 17144 26016 17196
rect 27160 17144 27212 17196
rect 27988 17187 28040 17196
rect 27988 17153 27997 17187
rect 27997 17153 28031 17187
rect 28031 17153 28040 17187
rect 27988 17144 28040 17153
rect 38200 17187 38252 17196
rect 38200 17153 38209 17187
rect 38209 17153 38243 17187
rect 38243 17153 38252 17187
rect 38200 17144 38252 17153
rect 17868 17076 17920 17128
rect 18420 17119 18472 17128
rect 18420 17085 18429 17119
rect 18429 17085 18463 17119
rect 18463 17085 18472 17119
rect 18420 17076 18472 17085
rect 19340 17076 19392 17128
rect 15292 17008 15344 17060
rect 23572 17076 23624 17128
rect 24860 17076 24912 17128
rect 25504 17076 25556 17128
rect 20260 16940 20312 16992
rect 20628 16940 20680 16992
rect 21916 16940 21968 16992
rect 22008 16940 22060 16992
rect 25136 16940 25188 16992
rect 26424 17008 26476 17060
rect 38016 17051 38068 17060
rect 38016 17017 38025 17051
rect 38025 17017 38059 17051
rect 38059 17017 38068 17051
rect 38016 17008 38068 17017
rect 27068 16940 27120 16992
rect 27160 16940 27212 16992
rect 29276 16940 29328 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 12900 16600 12952 16652
rect 14648 16600 14700 16652
rect 20444 16668 20496 16720
rect 21088 16668 21140 16720
rect 22008 16668 22060 16720
rect 2872 16439 2924 16448
rect 2872 16405 2881 16439
rect 2881 16405 2915 16439
rect 2915 16405 2924 16439
rect 2872 16396 2924 16405
rect 17408 16532 17460 16584
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 21180 16643 21232 16652
rect 21180 16609 21189 16643
rect 21189 16609 21223 16643
rect 21223 16609 21232 16643
rect 21180 16600 21232 16609
rect 21364 16600 21416 16652
rect 22744 16736 22796 16788
rect 22652 16668 22704 16720
rect 24308 16736 24360 16788
rect 26056 16736 26108 16788
rect 26148 16736 26200 16788
rect 25596 16668 25648 16720
rect 26332 16668 26384 16720
rect 23664 16600 23716 16652
rect 24768 16643 24820 16652
rect 24768 16609 24777 16643
rect 24777 16609 24811 16643
rect 24811 16609 24820 16643
rect 24768 16600 24820 16609
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 19248 16532 19300 16584
rect 20076 16532 20128 16584
rect 28356 16643 28408 16652
rect 28356 16609 28365 16643
rect 28365 16609 28399 16643
rect 28399 16609 28408 16643
rect 28356 16600 28408 16609
rect 28816 16643 28868 16652
rect 28816 16609 28825 16643
rect 28825 16609 28859 16643
rect 28859 16609 28868 16643
rect 28816 16600 28868 16609
rect 19340 16464 19392 16516
rect 20628 16507 20680 16516
rect 20628 16473 20637 16507
rect 20637 16473 20671 16507
rect 20671 16473 20680 16507
rect 21732 16507 21784 16516
rect 20628 16464 20680 16473
rect 21732 16473 21741 16507
rect 21741 16473 21775 16507
rect 21775 16473 21784 16507
rect 21732 16464 21784 16473
rect 22376 16464 22428 16516
rect 23388 16507 23440 16516
rect 23388 16473 23397 16507
rect 23397 16473 23431 16507
rect 23431 16473 23440 16507
rect 23388 16464 23440 16473
rect 24952 16464 25004 16516
rect 25136 16507 25188 16516
rect 25136 16473 25145 16507
rect 25145 16473 25179 16507
rect 25179 16473 25188 16507
rect 25136 16464 25188 16473
rect 25688 16464 25740 16516
rect 26608 16464 26660 16516
rect 4620 16396 4672 16448
rect 15752 16396 15804 16448
rect 18052 16396 18104 16448
rect 21916 16396 21968 16448
rect 26792 16464 26844 16516
rect 27620 16464 27672 16516
rect 27160 16396 27212 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16124 2188 16176
rect 15752 16167 15804 16176
rect 15752 16133 15761 16167
rect 15761 16133 15795 16167
rect 15795 16133 15804 16167
rect 15752 16124 15804 16133
rect 17132 16124 17184 16176
rect 22468 16124 22520 16176
rect 25504 16192 25556 16244
rect 23848 16167 23900 16176
rect 23848 16133 23857 16167
rect 23857 16133 23891 16167
rect 23891 16133 23900 16167
rect 23848 16124 23900 16133
rect 26240 16124 26292 16176
rect 26424 16167 26476 16176
rect 26424 16133 26433 16167
rect 26433 16133 26467 16167
rect 26467 16133 26476 16167
rect 26424 16124 26476 16133
rect 26516 16167 26568 16176
rect 26516 16133 26525 16167
rect 26525 16133 26559 16167
rect 26559 16133 26568 16167
rect 26516 16124 26568 16133
rect 28724 16124 28776 16176
rect 10600 16056 10652 16108
rect 19248 16099 19300 16108
rect 10508 15988 10560 16040
rect 18420 15988 18472 16040
rect 16948 15920 17000 15972
rect 17684 15963 17736 15972
rect 17684 15929 17693 15963
rect 17693 15929 17727 15963
rect 17727 15929 17736 15963
rect 17684 15920 17736 15929
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 16396 15852 16448 15904
rect 17224 15852 17276 15904
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 20628 16056 20680 16108
rect 31392 16056 31444 16108
rect 38200 16099 38252 16108
rect 38200 16065 38209 16099
rect 38209 16065 38243 16099
rect 38243 16065 38252 16099
rect 38200 16056 38252 16065
rect 18604 15920 18656 15972
rect 20720 15963 20772 15972
rect 20720 15929 20729 15963
rect 20729 15929 20763 15963
rect 20763 15929 20772 15963
rect 20720 15920 20772 15929
rect 22192 15988 22244 16040
rect 23020 15988 23072 16040
rect 23664 15988 23716 16040
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 24952 15988 25004 16040
rect 25412 15988 25464 16040
rect 22652 15963 22704 15972
rect 22192 15852 22244 15904
rect 22652 15929 22661 15963
rect 22661 15929 22695 15963
rect 22695 15929 22704 15963
rect 22652 15920 22704 15929
rect 25504 15920 25556 15972
rect 25964 15963 26016 15972
rect 25964 15929 25973 15963
rect 25973 15929 26007 15963
rect 26007 15929 26016 15963
rect 25964 15920 26016 15929
rect 26240 15988 26292 16040
rect 27068 15988 27120 16040
rect 28080 16031 28132 16040
rect 28080 15997 28089 16031
rect 28089 15997 28123 16031
rect 28123 15997 28132 16031
rect 28080 15988 28132 15997
rect 29552 15920 29604 15972
rect 24768 15852 24820 15904
rect 26976 15852 27028 15904
rect 27620 15852 27672 15904
rect 29000 15852 29052 15904
rect 29460 15895 29512 15904
rect 29460 15861 29469 15895
rect 29469 15861 29503 15895
rect 29503 15861 29512 15895
rect 29460 15852 29512 15861
rect 38108 15895 38160 15904
rect 38108 15861 38117 15895
rect 38117 15861 38151 15895
rect 38151 15861 38160 15895
rect 38108 15852 38160 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 10508 15691 10560 15700
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 17132 15691 17184 15700
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 18052 15648 18104 15700
rect 21640 15648 21692 15700
rect 15384 15623 15436 15632
rect 15384 15589 15393 15623
rect 15393 15589 15427 15623
rect 15427 15589 15436 15623
rect 15384 15580 15436 15589
rect 17316 15580 17368 15632
rect 17684 15512 17736 15564
rect 4620 15444 4672 15496
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 19432 15512 19484 15564
rect 20444 15512 20496 15564
rect 20996 15555 21048 15564
rect 20996 15521 21005 15555
rect 21005 15521 21039 15555
rect 21039 15521 21048 15555
rect 20996 15512 21048 15521
rect 21456 15512 21508 15564
rect 22192 15580 22244 15632
rect 25688 15648 25740 15700
rect 25780 15648 25832 15700
rect 26056 15648 26108 15700
rect 36820 15648 36872 15700
rect 25228 15555 25280 15564
rect 25228 15521 25237 15555
rect 25237 15521 25271 15555
rect 25271 15521 25280 15555
rect 25596 15580 25648 15632
rect 25228 15512 25280 15521
rect 38108 15512 38160 15564
rect 21364 15444 21416 15496
rect 25780 15444 25832 15496
rect 26056 15444 26108 15496
rect 21732 15419 21784 15428
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 16672 15308 16724 15360
rect 18512 15308 18564 15360
rect 19156 15308 19208 15360
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 21732 15385 21741 15419
rect 21741 15385 21775 15419
rect 21775 15385 21784 15419
rect 21732 15376 21784 15385
rect 21916 15376 21968 15428
rect 22284 15308 22336 15360
rect 22836 15376 22888 15428
rect 23480 15419 23532 15428
rect 23480 15385 23489 15419
rect 23489 15385 23523 15419
rect 23523 15385 23532 15419
rect 23480 15376 23532 15385
rect 24492 15376 24544 15428
rect 26976 15419 27028 15428
rect 23572 15308 23624 15360
rect 25688 15308 25740 15360
rect 26700 15308 26752 15360
rect 26976 15385 26985 15419
rect 26985 15385 27019 15419
rect 27019 15385 27028 15419
rect 26976 15376 27028 15385
rect 28080 15376 28132 15428
rect 29736 15444 29788 15496
rect 30196 15376 30248 15428
rect 30380 15351 30432 15360
rect 30380 15317 30389 15351
rect 30389 15317 30423 15351
rect 30423 15317 30432 15351
rect 30380 15308 30432 15317
rect 31300 15308 31352 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 13636 15036 13688 15088
rect 14648 15011 14700 15020
rect 13912 14764 13964 14816
rect 14648 14977 14657 15011
rect 14657 14977 14691 15011
rect 14691 14977 14700 15011
rect 14648 14968 14700 14977
rect 15752 14832 15804 14884
rect 16580 14968 16632 15020
rect 16672 14968 16724 15020
rect 18512 15036 18564 15088
rect 19524 15079 19576 15088
rect 19524 15045 19533 15079
rect 19533 15045 19567 15079
rect 19567 15045 19576 15079
rect 19524 15036 19576 15045
rect 20352 15104 20404 15156
rect 22100 15147 22152 15156
rect 22100 15113 22109 15147
rect 22109 15113 22143 15147
rect 22143 15113 22152 15147
rect 22100 15104 22152 15113
rect 25228 15104 25280 15156
rect 24400 15079 24452 15088
rect 24400 15045 24409 15079
rect 24409 15045 24443 15079
rect 24443 15045 24452 15079
rect 24400 15036 24452 15045
rect 25136 15036 25188 15088
rect 28448 15104 28500 15156
rect 27068 15036 27120 15088
rect 28540 15036 28592 15088
rect 25044 15011 25096 15020
rect 16488 14900 16540 14952
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 18328 14900 18380 14952
rect 19248 14900 19300 14952
rect 19432 14943 19484 14952
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 16672 14764 16724 14816
rect 23664 14900 23716 14952
rect 25044 14977 25053 15011
rect 25053 14977 25087 15011
rect 25087 14977 25096 15011
rect 25044 14968 25096 14977
rect 29460 15104 29512 15156
rect 29920 15104 29972 15156
rect 25136 14900 25188 14952
rect 19984 14875 20036 14884
rect 19984 14841 19993 14875
rect 19993 14841 20027 14875
rect 20027 14841 20036 14875
rect 19984 14832 20036 14841
rect 24032 14832 24084 14884
rect 19340 14764 19392 14816
rect 20628 14807 20680 14816
rect 20628 14773 20637 14807
rect 20637 14773 20671 14807
rect 20671 14773 20680 14807
rect 20628 14764 20680 14773
rect 21272 14764 21324 14816
rect 29000 14968 29052 15020
rect 29368 14968 29420 15020
rect 30104 14968 30156 15020
rect 25596 14900 25648 14952
rect 26516 14943 26568 14952
rect 26516 14909 26525 14943
rect 26525 14909 26559 14943
rect 26559 14909 26568 14943
rect 26516 14900 26568 14909
rect 27344 14900 27396 14952
rect 28080 14943 28132 14952
rect 28080 14909 28089 14943
rect 28089 14909 28123 14943
rect 28123 14909 28132 14943
rect 28080 14900 28132 14909
rect 28356 14900 28408 14952
rect 30380 14900 30432 14952
rect 26332 14832 26384 14884
rect 27068 14832 27120 14884
rect 27804 14832 27856 14884
rect 27896 14832 27948 14884
rect 29552 14832 29604 14884
rect 27712 14764 27764 14816
rect 30288 14764 30340 14816
rect 31300 15104 31352 15156
rect 33968 15104 34020 15156
rect 38108 14764 38160 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 14188 14560 14240 14612
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 15384 14492 15436 14544
rect 14832 14356 14884 14408
rect 15844 14356 15896 14408
rect 18696 14560 18748 14612
rect 19524 14603 19576 14612
rect 19524 14569 19533 14603
rect 19533 14569 19567 14603
rect 19567 14569 19576 14603
rect 19524 14560 19576 14569
rect 19984 14560 20036 14612
rect 23848 14560 23900 14612
rect 24400 14560 24452 14612
rect 27344 14560 27396 14612
rect 20076 14492 20128 14544
rect 18144 14424 18196 14476
rect 19432 14424 19484 14476
rect 20352 14492 20404 14544
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17408 14356 17460 14408
rect 19616 14399 19668 14408
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 15384 14263 15436 14272
rect 15384 14229 15393 14263
rect 15393 14229 15427 14263
rect 15427 14229 15436 14263
rect 15384 14220 15436 14229
rect 18328 14288 18380 14340
rect 19156 14288 19208 14340
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20260 14424 20312 14476
rect 20260 14331 20312 14340
rect 20260 14297 20269 14331
rect 20269 14297 20303 14331
rect 20303 14297 20312 14331
rect 20260 14288 20312 14297
rect 20904 14331 20956 14340
rect 17960 14220 18012 14272
rect 20904 14297 20913 14331
rect 20913 14297 20947 14331
rect 20947 14297 20956 14331
rect 20904 14288 20956 14297
rect 20444 14220 20496 14272
rect 21272 14220 21324 14272
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 21824 14356 21876 14408
rect 25044 14492 25096 14544
rect 25320 14492 25372 14544
rect 26056 14492 26108 14544
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 25780 14424 25832 14476
rect 26148 14467 26200 14476
rect 26148 14433 26157 14467
rect 26157 14433 26191 14467
rect 26191 14433 26200 14467
rect 26148 14424 26200 14433
rect 26240 14424 26292 14476
rect 27160 14424 27212 14476
rect 25688 14356 25740 14408
rect 26700 14356 26752 14408
rect 22008 14220 22060 14272
rect 23296 14331 23348 14340
rect 23296 14297 23305 14331
rect 23305 14297 23339 14331
rect 23339 14297 23348 14331
rect 23296 14288 23348 14297
rect 23848 14288 23900 14340
rect 26148 14288 26200 14340
rect 26240 14288 26292 14340
rect 27344 14288 27396 14340
rect 29092 14492 29144 14544
rect 30012 14492 30064 14544
rect 28080 14424 28132 14476
rect 27804 14356 27856 14408
rect 28448 14399 28500 14408
rect 28448 14365 28457 14399
rect 28457 14365 28491 14399
rect 28491 14365 28500 14399
rect 28448 14356 28500 14365
rect 29920 14399 29972 14408
rect 29920 14365 29929 14399
rect 29929 14365 29963 14399
rect 29963 14365 29972 14399
rect 29920 14356 29972 14365
rect 30288 14288 30340 14340
rect 23388 14220 23440 14272
rect 24676 14263 24728 14272
rect 24676 14229 24685 14263
rect 24685 14229 24719 14263
rect 24719 14229 24728 14263
rect 24676 14220 24728 14229
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 25320 14220 25372 14272
rect 26056 14220 26108 14272
rect 27804 14220 27856 14272
rect 29736 14220 29788 14272
rect 30380 14220 30432 14272
rect 31208 14220 31260 14272
rect 36820 14220 36872 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 17408 14016 17460 14068
rect 22100 14016 22152 14068
rect 22192 14016 22244 14068
rect 13360 13948 13412 14000
rect 13636 13991 13688 14000
rect 13636 13957 13645 13991
rect 13645 13957 13679 13991
rect 13679 13957 13688 13991
rect 13636 13948 13688 13957
rect 14280 13991 14332 14000
rect 14280 13957 14289 13991
rect 14289 13957 14323 13991
rect 14323 13957 14332 13991
rect 14280 13948 14332 13957
rect 18144 13991 18196 14000
rect 18144 13957 18153 13991
rect 18153 13957 18187 13991
rect 18187 13957 18196 13991
rect 18144 13948 18196 13957
rect 19064 13991 19116 14000
rect 19064 13957 19073 13991
rect 19073 13957 19107 13991
rect 19107 13957 19116 13991
rect 19064 13948 19116 13957
rect 19156 13991 19208 14000
rect 19156 13957 19165 13991
rect 19165 13957 19199 13991
rect 19199 13957 19208 13991
rect 19156 13948 19208 13957
rect 20352 13948 20404 14000
rect 23388 13948 23440 14000
rect 24676 13948 24728 14000
rect 24768 13948 24820 14000
rect 26332 13991 26384 14000
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 15476 13923 15528 13932
rect 4068 13812 4120 13864
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 16580 13880 16632 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 19340 13880 19392 13932
rect 20444 13880 20496 13932
rect 21364 13880 21416 13932
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 25044 13880 25096 13932
rect 16304 13812 16356 13864
rect 16764 13812 16816 13864
rect 18144 13812 18196 13864
rect 18328 13812 18380 13864
rect 23848 13812 23900 13864
rect 25320 13812 25372 13864
rect 26332 13957 26341 13991
rect 26341 13957 26375 13991
rect 26375 13957 26384 13991
rect 26332 13948 26384 13957
rect 26424 13948 26476 14000
rect 27068 13948 27120 14000
rect 27252 14016 27304 14068
rect 27712 13991 27764 14000
rect 27712 13957 27721 13991
rect 27721 13957 27755 13991
rect 27755 13957 27764 13991
rect 27712 13948 27764 13957
rect 27804 13991 27856 14000
rect 27804 13957 27813 13991
rect 27813 13957 27847 13991
rect 27847 13957 27856 13991
rect 27804 13948 27856 13957
rect 13176 13787 13228 13796
rect 13176 13753 13185 13787
rect 13185 13753 13219 13787
rect 13219 13753 13228 13787
rect 13176 13744 13228 13753
rect 14740 13744 14792 13796
rect 18052 13744 18104 13796
rect 14188 13676 14240 13728
rect 21088 13744 21140 13796
rect 21180 13787 21232 13796
rect 21180 13753 21189 13787
rect 21189 13753 21223 13787
rect 21223 13753 21232 13787
rect 21180 13744 21232 13753
rect 23388 13744 23440 13796
rect 23664 13744 23716 13796
rect 23940 13744 23992 13796
rect 24584 13744 24636 13796
rect 27804 13812 27856 13864
rect 28080 13812 28132 13864
rect 28908 13855 28960 13864
rect 28908 13821 28917 13855
rect 28917 13821 28951 13855
rect 28951 13821 28960 13855
rect 28908 13812 28960 13821
rect 20536 13676 20588 13728
rect 24768 13676 24820 13728
rect 27160 13744 27212 13796
rect 28264 13744 28316 13796
rect 29184 13744 29236 13796
rect 29736 13923 29788 13932
rect 29736 13889 29745 13923
rect 29745 13889 29779 13923
rect 29779 13889 29788 13923
rect 29736 13880 29788 13889
rect 30196 14016 30248 14068
rect 30472 14016 30524 14068
rect 29920 13948 29972 14000
rect 29644 13855 29696 13864
rect 29644 13821 29653 13855
rect 29653 13821 29687 13855
rect 29687 13821 29696 13855
rect 29644 13812 29696 13821
rect 29828 13812 29880 13864
rect 31576 13812 31628 13864
rect 33140 13812 33192 13864
rect 38292 13855 38344 13864
rect 38292 13821 38301 13855
rect 38301 13821 38335 13855
rect 38335 13821 38344 13855
rect 38292 13812 38344 13821
rect 29736 13676 29788 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10600 13515 10652 13524
rect 10600 13481 10609 13515
rect 10609 13481 10643 13515
rect 10643 13481 10652 13515
rect 10600 13472 10652 13481
rect 14740 13404 14792 13456
rect 15476 13472 15528 13524
rect 16856 13472 16908 13524
rect 17960 13472 18012 13524
rect 19248 13472 19300 13524
rect 17224 13404 17276 13456
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 16120 13336 16172 13388
rect 15292 13268 15344 13320
rect 14372 13200 14424 13252
rect 13360 13132 13412 13184
rect 15752 13243 15804 13252
rect 15752 13209 15761 13243
rect 15761 13209 15795 13243
rect 15795 13209 15804 13243
rect 17132 13268 17184 13320
rect 18052 13336 18104 13388
rect 20168 13404 20220 13456
rect 20352 13472 20404 13524
rect 20444 13404 20496 13456
rect 20904 13404 20956 13456
rect 21640 13404 21692 13456
rect 22008 13472 22060 13524
rect 22560 13472 22612 13524
rect 28448 13472 28500 13524
rect 28632 13472 28684 13524
rect 31116 13515 31168 13524
rect 23388 13404 23440 13456
rect 19432 13336 19484 13388
rect 20536 13336 20588 13388
rect 15752 13200 15804 13209
rect 15384 13132 15436 13184
rect 18052 13200 18104 13252
rect 18972 13200 19024 13252
rect 20720 13200 20772 13252
rect 21272 13336 21324 13388
rect 22100 13200 22152 13252
rect 22284 13243 22336 13252
rect 22284 13209 22293 13243
rect 22293 13209 22327 13243
rect 22327 13209 22336 13243
rect 22744 13336 22796 13388
rect 23112 13336 23164 13388
rect 25596 13336 25648 13388
rect 25688 13336 25740 13388
rect 25964 13379 26016 13388
rect 25964 13345 25973 13379
rect 25973 13345 26007 13379
rect 26007 13345 26016 13379
rect 25964 13336 26016 13345
rect 26516 13336 26568 13388
rect 27528 13404 27580 13456
rect 29092 13404 29144 13456
rect 27436 13336 27488 13388
rect 31116 13481 31125 13515
rect 31125 13481 31159 13515
rect 31159 13481 31168 13515
rect 31116 13472 31168 13481
rect 38292 13515 38344 13524
rect 38292 13481 38301 13515
rect 38301 13481 38335 13515
rect 38335 13481 38344 13515
rect 38292 13472 38344 13481
rect 28264 13268 28316 13320
rect 29184 13311 29236 13320
rect 29184 13277 29193 13311
rect 29193 13277 29227 13311
rect 29227 13277 29236 13311
rect 31208 13336 31260 13388
rect 37096 13336 37148 13388
rect 29184 13268 29236 13277
rect 22836 13243 22888 13252
rect 22284 13200 22336 13209
rect 18512 13132 18564 13184
rect 22560 13132 22612 13184
rect 22836 13209 22845 13243
rect 22845 13209 22879 13243
rect 22879 13209 22888 13243
rect 22836 13200 22888 13209
rect 24768 13243 24820 13252
rect 24768 13209 24777 13243
rect 24777 13209 24811 13243
rect 24811 13209 24820 13243
rect 24768 13200 24820 13209
rect 24952 13200 25004 13252
rect 25964 13200 26016 13252
rect 26424 13132 26476 13184
rect 27620 13200 27672 13252
rect 27712 13200 27764 13252
rect 28908 13200 28960 13252
rect 30748 13268 30800 13320
rect 27896 13132 27948 13184
rect 28172 13132 28224 13184
rect 30196 13132 30248 13184
rect 30472 13175 30524 13184
rect 30472 13141 30481 13175
rect 30481 13141 30515 13175
rect 30515 13141 30524 13175
rect 30472 13132 30524 13141
rect 37924 13132 37976 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 13084 12928 13136 12980
rect 10968 12792 11020 12844
rect 13360 12792 13412 12844
rect 14188 12835 14240 12844
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 17960 12860 18012 12912
rect 22560 12928 22612 12980
rect 18972 12860 19024 12912
rect 19524 12860 19576 12912
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 15568 12792 15620 12844
rect 16396 12792 16448 12844
rect 17408 12792 17460 12844
rect 14372 12724 14424 12776
rect 14188 12656 14240 12708
rect 15476 12656 15528 12708
rect 16764 12724 16816 12776
rect 20076 12835 20128 12844
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 20260 12724 20312 12776
rect 17132 12656 17184 12708
rect 20812 12724 20864 12776
rect 22284 12860 22336 12912
rect 26424 12928 26476 12980
rect 27528 12928 27580 12980
rect 25596 12903 25648 12912
rect 25596 12869 25605 12903
rect 25605 12869 25639 12903
rect 25639 12869 25648 12903
rect 25596 12860 25648 12869
rect 29000 12928 29052 12980
rect 29092 12928 29144 12980
rect 30380 12928 30432 12980
rect 30932 12971 30984 12980
rect 30932 12937 30941 12971
rect 30941 12937 30975 12971
rect 30975 12937 30984 12971
rect 30932 12928 30984 12937
rect 21180 12792 21232 12844
rect 21456 12792 21508 12844
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 13636 12631 13688 12640
rect 13636 12597 13645 12631
rect 13645 12597 13679 12631
rect 13679 12597 13688 12631
rect 13636 12588 13688 12597
rect 15292 12588 15344 12640
rect 15936 12588 15988 12640
rect 16488 12588 16540 12640
rect 21180 12656 21232 12708
rect 22192 12724 22244 12776
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 24124 12724 24176 12776
rect 24492 12767 24544 12776
rect 24492 12733 24501 12767
rect 24501 12733 24535 12767
rect 24535 12733 24544 12767
rect 24492 12724 24544 12733
rect 26516 12724 26568 12776
rect 28448 12903 28500 12912
rect 28448 12869 28457 12903
rect 28457 12869 28491 12903
rect 28491 12869 28500 12903
rect 28448 12860 28500 12869
rect 29828 12860 29880 12912
rect 29736 12835 29788 12844
rect 29736 12801 29745 12835
rect 29745 12801 29779 12835
rect 29779 12801 29788 12835
rect 29736 12792 29788 12801
rect 31300 12860 31352 12912
rect 38016 12928 38068 12980
rect 31208 12792 31260 12844
rect 21088 12588 21140 12640
rect 27620 12656 27672 12708
rect 27804 12767 27856 12776
rect 27804 12733 27813 12767
rect 27813 12733 27847 12767
rect 27847 12733 27856 12767
rect 27804 12724 27856 12733
rect 28172 12724 28224 12776
rect 28816 12767 28868 12776
rect 28816 12733 28825 12767
rect 28825 12733 28859 12767
rect 28859 12733 28868 12767
rect 28816 12724 28868 12733
rect 29460 12724 29512 12776
rect 33232 12835 33284 12844
rect 33232 12801 33241 12835
rect 33241 12801 33275 12835
rect 33275 12801 33284 12835
rect 33232 12792 33284 12801
rect 23480 12588 23532 12640
rect 24676 12588 24728 12640
rect 27528 12588 27580 12640
rect 30196 12588 30248 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 16488 12384 16540 12436
rect 16856 12316 16908 12368
rect 17408 12384 17460 12436
rect 18328 12384 18380 12436
rect 18604 12384 18656 12436
rect 21088 12384 21140 12436
rect 21548 12384 21600 12436
rect 21732 12384 21784 12436
rect 18972 12316 19024 12368
rect 22744 12316 22796 12368
rect 25964 12316 26016 12368
rect 15016 12248 15068 12300
rect 18236 12291 18288 12300
rect 18236 12257 18245 12291
rect 18245 12257 18279 12291
rect 18279 12257 18288 12291
rect 18236 12248 18288 12257
rect 14096 12180 14148 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 13728 12112 13780 12164
rect 15384 12155 15436 12164
rect 15384 12121 15393 12155
rect 15393 12121 15427 12155
rect 15427 12121 15436 12155
rect 15384 12112 15436 12121
rect 15476 12155 15528 12164
rect 15476 12121 15485 12155
rect 15485 12121 15519 12155
rect 15519 12121 15528 12155
rect 15476 12112 15528 12121
rect 16304 12112 16356 12164
rect 16672 12155 16724 12164
rect 16672 12121 16681 12155
rect 16681 12121 16715 12155
rect 16715 12121 16724 12155
rect 16672 12112 16724 12121
rect 17316 12112 17368 12164
rect 18972 12112 19024 12164
rect 20168 12044 20220 12096
rect 21548 12248 21600 12300
rect 22008 12248 22060 12300
rect 23296 12248 23348 12300
rect 25412 12248 25464 12300
rect 26424 12291 26476 12300
rect 26424 12257 26433 12291
rect 26433 12257 26467 12291
rect 26467 12257 26476 12291
rect 26424 12248 26476 12257
rect 23572 12180 23624 12232
rect 21180 12155 21232 12164
rect 21180 12121 21189 12155
rect 21189 12121 21223 12155
rect 21223 12121 21232 12155
rect 21180 12112 21232 12121
rect 21548 12112 21600 12164
rect 21364 12044 21416 12096
rect 23848 12112 23900 12164
rect 22836 12044 22888 12096
rect 25780 12155 25832 12164
rect 25780 12121 25789 12155
rect 25789 12121 25823 12155
rect 25823 12121 25832 12155
rect 25780 12112 25832 12121
rect 29644 12384 29696 12436
rect 27068 12359 27120 12368
rect 27068 12325 27077 12359
rect 27077 12325 27111 12359
rect 27111 12325 27120 12359
rect 27068 12316 27120 12325
rect 28816 12359 28868 12368
rect 28816 12325 28825 12359
rect 28825 12325 28859 12359
rect 28859 12325 28868 12359
rect 28816 12316 28868 12325
rect 27344 12248 27396 12300
rect 28724 12248 28776 12300
rect 29736 12180 29788 12232
rect 27528 12155 27580 12164
rect 27528 12121 27537 12155
rect 27537 12121 27571 12155
rect 27571 12121 27580 12155
rect 27528 12112 27580 12121
rect 27620 12112 27672 12164
rect 29644 12112 29696 12164
rect 30196 12180 30248 12232
rect 31024 12223 31076 12232
rect 31024 12189 31033 12223
rect 31033 12189 31067 12223
rect 31067 12189 31076 12223
rect 31024 12180 31076 12189
rect 31116 12223 31168 12232
rect 31116 12189 31125 12223
rect 31125 12189 31159 12223
rect 31159 12189 31168 12223
rect 31116 12180 31168 12189
rect 30564 12112 30616 12164
rect 27436 12044 27488 12096
rect 27712 12044 27764 12096
rect 31208 12044 31260 12096
rect 31484 12044 31536 12096
rect 31668 12087 31720 12096
rect 31668 12053 31677 12087
rect 31677 12053 31711 12087
rect 31711 12053 31720 12087
rect 31668 12044 31720 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 13728 11883 13780 11892
rect 13728 11849 13737 11883
rect 13737 11849 13771 11883
rect 13771 11849 13780 11883
rect 13728 11840 13780 11849
rect 11980 11815 12032 11824
rect 11980 11781 11989 11815
rect 11989 11781 12023 11815
rect 12023 11781 12032 11815
rect 11980 11772 12032 11781
rect 16304 11815 16356 11824
rect 16304 11781 16313 11815
rect 16313 11781 16347 11815
rect 16347 11781 16356 11815
rect 16304 11772 16356 11781
rect 13452 11704 13504 11756
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 14648 11636 14700 11688
rect 17408 11772 17460 11824
rect 17776 11815 17828 11824
rect 17776 11781 17785 11815
rect 17785 11781 17819 11815
rect 17819 11781 17828 11815
rect 17776 11772 17828 11781
rect 20260 11840 20312 11892
rect 21548 11840 21600 11892
rect 23848 11840 23900 11892
rect 26056 11840 26108 11892
rect 26332 11840 26384 11892
rect 19156 11772 19208 11824
rect 20352 11772 20404 11824
rect 22100 11772 22152 11824
rect 22744 11772 22796 11824
rect 23388 11772 23440 11824
rect 24584 11772 24636 11824
rect 27160 11815 27212 11824
rect 27160 11781 27169 11815
rect 27169 11781 27203 11815
rect 27203 11781 27212 11815
rect 27160 11772 27212 11781
rect 31116 11840 31168 11892
rect 31576 11883 31628 11892
rect 31576 11849 31585 11883
rect 31585 11849 31619 11883
rect 31619 11849 31628 11883
rect 31576 11840 31628 11849
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 27068 11704 27120 11756
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 17408 11636 17460 11688
rect 16580 11568 16632 11620
rect 17960 11636 18012 11688
rect 18972 11636 19024 11688
rect 19432 11679 19484 11688
rect 19432 11645 19441 11679
rect 19441 11645 19475 11679
rect 19475 11645 19484 11679
rect 19432 11636 19484 11645
rect 21180 11636 21232 11688
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 23848 11636 23900 11688
rect 25044 11636 25096 11688
rect 27804 11679 27856 11688
rect 18604 11568 18656 11620
rect 15108 11500 15160 11552
rect 20720 11568 20772 11620
rect 27804 11645 27813 11679
rect 27813 11645 27847 11679
rect 27847 11645 27856 11679
rect 27804 11636 27856 11645
rect 18880 11500 18932 11552
rect 21364 11500 21416 11552
rect 21548 11500 21600 11552
rect 27252 11568 27304 11620
rect 29184 11772 29236 11824
rect 29460 11772 29512 11824
rect 29736 11704 29788 11756
rect 32312 11772 32364 11824
rect 30932 11747 30984 11756
rect 30932 11713 30941 11747
rect 30941 11713 30975 11747
rect 30975 11713 30984 11747
rect 30932 11704 30984 11713
rect 31208 11704 31260 11756
rect 38200 11747 38252 11756
rect 28448 11636 28500 11688
rect 30196 11636 30248 11688
rect 31116 11636 31168 11688
rect 38200 11713 38209 11747
rect 38209 11713 38243 11747
rect 38243 11713 38252 11747
rect 38200 11704 38252 11713
rect 23020 11500 23072 11552
rect 28264 11500 28316 11552
rect 29092 11500 29144 11552
rect 32312 11543 32364 11552
rect 32312 11509 32321 11543
rect 32321 11509 32355 11543
rect 32355 11509 32364 11543
rect 32312 11500 32364 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 8944 11296 8996 11348
rect 17776 11296 17828 11348
rect 18052 11296 18104 11348
rect 19340 11296 19392 11348
rect 23572 11296 23624 11348
rect 27712 11339 27764 11348
rect 27712 11305 27721 11339
rect 27721 11305 27755 11339
rect 27755 11305 27764 11339
rect 27712 11296 27764 11305
rect 27804 11296 27856 11348
rect 14188 11228 14240 11280
rect 17316 11271 17368 11280
rect 15384 11160 15436 11212
rect 17316 11237 17325 11271
rect 17325 11237 17359 11271
rect 17359 11237 17368 11271
rect 17316 11228 17368 11237
rect 18972 11228 19024 11280
rect 16764 11203 16816 11212
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14464 11092 14516 11144
rect 15476 11092 15528 11144
rect 16764 11169 16773 11203
rect 16773 11169 16807 11203
rect 16807 11169 16816 11203
rect 16764 11160 16816 11169
rect 17684 11160 17736 11212
rect 18604 11160 18656 11212
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 15384 11024 15436 11076
rect 18328 11092 18380 11144
rect 16396 11024 16448 11076
rect 16212 10999 16264 11008
rect 16212 10965 16221 10999
rect 16221 10965 16255 10999
rect 16255 10965 16264 10999
rect 16212 10956 16264 10965
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 19432 11160 19484 11212
rect 20352 11228 20404 11280
rect 20444 11228 20496 11280
rect 22008 11228 22060 11280
rect 22560 11228 22612 11280
rect 19524 11092 19576 11144
rect 20812 11135 20864 11144
rect 20812 11101 20821 11135
rect 20821 11101 20855 11135
rect 20855 11101 20864 11135
rect 20812 11092 20864 11101
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 26240 11160 26292 11212
rect 26332 11160 26384 11212
rect 29000 11296 29052 11348
rect 29184 11228 29236 11280
rect 30472 11228 30524 11280
rect 33508 11228 33560 11280
rect 32404 11160 32456 11212
rect 23848 11092 23900 11101
rect 29736 11092 29788 11144
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30380 11135 30432 11144
rect 30380 11101 30389 11135
rect 30389 11101 30423 11135
rect 30423 11101 30432 11135
rect 30380 11092 30432 11101
rect 33416 11135 33468 11144
rect 33416 11101 33425 11135
rect 33425 11101 33459 11135
rect 33459 11101 33468 11135
rect 33416 11092 33468 11101
rect 16856 11024 16908 11033
rect 17132 10956 17184 11008
rect 18604 10956 18656 11008
rect 20996 11024 21048 11076
rect 22192 11024 22244 11076
rect 23296 11024 23348 11076
rect 25136 11067 25188 11076
rect 22100 10956 22152 11008
rect 22836 10956 22888 11008
rect 25136 11033 25145 11067
rect 25145 11033 25179 11067
rect 25179 11033 25188 11067
rect 25136 11024 25188 11033
rect 25228 11067 25280 11076
rect 25228 11033 25237 11067
rect 25237 11033 25271 11067
rect 25271 11033 25280 11067
rect 25228 11024 25280 11033
rect 27528 11024 27580 11076
rect 29184 11024 29236 11076
rect 30012 11024 30064 11076
rect 31668 11024 31720 11076
rect 26056 10956 26108 11008
rect 30288 10956 30340 11008
rect 30472 10999 30524 11008
rect 30472 10965 30481 10999
rect 30481 10965 30515 10999
rect 30515 10965 30524 10999
rect 30472 10956 30524 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 12900 10752 12952 10804
rect 13268 10752 13320 10804
rect 16580 10752 16632 10804
rect 22100 10752 22152 10804
rect 14280 10684 14332 10736
rect 15384 10684 15436 10736
rect 20812 10684 20864 10736
rect 21272 10727 21324 10736
rect 21272 10693 21281 10727
rect 21281 10693 21315 10727
rect 21315 10693 21324 10727
rect 21272 10684 21324 10693
rect 21456 10684 21508 10736
rect 21640 10684 21692 10736
rect 23480 10752 23532 10804
rect 23848 10752 23900 10804
rect 24032 10752 24084 10804
rect 23572 10727 23624 10736
rect 23572 10693 23581 10727
rect 23581 10693 23615 10727
rect 23615 10693 23624 10727
rect 23572 10684 23624 10693
rect 1584 10616 1636 10668
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 13636 10616 13688 10668
rect 15108 10616 15160 10668
rect 16580 10616 16632 10668
rect 17776 10616 17828 10668
rect 21364 10616 21416 10668
rect 25044 10727 25096 10736
rect 25044 10693 25053 10727
rect 25053 10693 25087 10727
rect 25087 10693 25096 10727
rect 25044 10684 25096 10693
rect 25504 10684 25556 10736
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 16028 10548 16080 10600
rect 18144 10548 18196 10600
rect 16672 10480 16724 10532
rect 17868 10480 17920 10532
rect 18328 10548 18380 10600
rect 19432 10548 19484 10600
rect 20260 10591 20312 10600
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 16212 10412 16264 10464
rect 19616 10412 19668 10464
rect 20260 10557 20269 10591
rect 20269 10557 20303 10591
rect 20303 10557 20312 10591
rect 20260 10548 20312 10557
rect 20444 10548 20496 10600
rect 22100 10548 22152 10600
rect 20904 10480 20956 10532
rect 27620 10752 27672 10804
rect 28448 10752 28500 10804
rect 28724 10752 28776 10804
rect 30932 10752 30984 10804
rect 31668 10795 31720 10804
rect 31668 10761 31677 10795
rect 31677 10761 31711 10795
rect 31711 10761 31720 10795
rect 31668 10752 31720 10761
rect 33416 10752 33468 10804
rect 27436 10684 27488 10736
rect 23204 10548 23256 10600
rect 22468 10412 22520 10464
rect 22836 10412 22888 10464
rect 24216 10548 24268 10600
rect 27252 10548 27304 10600
rect 28540 10548 28592 10600
rect 29368 10548 29420 10600
rect 30012 10591 30064 10600
rect 30012 10557 30021 10591
rect 30021 10557 30055 10591
rect 30055 10557 30064 10591
rect 30012 10548 30064 10557
rect 33140 10684 33192 10736
rect 38292 10659 38344 10668
rect 38292 10625 38301 10659
rect 38301 10625 38335 10659
rect 38335 10625 38344 10659
rect 38292 10616 38344 10625
rect 30196 10412 30248 10464
rect 30932 10412 30984 10464
rect 32036 10412 32088 10464
rect 33140 10412 33192 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 1768 10208 1820 10260
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 12532 10208 12584 10260
rect 15568 10208 15620 10260
rect 13360 10140 13412 10192
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 14556 10004 14608 10056
rect 14740 10004 14792 10056
rect 14832 10004 14884 10056
rect 15476 10004 15528 10056
rect 20628 10208 20680 10260
rect 20812 10251 20864 10260
rect 20812 10217 20821 10251
rect 20821 10217 20855 10251
rect 20855 10217 20864 10251
rect 20812 10208 20864 10217
rect 23664 10208 23716 10260
rect 17224 10183 17276 10192
rect 17224 10149 17233 10183
rect 17233 10149 17267 10183
rect 17267 10149 17276 10183
rect 17224 10140 17276 10149
rect 17776 10140 17828 10192
rect 19616 10140 19668 10192
rect 20444 10140 20496 10192
rect 18512 10115 18564 10124
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 25504 10140 25556 10192
rect 16672 9979 16724 9988
rect 16672 9945 16681 9979
rect 16681 9945 16715 9979
rect 16715 9945 16724 9979
rect 16672 9936 16724 9945
rect 16764 9979 16816 9988
rect 16764 9945 16773 9979
rect 16773 9945 16807 9979
rect 16807 9945 16816 9979
rect 17868 9979 17920 9988
rect 16764 9936 16816 9945
rect 17868 9945 17877 9979
rect 17877 9945 17911 9979
rect 17911 9945 17920 9979
rect 17868 9936 17920 9945
rect 17960 9979 18012 9988
rect 17960 9945 17969 9979
rect 17969 9945 18003 9979
rect 18003 9945 18012 9979
rect 17960 9936 18012 9945
rect 18144 9936 18196 9988
rect 23848 10072 23900 10124
rect 24492 10072 24544 10124
rect 26792 10208 26844 10260
rect 27620 10208 27672 10260
rect 27988 10208 28040 10260
rect 28724 10208 28776 10260
rect 28908 10251 28960 10260
rect 28908 10217 28917 10251
rect 28917 10217 28951 10251
rect 28951 10217 28960 10251
rect 28908 10208 28960 10217
rect 30288 10208 30340 10260
rect 32036 10251 32088 10260
rect 27252 10140 27304 10192
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 22008 10004 22060 10056
rect 23572 10004 23624 10056
rect 26240 10072 26292 10124
rect 27160 10115 27212 10124
rect 27160 10081 27169 10115
rect 27169 10081 27203 10115
rect 27203 10081 27212 10115
rect 27160 10072 27212 10081
rect 28080 10072 28132 10124
rect 30196 10140 30248 10192
rect 32036 10217 32045 10251
rect 32045 10217 32079 10251
rect 32079 10217 32088 10251
rect 32036 10208 32088 10217
rect 32312 10140 32364 10192
rect 30012 10072 30064 10124
rect 29644 10004 29696 10056
rect 19340 9936 19392 9988
rect 19616 9936 19668 9988
rect 19984 9979 20036 9988
rect 19984 9945 19993 9979
rect 19993 9945 20027 9979
rect 20027 9945 20036 9979
rect 19984 9936 20036 9945
rect 20536 9936 20588 9988
rect 20720 9936 20772 9988
rect 21272 9936 21324 9988
rect 23756 9936 23808 9988
rect 24860 9936 24912 9988
rect 26792 9936 26844 9988
rect 27988 9936 28040 9988
rect 33140 10072 33192 10124
rect 15752 9868 15804 9920
rect 18328 9868 18380 9920
rect 18604 9868 18656 9920
rect 24032 9868 24084 9920
rect 24124 9868 24176 9920
rect 24768 9868 24820 9920
rect 28080 9868 28132 9920
rect 28448 9868 28500 9920
rect 29552 9868 29604 9920
rect 29736 9868 29788 9920
rect 30472 9868 30524 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 6828 9664 6880 9716
rect 9220 9664 9272 9716
rect 11980 9596 12032 9648
rect 14740 9664 14792 9716
rect 20812 9664 20864 9716
rect 20904 9664 20956 9716
rect 22468 9664 22520 9716
rect 15844 9596 15896 9648
rect 17684 9639 17736 9648
rect 17684 9605 17693 9639
rect 17693 9605 17727 9639
rect 17727 9605 17736 9639
rect 17684 9596 17736 9605
rect 18328 9639 18380 9648
rect 18328 9605 18337 9639
rect 18337 9605 18371 9639
rect 18371 9605 18380 9639
rect 18328 9596 18380 9605
rect 18880 9596 18932 9648
rect 22284 9596 22336 9648
rect 22376 9596 22428 9648
rect 24768 9664 24820 9716
rect 25688 9664 25740 9716
rect 34796 9664 34848 9716
rect 24124 9596 24176 9648
rect 25596 9596 25648 9648
rect 25964 9596 26016 9648
rect 27528 9596 27580 9648
rect 27620 9596 27672 9648
rect 29644 9639 29696 9648
rect 29644 9605 29653 9639
rect 29653 9605 29687 9639
rect 29687 9605 29696 9639
rect 29644 9596 29696 9605
rect 30012 9596 30064 9648
rect 30564 9596 30616 9648
rect 30656 9596 30708 9648
rect 32772 9596 32824 9648
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 13912 9528 13964 9580
rect 14004 9392 14056 9444
rect 21732 9528 21784 9580
rect 26240 9528 26292 9580
rect 15660 9503 15712 9512
rect 15660 9469 15669 9503
rect 15669 9469 15703 9503
rect 15703 9469 15712 9503
rect 15660 9460 15712 9469
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 17132 9460 17184 9512
rect 17868 9460 17920 9512
rect 17960 9392 18012 9444
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 17132 9324 17184 9376
rect 18236 9324 18288 9376
rect 22560 9392 22612 9444
rect 21364 9324 21416 9376
rect 23204 9460 23256 9512
rect 23572 9460 23624 9512
rect 23940 9460 23992 9512
rect 26700 9460 26752 9512
rect 27712 9528 27764 9580
rect 32404 9571 32456 9580
rect 32404 9537 32413 9571
rect 32413 9537 32447 9571
rect 32447 9537 32456 9571
rect 32404 9528 32456 9537
rect 33140 9571 33192 9580
rect 27344 9460 27396 9512
rect 28080 9460 28132 9512
rect 29920 9503 29972 9512
rect 29920 9469 29929 9503
rect 29929 9469 29963 9503
rect 29963 9469 29972 9503
rect 29920 9460 29972 9469
rect 33140 9537 33149 9571
rect 33149 9537 33183 9571
rect 33183 9537 33192 9571
rect 33140 9528 33192 9537
rect 36084 9392 36136 9444
rect 29092 9324 29144 9376
rect 29184 9324 29236 9376
rect 30656 9324 30708 9376
rect 30932 9367 30984 9376
rect 30932 9333 30941 9367
rect 30941 9333 30975 9367
rect 30975 9333 30984 9367
rect 30932 9324 30984 9333
rect 33048 9367 33100 9376
rect 33048 9333 33057 9367
rect 33057 9333 33091 9367
rect 33091 9333 33100 9367
rect 33048 9324 33100 9333
rect 33600 9367 33652 9376
rect 33600 9333 33609 9367
rect 33609 9333 33643 9367
rect 33643 9333 33652 9367
rect 33600 9324 33652 9333
rect 37556 9367 37608 9376
rect 37556 9333 37565 9367
rect 37565 9333 37599 9367
rect 37599 9333 37608 9367
rect 37556 9324 37608 9333
rect 38292 9367 38344 9376
rect 38292 9333 38301 9367
rect 38301 9333 38335 9367
rect 38335 9333 38344 9367
rect 38292 9324 38344 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 13728 9120 13780 9172
rect 20628 9120 20680 9172
rect 17868 9052 17920 9104
rect 17960 9052 18012 9104
rect 19708 9052 19760 9104
rect 19984 9052 20036 9104
rect 20996 9052 21048 9104
rect 22100 9120 22152 9172
rect 22652 9120 22704 9172
rect 23204 9052 23256 9104
rect 26608 9120 26660 9172
rect 26700 9120 26752 9172
rect 4068 8984 4120 9036
rect 15936 8984 15988 9036
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 18696 9027 18748 9036
rect 18696 8993 18705 9027
rect 18705 8993 18739 9027
rect 18739 8993 18748 9027
rect 18696 8984 18748 8993
rect 21180 8984 21232 9036
rect 21364 8984 21416 9036
rect 23480 8984 23532 9036
rect 24032 8984 24084 9036
rect 27344 9052 27396 9104
rect 29368 9120 29420 9172
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 12440 8916 12492 8968
rect 15292 8916 15344 8968
rect 14004 8848 14056 8900
rect 15568 8891 15620 8900
rect 15568 8857 15577 8891
rect 15577 8857 15611 8891
rect 15611 8857 15620 8891
rect 15568 8848 15620 8857
rect 16488 8848 16540 8900
rect 16856 8848 16908 8900
rect 18236 8891 18288 8900
rect 18236 8857 18245 8891
rect 18245 8857 18279 8891
rect 18279 8857 18288 8891
rect 18236 8848 18288 8857
rect 18328 8891 18380 8900
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 19340 8848 19392 8900
rect 16580 8780 16632 8832
rect 17316 8780 17368 8832
rect 19708 8848 19760 8900
rect 20996 8848 21048 8900
rect 24308 8916 24360 8968
rect 29920 8984 29972 9036
rect 32772 9052 32824 9104
rect 30932 8984 30984 9036
rect 31576 9027 31628 9036
rect 31576 8993 31585 9027
rect 31585 8993 31619 9027
rect 31619 8993 31628 9027
rect 31576 8984 31628 8993
rect 36084 8959 36136 8968
rect 21088 8780 21140 8832
rect 21548 8848 21600 8900
rect 22560 8848 22612 8900
rect 22928 8780 22980 8832
rect 23204 8780 23256 8832
rect 24584 8780 24636 8832
rect 24860 8848 24912 8900
rect 26240 8848 26292 8900
rect 36084 8925 36093 8959
rect 36093 8925 36127 8959
rect 36127 8925 36136 8959
rect 36084 8916 36136 8925
rect 37556 8959 37608 8968
rect 37556 8925 37565 8959
rect 37565 8925 37599 8959
rect 37599 8925 37608 8959
rect 37556 8916 37608 8925
rect 25504 8780 25556 8832
rect 28356 8848 28408 8900
rect 29184 8848 29236 8900
rect 29644 8848 29696 8900
rect 30564 8848 30616 8900
rect 31300 8891 31352 8900
rect 31300 8857 31309 8891
rect 31309 8857 31343 8891
rect 31343 8857 31352 8891
rect 31300 8848 31352 8857
rect 32588 8891 32640 8900
rect 32588 8857 32597 8891
rect 32597 8857 32631 8891
rect 32631 8857 32640 8891
rect 32588 8848 32640 8857
rect 33600 8848 33652 8900
rect 35992 8891 36044 8900
rect 35992 8857 36001 8891
rect 36001 8857 36035 8891
rect 36035 8857 36044 8891
rect 35992 8848 36044 8857
rect 26608 8780 26660 8832
rect 30288 8780 30340 8832
rect 30932 8780 30984 8832
rect 32128 8780 32180 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 15292 8576 15344 8628
rect 15844 8576 15896 8628
rect 17224 8576 17276 8628
rect 13912 8551 13964 8560
rect 13912 8517 13921 8551
rect 13921 8517 13955 8551
rect 13955 8517 13964 8551
rect 13912 8508 13964 8517
rect 14648 8440 14700 8492
rect 17592 8508 17644 8560
rect 17132 8483 17184 8492
rect 14832 8372 14884 8424
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17868 8508 17920 8560
rect 20812 8576 20864 8628
rect 21640 8576 21692 8628
rect 23296 8576 23348 8628
rect 25596 8576 25648 8628
rect 27712 8576 27764 8628
rect 19340 8508 19392 8560
rect 20720 8508 20772 8560
rect 21088 8508 21140 8560
rect 21732 8508 21784 8560
rect 22192 8508 22244 8560
rect 23664 8508 23716 8560
rect 25044 8508 25096 8560
rect 20352 8440 20404 8492
rect 20628 8440 20680 8492
rect 22284 8440 22336 8492
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 17684 8372 17736 8424
rect 13636 8304 13688 8356
rect 14096 8304 14148 8356
rect 17132 8304 17184 8356
rect 19616 8372 19668 8424
rect 20168 8372 20220 8424
rect 21456 8372 21508 8424
rect 21732 8372 21784 8424
rect 21916 8372 21968 8424
rect 24676 8372 24728 8424
rect 29552 8508 29604 8560
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 29368 8440 29420 8492
rect 26884 8372 26936 8424
rect 27528 8372 27580 8424
rect 29276 8372 29328 8424
rect 30564 8508 30616 8560
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 36820 8440 36872 8492
rect 19156 8347 19208 8356
rect 2044 8236 2096 8288
rect 6828 8236 6880 8288
rect 15016 8236 15068 8288
rect 19156 8313 19165 8347
rect 19165 8313 19199 8347
rect 19199 8313 19208 8347
rect 19156 8304 19208 8313
rect 19340 8304 19392 8356
rect 22560 8304 22612 8356
rect 19248 8236 19300 8288
rect 20628 8236 20680 8288
rect 21456 8236 21508 8288
rect 25780 8236 25832 8288
rect 25872 8236 25924 8288
rect 28632 8236 28684 8288
rect 28724 8236 28776 8288
rect 29552 8304 29604 8356
rect 29276 8236 29328 8288
rect 29736 8236 29788 8288
rect 37188 8372 37240 8424
rect 30840 8304 30892 8356
rect 31576 8304 31628 8356
rect 32588 8304 32640 8356
rect 34520 8304 34572 8356
rect 36360 8347 36412 8356
rect 36360 8313 36369 8347
rect 36369 8313 36403 8347
rect 36403 8313 36412 8347
rect 36360 8304 36412 8313
rect 33600 8236 33652 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 18144 8032 18196 8084
rect 19064 8032 19116 8084
rect 19616 8032 19668 8084
rect 20168 8032 20220 8084
rect 20720 8075 20772 8084
rect 20720 8041 20729 8075
rect 20729 8041 20763 8075
rect 20763 8041 20772 8075
rect 20720 8032 20772 8041
rect 21916 8032 21968 8084
rect 22008 8032 22060 8084
rect 24308 8032 24360 8084
rect 16580 7964 16632 8016
rect 15200 7896 15252 7948
rect 16396 7896 16448 7948
rect 18880 7964 18932 8016
rect 17776 7939 17828 7948
rect 17776 7905 17785 7939
rect 17785 7905 17819 7939
rect 17819 7905 17828 7939
rect 17776 7896 17828 7905
rect 18420 7896 18472 7948
rect 18788 7896 18840 7948
rect 21456 7896 21508 7948
rect 23480 7896 23532 7948
rect 12440 7828 12492 7880
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15292 7828 15344 7880
rect 19248 7828 19300 7880
rect 21180 7828 21232 7880
rect 24032 7871 24084 7880
rect 24032 7837 24041 7871
rect 24041 7837 24075 7871
rect 24075 7837 24084 7871
rect 24032 7828 24084 7837
rect 28264 8032 28316 8084
rect 31208 7964 31260 8016
rect 36084 8032 36136 8084
rect 27528 7896 27580 7948
rect 26700 7871 26752 7880
rect 26700 7837 26709 7871
rect 26709 7837 26743 7871
rect 26743 7837 26752 7871
rect 30380 7896 30432 7948
rect 36636 7939 36688 7948
rect 26700 7828 26752 7837
rect 36636 7905 36645 7939
rect 36645 7905 36679 7939
rect 36679 7905 36688 7939
rect 36636 7896 36688 7905
rect 36084 7828 36136 7880
rect 37832 7871 37884 7880
rect 37832 7837 37841 7871
rect 37841 7837 37875 7871
rect 37875 7837 37884 7871
rect 37832 7828 37884 7837
rect 13452 7692 13504 7744
rect 14556 7760 14608 7812
rect 16120 7760 16172 7812
rect 16396 7760 16448 7812
rect 14648 7692 14700 7744
rect 18788 7760 18840 7812
rect 19984 7803 20036 7812
rect 19984 7769 19993 7803
rect 19993 7769 20027 7803
rect 20027 7769 20036 7803
rect 19984 7760 20036 7769
rect 22652 7760 22704 7812
rect 23020 7760 23072 7812
rect 18144 7692 18196 7744
rect 20812 7692 20864 7744
rect 20904 7692 20956 7744
rect 21640 7692 21692 7744
rect 22744 7692 22796 7744
rect 25044 7760 25096 7812
rect 26332 7760 26384 7812
rect 28632 7760 28684 7812
rect 29460 7760 29512 7812
rect 31300 7760 31352 7812
rect 26240 7692 26292 7744
rect 31484 7692 31536 7744
rect 31944 7735 31996 7744
rect 31944 7701 31953 7735
rect 31953 7701 31987 7735
rect 31987 7701 31996 7735
rect 31944 7692 31996 7701
rect 33416 7692 33468 7744
rect 37464 7692 37516 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 14648 7488 14700 7540
rect 16396 7488 16448 7540
rect 16580 7488 16632 7540
rect 19156 7488 19208 7540
rect 19616 7488 19668 7540
rect 26332 7488 26384 7540
rect 26884 7488 26936 7540
rect 2044 7420 2096 7472
rect 15292 7420 15344 7472
rect 1584 7352 1636 7404
rect 12440 7352 12492 7404
rect 13820 7352 13872 7404
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 16672 7420 16724 7472
rect 16948 7463 17000 7472
rect 16948 7429 16957 7463
rect 16957 7429 16991 7463
rect 16991 7429 17000 7463
rect 16948 7420 17000 7429
rect 17132 7420 17184 7472
rect 19340 7420 19392 7472
rect 20168 7420 20220 7472
rect 23480 7420 23532 7472
rect 23848 7420 23900 7472
rect 24492 7463 24544 7472
rect 16028 7352 16080 7404
rect 16396 7352 16448 7404
rect 17592 7352 17644 7404
rect 19800 7352 19852 7404
rect 21272 7352 21324 7404
rect 21456 7352 21508 7404
rect 24492 7429 24501 7463
rect 24501 7429 24535 7463
rect 24535 7429 24544 7463
rect 24492 7420 24544 7429
rect 27252 7420 27304 7472
rect 28356 7488 28408 7540
rect 30656 7488 30708 7540
rect 34796 7488 34848 7540
rect 35532 7488 35584 7540
rect 36084 7488 36136 7540
rect 29000 7420 29052 7472
rect 29552 7420 29604 7472
rect 33140 7420 33192 7472
rect 37556 7420 37608 7472
rect 19524 7284 19576 7336
rect 19892 7284 19944 7336
rect 20168 7284 20220 7336
rect 22100 7284 22152 7336
rect 26792 7352 26844 7404
rect 27160 7395 27212 7404
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 38200 7352 38252 7404
rect 23664 7284 23716 7336
rect 25872 7284 25924 7336
rect 26240 7327 26292 7336
rect 26240 7293 26249 7327
rect 26249 7293 26283 7327
rect 26283 7293 26292 7327
rect 26240 7284 26292 7293
rect 26608 7284 26660 7336
rect 16672 7216 16724 7268
rect 17040 7216 17092 7268
rect 17776 7216 17828 7268
rect 12808 7148 12860 7200
rect 16120 7148 16172 7200
rect 18880 7216 18932 7268
rect 19248 7216 19300 7268
rect 21180 7216 21232 7268
rect 22468 7216 22520 7268
rect 27436 7216 27488 7268
rect 27528 7216 27580 7268
rect 31944 7284 31996 7336
rect 34612 7284 34664 7336
rect 34704 7284 34756 7336
rect 19616 7148 19668 7200
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 21088 7148 21140 7200
rect 21364 7191 21416 7200
rect 21364 7157 21373 7191
rect 21373 7157 21407 7191
rect 21407 7157 21416 7191
rect 21364 7148 21416 7157
rect 29000 7148 29052 7200
rect 30656 7216 30708 7268
rect 31576 7216 31628 7268
rect 32036 7216 32088 7268
rect 33416 7259 33468 7268
rect 33416 7225 33425 7259
rect 33425 7225 33459 7259
rect 33459 7225 33468 7259
rect 33416 7216 33468 7225
rect 35624 7216 35676 7268
rect 30840 7191 30892 7200
rect 30840 7157 30849 7191
rect 30849 7157 30883 7191
rect 30883 7157 30892 7191
rect 30840 7148 30892 7157
rect 32680 7148 32732 7200
rect 35716 7191 35768 7200
rect 35716 7157 35725 7191
rect 35725 7157 35759 7191
rect 35759 7157 35768 7191
rect 35716 7148 35768 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 14280 6944 14332 6996
rect 15016 6944 15068 6996
rect 26240 6944 26292 6996
rect 12808 6876 12860 6928
rect 15660 6808 15712 6860
rect 16212 6808 16264 6860
rect 16856 6808 16908 6860
rect 17960 6808 18012 6860
rect 18604 6808 18656 6860
rect 19248 6808 19300 6860
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 13360 6740 13412 6792
rect 13820 6740 13872 6792
rect 14188 6740 14240 6792
rect 15384 6740 15436 6792
rect 16120 6740 16172 6792
rect 16948 6740 17000 6792
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 18052 6740 18104 6792
rect 18972 6740 19024 6792
rect 20720 6876 20772 6928
rect 23388 6919 23440 6928
rect 20904 6808 20956 6860
rect 21364 6808 21416 6860
rect 23388 6885 23397 6919
rect 23397 6885 23431 6919
rect 23431 6885 23440 6919
rect 23388 6876 23440 6885
rect 23664 6876 23716 6928
rect 29000 6944 29052 6996
rect 29092 6944 29144 6996
rect 31484 6987 31536 6996
rect 31484 6953 31493 6987
rect 31493 6953 31527 6987
rect 31527 6953 31536 6987
rect 31484 6944 31536 6953
rect 32036 6987 32088 6996
rect 32036 6953 32045 6987
rect 32045 6953 32079 6987
rect 32079 6953 32088 6987
rect 32036 6944 32088 6953
rect 36084 6944 36136 6996
rect 37832 6944 37884 6996
rect 38200 6987 38252 6996
rect 38200 6953 38209 6987
rect 38209 6953 38243 6987
rect 38243 6953 38252 6987
rect 38200 6944 38252 6953
rect 24952 6808 25004 6860
rect 25504 6851 25556 6860
rect 25504 6817 25513 6851
rect 25513 6817 25547 6851
rect 25547 6817 25556 6851
rect 25504 6808 25556 6817
rect 24032 6783 24084 6792
rect 13636 6715 13688 6724
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 17040 6672 17092 6724
rect 19340 6672 19392 6724
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 19800 6672 19852 6724
rect 21548 6672 21600 6724
rect 21640 6672 21692 6724
rect 23940 6715 23992 6724
rect 20720 6604 20772 6656
rect 20996 6604 21048 6656
rect 23940 6681 23949 6715
rect 23949 6681 23983 6715
rect 23983 6681 23992 6715
rect 23940 6672 23992 6681
rect 25136 6740 25188 6792
rect 26056 6672 26108 6724
rect 26608 6808 26660 6860
rect 27160 6808 27212 6860
rect 31576 6808 31628 6860
rect 34612 6808 34664 6860
rect 35440 6851 35492 6860
rect 35440 6817 35449 6851
rect 35449 6817 35483 6851
rect 35483 6817 35492 6851
rect 35440 6808 35492 6817
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 30288 6672 30340 6724
rect 30472 6672 30524 6724
rect 24492 6604 24544 6656
rect 27988 6647 28040 6656
rect 27988 6613 27997 6647
rect 27997 6613 28031 6647
rect 28031 6613 28040 6647
rect 27988 6604 28040 6613
rect 32496 6604 32548 6656
rect 33416 6604 33468 6656
rect 33692 6604 33744 6656
rect 35808 6604 35860 6656
rect 36636 6647 36688 6656
rect 36636 6613 36645 6647
rect 36645 6613 36679 6647
rect 36679 6613 36688 6647
rect 36636 6604 36688 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 12532 6400 12584 6452
rect 13452 6400 13504 6452
rect 13912 6400 13964 6452
rect 16580 6400 16632 6452
rect 16948 6400 17000 6452
rect 19340 6400 19392 6452
rect 19984 6400 20036 6452
rect 22284 6400 22336 6452
rect 15752 6375 15804 6384
rect 15752 6341 15761 6375
rect 15761 6341 15795 6375
rect 15795 6341 15804 6375
rect 18328 6375 18380 6384
rect 15752 6332 15804 6341
rect 18328 6341 18337 6375
rect 18337 6341 18371 6375
rect 18371 6341 18380 6375
rect 18328 6332 18380 6341
rect 18420 6332 18472 6384
rect 20076 6332 20128 6384
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13360 6264 13412 6316
rect 14464 6264 14516 6316
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 15384 6196 15436 6248
rect 16672 6196 16724 6248
rect 17684 6196 17736 6248
rect 19432 6196 19484 6248
rect 16028 6128 16080 6180
rect 14280 6060 14332 6112
rect 18788 6128 18840 6180
rect 16856 6060 16908 6112
rect 22100 6332 22152 6384
rect 23664 6332 23716 6384
rect 20352 6307 20404 6316
rect 20352 6273 20361 6307
rect 20361 6273 20395 6307
rect 20395 6273 20404 6307
rect 20352 6264 20404 6273
rect 20444 6264 20496 6316
rect 23848 6307 23900 6316
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 20812 6196 20864 6248
rect 23020 6196 23072 6248
rect 23480 6196 23532 6248
rect 24676 6264 24728 6316
rect 24584 6239 24636 6248
rect 24584 6205 24593 6239
rect 24593 6205 24627 6239
rect 24627 6205 24636 6239
rect 24584 6196 24636 6205
rect 24860 6332 24912 6384
rect 26056 6400 26108 6452
rect 26516 6400 26568 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 28448 6400 28500 6452
rect 28816 6400 28868 6452
rect 29368 6332 29420 6384
rect 29828 6332 29880 6384
rect 30012 6332 30064 6384
rect 31576 6332 31628 6384
rect 33600 6400 33652 6452
rect 38016 6375 38068 6384
rect 38016 6341 38025 6375
rect 38025 6341 38059 6375
rect 38059 6341 38068 6375
rect 38016 6332 38068 6341
rect 26240 6196 26292 6248
rect 26608 6239 26660 6248
rect 26608 6205 26617 6239
rect 26617 6205 26651 6239
rect 26651 6205 26660 6239
rect 26608 6196 26660 6205
rect 23940 6128 23992 6180
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 21732 6060 21784 6112
rect 24860 6060 24912 6112
rect 30288 6264 30340 6316
rect 30564 6264 30616 6316
rect 34060 6264 34112 6316
rect 35440 6307 35492 6316
rect 35440 6273 35449 6307
rect 35449 6273 35483 6307
rect 35483 6273 35492 6307
rect 35440 6264 35492 6273
rect 38200 6307 38252 6316
rect 38200 6273 38209 6307
rect 38209 6273 38243 6307
rect 38243 6273 38252 6307
rect 38200 6264 38252 6273
rect 29736 6239 29788 6248
rect 29736 6205 29745 6239
rect 29745 6205 29779 6239
rect 29779 6205 29788 6239
rect 29736 6196 29788 6205
rect 31944 6196 31996 6248
rect 31576 6128 31628 6180
rect 33140 6128 33192 6180
rect 33416 6171 33468 6180
rect 33416 6137 33425 6171
rect 33425 6137 33459 6171
rect 33459 6137 33468 6171
rect 33416 6128 33468 6137
rect 29276 6060 29328 6112
rect 30380 6060 30432 6112
rect 32496 6060 32548 6112
rect 34520 6103 34572 6112
rect 34520 6069 34529 6103
rect 34529 6069 34563 6103
rect 34563 6069 34572 6103
rect 34520 6060 34572 6069
rect 35348 6103 35400 6112
rect 35348 6069 35357 6103
rect 35357 6069 35391 6103
rect 35391 6069 35400 6103
rect 35348 6060 35400 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 13268 5856 13320 5908
rect 13728 5856 13780 5908
rect 15384 5856 15436 5908
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 16028 5856 16080 5908
rect 16856 5856 16908 5908
rect 20168 5856 20220 5908
rect 20352 5856 20404 5908
rect 14740 5788 14792 5840
rect 15936 5788 15988 5840
rect 16672 5788 16724 5840
rect 17592 5831 17644 5840
rect 17592 5797 17601 5831
rect 17601 5797 17635 5831
rect 17635 5797 17644 5831
rect 17592 5788 17644 5797
rect 17684 5788 17736 5840
rect 13636 5652 13688 5704
rect 14464 5652 14516 5704
rect 17960 5720 18012 5772
rect 18144 5788 18196 5840
rect 20628 5788 20680 5840
rect 20812 5831 20864 5840
rect 20812 5797 20821 5831
rect 20821 5797 20855 5831
rect 20855 5797 20864 5831
rect 20812 5788 20864 5797
rect 20996 5788 21048 5840
rect 21364 5788 21416 5840
rect 24032 5856 24084 5908
rect 31576 5856 31628 5908
rect 31668 5856 31720 5908
rect 24400 5788 24452 5840
rect 26332 5831 26384 5840
rect 26332 5797 26341 5831
rect 26341 5797 26375 5831
rect 26375 5797 26384 5831
rect 26332 5788 26384 5797
rect 28908 5831 28960 5840
rect 28908 5797 28917 5831
rect 28917 5797 28951 5831
rect 28951 5797 28960 5831
rect 28908 5788 28960 5797
rect 31392 5788 31444 5840
rect 19156 5720 19208 5772
rect 23664 5720 23716 5772
rect 23848 5720 23900 5772
rect 24860 5763 24912 5772
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 24952 5720 25004 5772
rect 29736 5763 29788 5772
rect 29736 5729 29745 5763
rect 29745 5729 29779 5763
rect 29779 5729 29788 5763
rect 29736 5720 29788 5729
rect 30012 5763 30064 5772
rect 30012 5729 30021 5763
rect 30021 5729 30055 5763
rect 30055 5729 30064 5763
rect 30012 5720 30064 5729
rect 31024 5720 31076 5772
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16212 5627 16264 5636
rect 16212 5593 16221 5627
rect 16221 5593 16255 5627
rect 16255 5593 16264 5627
rect 16212 5584 16264 5593
rect 16580 5584 16632 5636
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 24032 5695 24084 5704
rect 19156 5584 19208 5636
rect 20904 5584 20956 5636
rect 21272 5584 21324 5636
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 26332 5652 26384 5704
rect 26608 5652 26660 5704
rect 21548 5584 21600 5636
rect 21916 5584 21968 5636
rect 22376 5584 22428 5636
rect 23204 5584 23256 5636
rect 25320 5584 25372 5636
rect 28724 5584 28776 5636
rect 31944 5763 31996 5772
rect 31944 5729 31953 5763
rect 31953 5729 31987 5763
rect 31987 5729 31996 5763
rect 31944 5720 31996 5729
rect 35624 5856 35676 5908
rect 37096 5899 37148 5908
rect 37096 5865 37105 5899
rect 37105 5865 37139 5899
rect 37139 5865 37148 5899
rect 37096 5856 37148 5865
rect 38108 5856 38160 5908
rect 34520 5788 34572 5840
rect 35808 5788 35860 5840
rect 34060 5720 34112 5772
rect 9220 5516 9272 5568
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 18788 5516 18840 5568
rect 20444 5516 20496 5568
rect 20536 5516 20588 5568
rect 22652 5516 22704 5568
rect 23296 5516 23348 5568
rect 24400 5516 24452 5568
rect 31024 5516 31076 5568
rect 34704 5584 34756 5636
rect 34796 5516 34848 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 14096 5312 14148 5364
rect 15752 5312 15804 5364
rect 16948 5355 17000 5364
rect 16948 5321 16957 5355
rect 16957 5321 16991 5355
rect 16991 5321 17000 5355
rect 16948 5312 17000 5321
rect 18144 5312 18196 5364
rect 23756 5355 23808 5364
rect 17132 5244 17184 5296
rect 18052 5244 18104 5296
rect 18696 5244 18748 5296
rect 18972 5244 19024 5296
rect 20812 5244 20864 5296
rect 20904 5244 20956 5296
rect 23756 5321 23765 5355
rect 23765 5321 23799 5355
rect 23799 5321 23808 5355
rect 23756 5312 23808 5321
rect 23848 5312 23900 5364
rect 24952 5312 25004 5364
rect 25044 5312 25096 5364
rect 30012 5355 30064 5364
rect 10324 5176 10376 5228
rect 12440 5176 12492 5228
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 16028 5219 16080 5228
rect 15200 5108 15252 5160
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 19248 5176 19300 5228
rect 18236 5108 18288 5160
rect 20444 5108 20496 5160
rect 17684 5040 17736 5092
rect 17960 5083 18012 5092
rect 17960 5049 17969 5083
rect 17969 5049 18003 5083
rect 18003 5049 18012 5083
rect 17960 5040 18012 5049
rect 18788 5040 18840 5092
rect 19984 5040 20036 5092
rect 21180 5176 21232 5228
rect 21364 5176 21416 5228
rect 24492 5176 24544 5228
rect 26332 5244 26384 5296
rect 26608 5287 26660 5296
rect 26608 5253 26617 5287
rect 26617 5253 26651 5287
rect 26651 5253 26660 5287
rect 26608 5244 26660 5253
rect 28080 5244 28132 5296
rect 30012 5321 30021 5355
rect 30021 5321 30055 5355
rect 30055 5321 30064 5355
rect 30012 5312 30064 5321
rect 34612 5312 34664 5364
rect 35808 5312 35860 5364
rect 37924 5244 37976 5296
rect 27344 5219 27396 5228
rect 22008 5151 22060 5160
rect 22008 5117 22017 5151
rect 22017 5117 22051 5151
rect 22051 5117 22060 5151
rect 22008 5108 22060 5117
rect 24584 5108 24636 5160
rect 25136 5108 25188 5160
rect 23756 5040 23808 5092
rect 27344 5185 27353 5219
rect 27353 5185 27387 5219
rect 27387 5185 27396 5219
rect 27344 5176 27396 5185
rect 26332 5108 26384 5160
rect 29184 5108 29236 5160
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 18236 4972 18288 5024
rect 18696 4972 18748 5024
rect 21180 4972 21232 5024
rect 22744 4972 22796 5024
rect 22836 4972 22888 5024
rect 30104 5176 30156 5228
rect 31484 5176 31536 5228
rect 32496 5219 32548 5228
rect 32496 5185 32505 5219
rect 32505 5185 32539 5219
rect 32539 5185 32548 5219
rect 32496 5176 32548 5185
rect 36636 5176 36688 5228
rect 38200 5219 38252 5228
rect 38200 5185 38209 5219
rect 38209 5185 38243 5219
rect 38243 5185 38252 5219
rect 38200 5176 38252 5185
rect 30380 5108 30432 5160
rect 30564 5108 30616 5160
rect 32312 5040 32364 5092
rect 32128 4972 32180 5024
rect 32772 4972 32824 5024
rect 32864 4972 32916 5024
rect 34796 4972 34848 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10324 4811 10376 4820
rect 10324 4777 10333 4811
rect 10333 4777 10367 4811
rect 10367 4777 10376 4811
rect 10324 4768 10376 4777
rect 18144 4768 18196 4820
rect 18420 4768 18472 4820
rect 18696 4768 18748 4820
rect 21916 4768 21968 4820
rect 22100 4768 22152 4820
rect 23940 4768 23992 4820
rect 24768 4768 24820 4820
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 15936 4632 15988 4684
rect 16856 4632 16908 4684
rect 17500 4700 17552 4752
rect 17592 4700 17644 4752
rect 20904 4700 20956 4752
rect 21640 4700 21692 4752
rect 30656 4768 30708 4820
rect 33232 4768 33284 4820
rect 17316 4632 17368 4684
rect 18972 4632 19024 4684
rect 20260 4632 20312 4684
rect 21272 4632 21324 4684
rect 22008 4632 22060 4684
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 13636 4564 13688 4616
rect 15660 4601 15712 4616
rect 15660 4567 15677 4601
rect 15677 4567 15711 4601
rect 15711 4567 15712 4601
rect 15660 4564 15712 4567
rect 14096 4428 14148 4480
rect 14648 4428 14700 4480
rect 16580 4428 16632 4480
rect 17224 4428 17276 4480
rect 17316 4428 17368 4480
rect 17960 4496 18012 4548
rect 19248 4564 19300 4616
rect 20720 4564 20772 4616
rect 17776 4428 17828 4480
rect 18880 4428 18932 4480
rect 19432 4428 19484 4480
rect 22560 4496 22612 4548
rect 25964 4632 26016 4684
rect 26424 4632 26476 4684
rect 32680 4700 32732 4752
rect 31392 4632 31444 4684
rect 23848 4564 23900 4616
rect 24952 4564 25004 4616
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 26332 4564 26384 4573
rect 29000 4564 29052 4616
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 31300 4564 31352 4616
rect 23940 4471 23992 4480
rect 23940 4437 23949 4471
rect 23949 4437 23983 4471
rect 23983 4437 23992 4471
rect 23940 4428 23992 4437
rect 25044 4428 25096 4480
rect 26240 4428 26292 4480
rect 28908 4496 28960 4548
rect 32312 4607 32364 4616
rect 32312 4573 32321 4607
rect 32321 4573 32355 4607
rect 32355 4573 32364 4607
rect 32312 4564 32364 4573
rect 33324 4632 33376 4684
rect 34060 4564 34112 4616
rect 34520 4564 34572 4616
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 33416 4496 33468 4548
rect 36084 4496 36136 4548
rect 31576 4428 31628 4480
rect 33508 4428 33560 4480
rect 34152 4471 34204 4480
rect 34152 4437 34161 4471
rect 34161 4437 34195 4471
rect 34195 4437 34204 4471
rect 34152 4428 34204 4437
rect 34888 4471 34940 4480
rect 34888 4437 34897 4471
rect 34897 4437 34931 4471
rect 34931 4437 34940 4471
rect 34888 4428 34940 4437
rect 36268 4428 36320 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 14648 4199 14700 4208
rect 14648 4165 14657 4199
rect 14657 4165 14691 4199
rect 14691 4165 14700 4199
rect 14648 4156 14700 4165
rect 9956 4088 10008 4140
rect 14096 4088 14148 4140
rect 14464 4088 14516 4140
rect 15660 4156 15712 4208
rect 16488 4156 16540 4208
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 17040 4224 17092 4276
rect 17960 4156 18012 4208
rect 19984 4224 20036 4276
rect 22100 4224 22152 4276
rect 22192 4267 22244 4276
rect 22192 4233 22201 4267
rect 22201 4233 22235 4267
rect 22235 4233 22244 4267
rect 22192 4224 22244 4233
rect 25044 4224 25096 4276
rect 25136 4224 25188 4276
rect 28724 4224 28776 4276
rect 23940 4156 23992 4208
rect 24400 4199 24452 4208
rect 24400 4165 24409 4199
rect 24409 4165 24443 4199
rect 24443 4165 24452 4199
rect 24400 4156 24452 4165
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18972 4131 19024 4140
rect 18144 4020 18196 4072
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19616 4088 19668 4140
rect 23112 4088 23164 4140
rect 26332 4156 26384 4208
rect 26608 4199 26660 4208
rect 26608 4165 26617 4199
rect 26617 4165 26651 4199
rect 26651 4165 26660 4199
rect 26608 4156 26660 4165
rect 32864 4224 32916 4276
rect 33416 4267 33468 4276
rect 33416 4233 33425 4267
rect 33425 4233 33459 4267
rect 33459 4233 33468 4267
rect 33416 4224 33468 4233
rect 34060 4224 34112 4276
rect 37372 4224 37424 4276
rect 36268 4156 36320 4208
rect 25872 4088 25924 4140
rect 24676 4063 24728 4072
rect 24676 4029 24685 4063
rect 24685 4029 24719 4063
rect 24719 4029 24728 4063
rect 24676 4020 24728 4029
rect 25136 4020 25188 4072
rect 13912 3952 13964 4004
rect 19432 3952 19484 4004
rect 21272 3952 21324 4004
rect 18052 3884 18104 3936
rect 18236 3884 18288 3936
rect 20536 3884 20588 3936
rect 20904 3884 20956 3936
rect 22100 3952 22152 4004
rect 22284 3952 22336 4004
rect 24768 3952 24820 4004
rect 25872 3952 25924 4004
rect 25964 3952 26016 4004
rect 27344 4020 27396 4072
rect 29000 4088 29052 4140
rect 31484 4088 31536 4140
rect 33232 4088 33284 4140
rect 29368 4063 29420 4072
rect 29368 4029 29377 4063
rect 29377 4029 29411 4063
rect 29411 4029 29420 4063
rect 29368 4020 29420 4029
rect 31208 4020 31260 4072
rect 32128 4020 32180 4072
rect 21456 3927 21508 3936
rect 21456 3893 21465 3927
rect 21465 3893 21499 3927
rect 21499 3893 21508 3927
rect 21456 3884 21508 3893
rect 24032 3884 24084 3936
rect 31668 3952 31720 4004
rect 31944 3952 31996 4004
rect 37832 4088 37884 4140
rect 37556 4020 37608 4072
rect 38108 4020 38160 4072
rect 34336 3952 34388 4004
rect 36636 3952 36688 4004
rect 28448 3884 28500 3936
rect 28632 3927 28684 3936
rect 28632 3893 28653 3927
rect 28653 3893 28684 3927
rect 28632 3884 28684 3893
rect 31116 3884 31168 3936
rect 31484 3884 31536 3936
rect 33508 3884 33560 3936
rect 33876 3927 33928 3936
rect 33876 3893 33885 3927
rect 33885 3893 33919 3927
rect 33919 3893 33928 3927
rect 33876 3884 33928 3893
rect 34888 3884 34940 3936
rect 36084 3927 36136 3936
rect 36084 3893 36093 3927
rect 36093 3893 36127 3927
rect 36127 3893 36136 3927
rect 36084 3884 36136 3893
rect 38200 3927 38252 3936
rect 38200 3893 38209 3927
rect 38209 3893 38243 3927
rect 38243 3893 38252 3927
rect 38200 3884 38252 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 14096 3680 14148 3732
rect 17224 3680 17276 3732
rect 17684 3680 17736 3732
rect 19432 3680 19484 3732
rect 19616 3723 19668 3732
rect 19616 3689 19625 3723
rect 19625 3689 19659 3723
rect 19659 3689 19668 3723
rect 19616 3680 19668 3689
rect 19892 3680 19944 3732
rect 21916 3680 21968 3732
rect 22192 3680 22244 3732
rect 28448 3680 28500 3732
rect 31576 3680 31628 3732
rect 31668 3680 31720 3732
rect 33876 3680 33928 3732
rect 15936 3612 15988 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 12440 3476 12492 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 16488 3544 16540 3596
rect 18144 3544 18196 3596
rect 20996 3544 21048 3596
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 22928 3612 22980 3664
rect 23112 3612 23164 3664
rect 24952 3612 25004 3664
rect 31116 3612 31168 3664
rect 31760 3612 31812 3664
rect 33232 3612 33284 3664
rect 33692 3655 33744 3664
rect 33692 3621 33701 3655
rect 33701 3621 33735 3655
rect 33735 3621 33744 3655
rect 33692 3612 33744 3621
rect 33968 3612 34020 3664
rect 21640 3544 21692 3596
rect 21916 3544 21968 3596
rect 26332 3587 26384 3596
rect 26332 3553 26341 3587
rect 26341 3553 26375 3587
rect 26375 3553 26384 3587
rect 26332 3544 26384 3553
rect 29736 3587 29788 3596
rect 29736 3553 29745 3587
rect 29745 3553 29779 3587
rect 29779 3553 29788 3587
rect 29736 3544 29788 3553
rect 31208 3544 31260 3596
rect 37372 3612 37424 3664
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 16672 3408 16724 3460
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18696 3451 18748 3460
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 17132 3340 17184 3392
rect 18696 3417 18705 3451
rect 18705 3417 18739 3451
rect 18739 3417 18748 3451
rect 18696 3408 18748 3417
rect 19340 3408 19392 3460
rect 23756 3476 23808 3528
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 37556 3519 37608 3528
rect 37556 3485 37565 3519
rect 37565 3485 37599 3519
rect 37599 3485 37608 3519
rect 37556 3476 37608 3485
rect 38292 3476 38344 3528
rect 39304 3476 39356 3528
rect 22928 3408 22980 3460
rect 23480 3408 23532 3460
rect 25320 3408 25372 3460
rect 25780 3408 25832 3460
rect 19892 3340 19944 3392
rect 19984 3340 20036 3392
rect 23848 3383 23900 3392
rect 23848 3349 23857 3383
rect 23857 3349 23891 3383
rect 23891 3349 23900 3383
rect 23848 3340 23900 3349
rect 24400 3340 24452 3392
rect 26148 3340 26200 3392
rect 26884 3340 26936 3392
rect 31944 3408 31996 3460
rect 32220 3451 32272 3460
rect 32220 3417 32229 3451
rect 32229 3417 32263 3451
rect 32263 3417 32272 3451
rect 32220 3408 32272 3417
rect 34152 3408 34204 3460
rect 34244 3451 34296 3460
rect 34244 3417 34253 3451
rect 34253 3417 34287 3451
rect 34287 3417 34296 3451
rect 34244 3408 34296 3417
rect 36084 3451 36136 3460
rect 36084 3417 36093 3451
rect 36093 3417 36127 3451
rect 36127 3417 36136 3451
rect 36084 3408 36136 3417
rect 31392 3340 31444 3392
rect 31576 3340 31628 3392
rect 33600 3340 33652 3392
rect 33692 3340 33744 3392
rect 36360 3340 36412 3392
rect 37556 3340 37608 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 10048 3136 10100 3188
rect 12992 3136 13044 3188
rect 14280 3068 14332 3120
rect 14464 3068 14516 3120
rect 17132 3111 17184 3120
rect 17132 3077 17141 3111
rect 17141 3077 17175 3111
rect 17175 3077 17184 3111
rect 17132 3068 17184 3077
rect 18236 3068 18288 3120
rect 18604 3068 18656 3120
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 14004 2932 14056 2984
rect 31760 3136 31812 3188
rect 31944 3136 31996 3188
rect 33232 3136 33284 3188
rect 33600 3136 33652 3188
rect 36084 3136 36136 3188
rect 18788 3068 18840 3120
rect 21272 3068 21324 3120
rect 23296 3068 23348 3120
rect 24308 3068 24360 3120
rect 24584 3111 24636 3120
rect 24584 3077 24593 3111
rect 24593 3077 24627 3111
rect 24627 3077 24636 3111
rect 24584 3068 24636 3077
rect 24860 3068 24912 3120
rect 26332 3068 26384 3120
rect 18880 3000 18932 3052
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 27344 3068 27396 3120
rect 28816 3068 28868 3120
rect 29552 3068 29604 3120
rect 31116 3068 31168 3120
rect 31300 3068 31352 3120
rect 36636 3068 36688 3120
rect 21456 3000 21508 3009
rect 27068 3000 27120 3052
rect 28724 3000 28776 3052
rect 15200 2932 15252 2984
rect 12716 2864 12768 2916
rect 16120 2864 16172 2916
rect 16304 2932 16356 2984
rect 22836 2932 22888 2984
rect 26240 2932 26292 2984
rect 26700 2932 26752 2984
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 7564 2796 7616 2848
rect 12440 2796 12492 2848
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 15476 2796 15528 2848
rect 16212 2839 16264 2848
rect 16212 2805 16221 2839
rect 16221 2805 16255 2839
rect 16255 2805 16264 2839
rect 16212 2796 16264 2805
rect 17500 2864 17552 2916
rect 17776 2864 17828 2916
rect 19432 2796 19484 2848
rect 24952 2864 25004 2916
rect 28632 2932 28684 2984
rect 28908 2932 28960 2984
rect 29644 2932 29696 2984
rect 35532 3000 35584 3052
rect 36360 3000 36412 3052
rect 31300 2932 31352 2984
rect 21364 2796 21416 2848
rect 22284 2839 22336 2848
rect 22284 2805 22314 2839
rect 22314 2805 22336 2839
rect 22284 2796 22336 2805
rect 29000 2864 29052 2916
rect 30380 2864 30432 2916
rect 32128 2932 32180 2984
rect 31760 2864 31812 2916
rect 31852 2864 31904 2916
rect 35348 2932 35400 2984
rect 26700 2796 26752 2848
rect 34152 2796 34204 2848
rect 37556 2839 37608 2848
rect 37556 2805 37565 2839
rect 37565 2805 37599 2839
rect 37599 2805 37608 2839
rect 37556 2796 37608 2805
rect 38292 2796 38344 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 12256 2592 12308 2644
rect 13912 2592 13964 2644
rect 20 2524 72 2576
rect 2412 2388 2464 2440
rect 8668 2524 8720 2576
rect 12992 2524 13044 2576
rect 13636 2524 13688 2576
rect 4620 2456 4672 2508
rect 9220 2456 9272 2508
rect 17776 2592 17828 2644
rect 19340 2592 19392 2644
rect 19432 2592 19484 2644
rect 28540 2592 28592 2644
rect 28632 2592 28684 2644
rect 16856 2524 16908 2576
rect 23388 2524 23440 2576
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 7564 2388 7616 2440
rect 9680 2388 9732 2440
rect 12440 2388 12492 2440
rect 14832 2388 14884 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 8392 2252 8444 2304
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 18880 2456 18932 2508
rect 21456 2499 21508 2508
rect 21456 2465 21465 2499
rect 21465 2465 21499 2499
rect 21499 2465 21508 2499
rect 21456 2456 21508 2465
rect 24676 2499 24728 2508
rect 24676 2465 24685 2499
rect 24685 2465 24719 2499
rect 24719 2465 24728 2499
rect 24676 2456 24728 2465
rect 25964 2524 26016 2576
rect 26884 2524 26936 2576
rect 28908 2456 28960 2508
rect 11612 2252 11664 2304
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 13544 2252 13596 2304
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 18512 2388 18564 2440
rect 27068 2388 27120 2440
rect 33416 2592 33468 2644
rect 33692 2592 33744 2644
rect 34428 2592 34480 2644
rect 37556 2592 37608 2644
rect 38200 2635 38252 2644
rect 38200 2601 38209 2635
rect 38209 2601 38243 2635
rect 38243 2601 38252 2635
rect 38200 2592 38252 2601
rect 32680 2524 32732 2576
rect 32128 2456 32180 2508
rect 34244 2524 34296 2576
rect 37096 2524 37148 2576
rect 16396 2320 16448 2372
rect 16764 2252 16816 2304
rect 18696 2252 18748 2304
rect 20168 2320 20220 2372
rect 21180 2363 21232 2372
rect 21180 2329 21189 2363
rect 21189 2329 21223 2363
rect 21223 2329 21232 2363
rect 21180 2320 21232 2329
rect 21272 2320 21324 2372
rect 22744 2320 22796 2372
rect 24952 2363 25004 2372
rect 24952 2329 24961 2363
rect 24961 2329 24995 2363
rect 24995 2329 25004 2363
rect 24952 2320 25004 2329
rect 21916 2252 21968 2304
rect 22468 2252 22520 2304
rect 25964 2252 26016 2304
rect 27620 2252 27672 2304
rect 31116 2320 31168 2372
rect 29276 2252 29328 2304
rect 30288 2252 30340 2304
rect 31392 2252 31444 2304
rect 32772 2320 32824 2372
rect 34336 2388 34388 2440
rect 35440 2388 35492 2440
rect 35716 2388 35768 2440
rect 37464 2431 37516 2440
rect 34428 2320 34480 2372
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 35716 2295 35768 2304
rect 35716 2261 35725 2295
rect 35725 2261 35759 2295
rect 35759 2261 35768 2295
rect 35716 2252 35768 2261
rect 37188 2252 37240 2304
rect 37372 2252 37424 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 15292 2048 15344 2100
rect 24860 2048 24912 2100
rect 25872 2048 25924 2100
rect 35716 2048 35768 2100
rect 16120 1980 16172 2032
rect 19432 1980 19484 2032
rect 27620 1980 27672 2032
rect 30932 1980 30984 2032
rect 16212 1912 16264 1964
rect 21180 1912 21232 1964
rect 13084 1844 13136 1896
rect 21088 1844 21140 1896
rect 28540 1912 28592 1964
rect 38016 1912 38068 1964
rect 23204 1844 23256 1896
<< metal2 >>
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 2962 39536 3018 39545
rect 2962 39471 3018 39480
rect 1320 37126 1348 39200
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 2608 37210 2636 39200
rect 2870 37496 2926 37505
rect 2870 37431 2926 37440
rect 1308 37120 1360 37126
rect 1308 37062 1360 37068
rect 1674 36136 1730 36145
rect 1674 36071 1730 36080
rect 1688 36038 1716 36071
rect 1676 36032 1728 36038
rect 1676 35974 1728 35980
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 1688 34105 1716 34342
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1596 32065 1624 32370
rect 1582 32056 1638 32065
rect 1582 31991 1584 32000
rect 1636 31991 1638 32000
rect 1584 31962 1636 31968
rect 1674 30696 1730 30705
rect 1674 30631 1676 30640
rect 1728 30631 1730 30640
rect 1676 30602 1728 30608
rect 1688 30394 1716 30602
rect 1676 30388 1728 30394
rect 1676 30330 1728 30336
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1596 28694 1624 29106
rect 1584 28688 1636 28694
rect 1582 28656 1584 28665
rect 1636 28656 1638 28665
rect 1582 28591 1638 28600
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26625 1716 26726
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1780 26042 1808 37198
rect 2608 37182 2820 37210
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2884 36854 2912 37431
rect 2872 36848 2924 36854
rect 2872 36790 2924 36796
rect 2044 36644 2096 36650
rect 2044 36586 2096 36592
rect 1860 36168 1912 36174
rect 1860 36110 1912 36116
rect 1872 34746 1900 36110
rect 1860 34740 1912 34746
rect 1860 34682 1912 34688
rect 1860 30660 1912 30666
rect 1860 30602 1912 30608
rect 1768 26036 1820 26042
rect 1768 25978 1820 25984
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1596 24954 1624 25191
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23225 1716 23462
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21185 1716 21286
rect 1674 21176 1730 21185
rect 1780 21146 1808 21490
rect 1674 21111 1730 21120
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1872 20262 1900 30602
rect 2056 26926 2084 36586
rect 2884 36378 2912 36790
rect 2976 36786 3004 39471
rect 4526 39200 4582 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28354 39200 28410 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4068 37256 4120 37262
rect 4068 37198 4120 37204
rect 2964 36780 3016 36786
rect 2964 36722 3016 36728
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 2136 34604 2188 34610
rect 2136 34546 2188 34552
rect 2148 33862 2176 34546
rect 2136 33856 2188 33862
rect 2136 33798 2188 33804
rect 2044 26920 2096 26926
rect 2044 26862 2096 26868
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1964 20942 1992 25230
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1688 19718 1716 19751
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1964 18290 1992 20878
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1596 17814 1624 18226
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1674 14376 1730 14385
rect 1674 14311 1730 14320
rect 1688 14278 1716 14311
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10305 1624 10610
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1582 10296 1638 10305
rect 1780 10266 1808 10406
rect 1582 10231 1584 10240
rect 1636 10231 1638 10240
rect 1768 10260 1820 10266
rect 1584 10202 1636 10208
rect 1768 10202 1820 10208
rect 1584 8968 1636 8974
rect 1582 8936 1584 8945
rect 1636 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8634 1624 8871
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2056 8294 2084 25842
rect 2148 16182 2176 33798
rect 4080 30122 4108 37198
rect 4632 37126 4660 37726
rect 6472 37126 6500 39200
rect 7760 37262 7788 39200
rect 9692 37262 9720 39200
rect 7288 37256 7340 37262
rect 7288 37198 7340 37204
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 5448 37120 5500 37126
rect 5448 37062 5500 37068
rect 6460 37120 6512 37126
rect 6460 37062 6512 37068
rect 5460 36922 5488 37062
rect 5448 36916 5500 36922
rect 5448 36858 5500 36864
rect 7300 36582 7328 37198
rect 11624 37126 11652 39200
rect 11980 37256 12032 37262
rect 11980 37198 12032 37204
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 9956 37120 10008 37126
rect 9956 37062 10008 37068
rect 11612 37120 11664 37126
rect 11612 37062 11664 37068
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30116 4120 30122
rect 4068 30058 4120 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2884 16454 2912 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 6840 21146 6868 26930
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4724 18970 4752 19790
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 8036 18630 8064 37062
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 2136 16176 2188 16182
rect 2136 16118 2188 16124
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15502 4660 16390
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 9042 4108 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2056 7478 2084 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4865 1716 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 1674 4856 1730 4865
rect 4214 4859 4522 4868
rect 1674 4791 1730 4800
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1584 3528 1636 3534
rect 1582 3496 1584 3505
rect 1636 3496 1638 3505
rect 1582 3431 1638 3440
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1780 3398 1808 3431
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 2424 2446 2452 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2514 4660 15438
rect 8956 11354 8984 20742
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9232 9722 9260 10610
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 6840 8294 6868 9658
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 7576 2446 7604 2790
rect 8680 2582 8708 9318
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 9232 2514 9260 5510
rect 9968 4146 9996 37062
rect 11992 24138 12020 37198
rect 12912 37126 12940 39200
rect 14556 37392 14608 37398
rect 14556 37334 14608 37340
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 13280 36582 13308 37198
rect 13268 36576 13320 36582
rect 13268 36518 13320 36524
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 12452 29102 12480 29990
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 13280 21418 13308 36518
rect 14568 26234 14596 37334
rect 14844 37330 14872 39200
rect 16776 37482 16804 39200
rect 16684 37454 16804 37482
rect 18064 37466 18092 39200
rect 18052 37460 18104 37466
rect 16684 37330 16712 37454
rect 18052 37402 18104 37408
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 16672 37324 16724 37330
rect 16672 37266 16724 37272
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 15212 36786 15240 37198
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 14476 26206 14596 26234
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 14476 20806 14504 26206
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 16658 12940 18566
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10520 15706 10548 15982
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10612 13530 10640 16050
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13174 13832 13230 13841
rect 13174 13767 13176 13776
rect 13228 13767 13230 13776
rect 13176 13738 13228 13744
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 13372 13190 13400 13942
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10980 10266 11008 12786
rect 12898 12472 12954 12481
rect 13096 12442 13124 12922
rect 13372 12850 13400 13126
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 12898 12407 12954 12416
rect 13084 12436 13136 12442
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11992 9654 12020 11766
rect 12912 11150 12940 12407
rect 13084 12378 13136 12384
rect 13464 11762 13492 20742
rect 15856 18426 15884 33254
rect 15948 28082 15976 36722
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13648 14006 13676 15030
rect 14660 15026 14688 16594
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12452 7886 12480 8910
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12452 7410 12480 7822
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10336 4826 10364 5170
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10428 4457 10456 4558
rect 10414 4448 10470 4457
rect 10414 4383 10470 4392
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10060 2650 10088 3130
rect 12268 2650 12296 6734
rect 12452 5234 12480 7346
rect 12544 6458 12572 10202
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12452 3534 12480 5170
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12728 2922 12756 10950
rect 12912 10810 12940 11086
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6934 12848 7142
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5953 13216 6258
rect 13174 5944 13230 5953
rect 13280 5914 13308 10746
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13372 8634 13400 10134
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6322 13400 6734
rect 13464 6458 13492 7686
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13174 5879 13230 5888
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 12452 2446 12480 2790
rect 13004 2582 13032 3130
rect 13556 2774 13584 11086
rect 13648 10674 13676 12582
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11898 13768 12106
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13924 9586 13952 14758
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14200 13938 14228 14554
rect 14844 14414 14872 15302
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14280 14000 14332 14006
rect 14278 13968 14280 13977
rect 14332 13968 14334 13977
rect 14188 13932 14240 13938
rect 14108 13892 14188 13920
rect 14108 12238 14136 13892
rect 14278 13903 14334 13912
rect 14188 13874 14240 13880
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14200 12850 14228 13670
rect 14384 13394 14412 14214
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14752 13462 14780 13738
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14384 12782 14412 13194
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14200 11286 14228 12650
rect 14384 12434 14412 12718
rect 14292 12406 14412 12434
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14292 11150 14320 12406
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14476 11150 14504 11698
rect 14660 11694 14688 12174
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14292 10742 14320 11086
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13648 8362 13676 9522
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9178 13768 9318
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13818 8936 13874 8945
rect 13818 8871 13874 8880
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13634 8120 13690 8129
rect 13634 8055 13690 8064
rect 13648 6730 13676 8055
rect 13832 7562 13860 8871
rect 13924 8566 13952 9522
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 8906 14044 9386
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13910 8256 13966 8265
rect 13910 8191 13966 8200
rect 13740 7534 13860 7562
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13740 5914 13768 7534
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7041 13860 7346
rect 13818 7032 13874 7041
rect 13818 6967 13874 6976
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13636 5704 13688 5710
rect 13832 5692 13860 6734
rect 13924 6458 13952 8191
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13688 5664 13860 5692
rect 13636 5646 13688 5652
rect 13648 4622 13676 5646
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13924 2854 13952 3946
rect 14016 2990 14044 8842
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 5370 14136 8298
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 6798 14228 7346
rect 14292 7002 14320 8463
rect 14568 7818 14596 9998
rect 14660 8498 14688 11630
rect 14844 10062 14872 14350
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 12306 15056 13806
rect 15304 13326 15332 17002
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15396 14550 15424 15574
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12646 15332 13262
rect 15396 13190 15424 14214
rect 15488 13938 15516 18226
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15764 16182 15792 16390
rect 15752 16176 15804 16182
rect 15804 16136 15884 16164
rect 15752 16118 15804 16124
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15566 14104 15622 14113
rect 15566 14039 15568 14048
rect 15620 14039 15622 14048
rect 15568 14010 15620 14016
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15488 12850 15516 13466
rect 15764 13258 15792 14826
rect 15856 14414 15884 16136
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 16132 13394 16160 27814
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15502 16436 15846
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16500 14958 16528 18090
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16578 15056 16634 15065
rect 16684 15026 16712 15302
rect 16578 14991 16580 15000
rect 16632 14991 16634 15000
rect 16672 15020 16724 15026
rect 16580 14962 16632 14968
rect 16672 14962 16724 14968
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16304 13864 16356 13870
rect 16302 13832 16304 13841
rect 16356 13832 16358 13841
rect 16302 13767 16358 13776
rect 16394 13424 16450 13433
rect 16120 13388 16172 13394
rect 16394 13359 16450 13368
rect 16120 13330 16172 13336
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 16408 12850 16436 13359
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15488 12170 15516 12650
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 10674 15148 11494
rect 15396 11218 15424 12106
rect 15580 11370 15608 12786
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15488 11342 15608 11370
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15488 11150 15516 11342
rect 15566 11248 15622 11257
rect 15566 11183 15622 11192
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 10742 15424 11018
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14752 9722 14780 9998
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7546 14688 7686
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14108 4486 14136 5306
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 4049 14136 4082
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14108 3738 14136 3975
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14292 3126 14320 6054
rect 14476 5710 14504 6258
rect 14752 5846 14780 9658
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14844 7177 14872 8366
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 7886 15056 8230
rect 15212 7954 15240 10406
rect 15580 10266 15608 11183
rect 15672 10606 15700 11630
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15382 10160 15438 10169
rect 15382 10095 15384 10104
rect 15436 10095 15438 10104
rect 15384 10066 15436 10072
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15382 9616 15438 9625
rect 15382 9551 15438 9560
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 8634 15332 8910
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15304 7993 15332 8570
rect 15290 7984 15346 7993
rect 15200 7948 15252 7954
rect 15290 7919 15346 7928
rect 15200 7890 15252 7896
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15304 7478 15332 7822
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14830 7168 14886 7177
rect 14830 7103 14886 7112
rect 15028 7002 15056 7346
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15396 6798 15424 9551
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15396 5914 15424 6190
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 15198 5808 15254 5817
rect 15198 5743 15254 5752
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14476 5234 14504 5646
rect 14924 5568 14976 5574
rect 14922 5536 14924 5545
rect 14976 5536 14978 5545
rect 14922 5471 14978 5480
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 15212 5166 15240 5743
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 4214 14688 4422
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14476 3534 14504 4082
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14476 3126 14504 3470
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13556 2746 13676 2774
rect 13648 2582 13676 2746
rect 13924 2650 13952 2790
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 15212 2446 15240 2926
rect 15488 2854 15516 9998
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15580 5914 15608 8842
rect 15672 6866 15700 9454
rect 15764 9217 15792 9862
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15750 9208 15806 9217
rect 15750 9143 15806 9152
rect 15856 8634 15884 9590
rect 15948 9518 15976 12582
rect 16500 12442 16528 12582
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16316 11937 16344 12106
rect 16302 11928 16358 11937
rect 16302 11863 16358 11872
rect 16316 11830 16344 11863
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16592 11626 16620 13874
rect 16684 12170 16712 14758
rect 16776 13870 16804 37266
rect 18064 37262 18092 37402
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 19996 37126 20024 39200
rect 21928 37330 21956 39200
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 17500 36644 17552 36650
rect 17500 36586 17552 36592
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17420 16590 17448 17206
rect 17512 16794 17540 36586
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 18144 34536 18196 34542
rect 18144 34478 18196 34484
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16854 14104 16910 14113
rect 16854 14039 16910 14048
rect 16868 13938 16896 14039
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16854 13560 16910 13569
rect 16854 13495 16856 13504
rect 16908 13495 16910 13504
rect 16856 13466 16908 13472
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16776 11218 16804 12718
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16868 11082 16896 12310
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15948 9042 15976 9454
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 16040 7410 16068 10542
rect 16224 10470 16252 10950
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16210 10024 16266 10033
rect 16210 9959 16266 9968
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16132 7206 16160 7754
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16224 6866 16252 9959
rect 16408 7954 16436 11018
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16592 10674 16620 10746
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16578 10568 16634 10577
rect 16578 10503 16634 10512
rect 16672 10532 16724 10538
rect 16592 8922 16620 10503
rect 16672 10474 16724 10480
rect 16684 9994 16712 10474
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16776 9058 16804 9930
rect 16500 8906 16620 8922
rect 16488 8900 16620 8906
rect 16540 8894 16620 8900
rect 16684 9030 16804 9058
rect 16488 8842 16540 8848
rect 16580 8832 16632 8838
rect 16578 8800 16580 8809
rect 16632 8800 16634 8809
rect 16578 8735 16634 8744
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16408 7546 16436 7754
rect 16592 7546 16620 7958
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16684 7478 16712 9030
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15764 5370 15792 6326
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 16040 5914 16068 6122
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15948 4690 15976 5782
rect 16132 5710 16160 6734
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16210 5672 16266 5681
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 5137 16068 5170
rect 16026 5128 16082 5137
rect 16026 5063 16082 5072
rect 16132 4865 16160 5646
rect 16210 5607 16212 5616
rect 16264 5607 16266 5616
rect 16212 5578 16264 5584
rect 16118 4856 16174 4865
rect 16118 4791 16174 4800
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15672 4214 15700 4558
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15764 3233 15792 4626
rect 15934 4584 15990 4593
rect 15934 4519 15990 4528
rect 15948 3670 15976 4519
rect 16316 4457 16344 6258
rect 16302 4448 16358 4457
rect 16302 4383 16358 4392
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15750 3224 15806 3233
rect 15750 3159 15806 3168
rect 16316 2990 16344 4082
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 16132 2446 16160 2858
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 9692 800 9720 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 11624 800 11652 2246
rect 13096 1902 13124 2246
rect 13084 1896 13136 1902
rect 13084 1838 13136 1844
rect 13556 800 13584 2246
rect 14844 800 14872 2382
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 2106 15332 2246
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 16132 2038 16160 2382
rect 16120 2032 16172 2038
rect 16120 1974 16172 1980
rect 16224 1970 16252 2790
rect 16408 2378 16436 7346
rect 16578 7304 16634 7313
rect 16578 7239 16634 7248
rect 16672 7268 16724 7274
rect 16592 6458 16620 7239
rect 16672 7210 16724 7216
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16684 6254 16712 7210
rect 16868 6866 16896 8842
rect 16960 7478 16988 15914
rect 17144 15706 17172 16118
rect 17696 15978 17724 18294
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16561 17908 17070
rect 17866 16552 17922 16561
rect 17866 16487 17922 16496
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17236 15502 17264 15846
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17328 15042 17356 15574
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17236 15014 17356 15042
rect 17236 14414 17264 15014
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17038 13968 17094 13977
rect 17038 13903 17040 13912
rect 17092 13903 17094 13912
rect 17040 13874 17092 13880
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12714 17172 13262
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17038 12200 17094 12209
rect 17038 12135 17094 12144
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 17052 7274 17080 12135
rect 17144 11014 17172 12650
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17236 10198 17264 13398
rect 17328 12345 17356 14894
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17420 14074 17448 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17590 13696 17646 13705
rect 17590 13631 17646 13640
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17420 12442 17448 12786
rect 17408 12436 17460 12442
rect 17604 12434 17632 13631
rect 17696 12617 17724 15506
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17408 12378 17460 12384
rect 17512 12406 17632 12434
rect 17314 12336 17370 12345
rect 17314 12271 17370 12280
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 11286 17356 12106
rect 17408 11824 17460 11830
rect 17406 11792 17408 11801
rect 17460 11792 17462 11801
rect 17406 11727 17462 11736
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17144 9382 17172 9454
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17236 9058 17264 10134
rect 17314 9208 17370 9217
rect 17314 9143 17370 9152
rect 17144 9042 17264 9058
rect 17132 9036 17264 9042
rect 17184 9030 17264 9036
rect 17132 8978 17184 8984
rect 17328 8838 17356 9143
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17222 8664 17278 8673
rect 17222 8599 17224 8608
rect 17276 8599 17278 8608
rect 17224 8570 17276 8576
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 8362 17172 8434
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17420 7857 17448 11630
rect 17406 7848 17462 7857
rect 17406 7783 17462 7792
rect 17132 7472 17184 7478
rect 17132 7414 17184 7420
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17038 6760 17094 6769
rect 16960 6458 16988 6734
rect 17038 6695 17040 6704
rect 17092 6695 17094 6704
rect 17040 6666 17092 6672
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16592 5001 16620 5578
rect 16578 4992 16634 5001
rect 16578 4927 16634 4936
rect 16592 4486 16620 4927
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16500 3602 16528 4150
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16684 3466 16712 5782
rect 16946 5400 17002 5409
rect 16946 5335 16948 5344
rect 17000 5335 17002 5344
rect 16948 5306 17000 5312
rect 17144 5302 17172 7414
rect 17222 6896 17278 6905
rect 17222 6831 17278 6840
rect 17236 6798 17264 6831
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16854 4720 16910 4729
rect 16854 4655 16856 4664
rect 16908 4655 16910 4664
rect 16856 4626 16908 4632
rect 17052 4282 17080 5170
rect 17512 4758 17540 12406
rect 17696 11370 17724 12543
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17604 11342 17724 11370
rect 17788 11354 17816 11766
rect 17776 11348 17828 11354
rect 17604 8566 17632 11342
rect 17776 11290 17828 11296
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17696 9654 17724 11154
rect 17774 10704 17830 10713
rect 17774 10639 17776 10648
rect 17828 10639 17830 10648
rect 17776 10610 17828 10616
rect 17880 10538 17908 16487
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 15706 18092 16390
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 18064 15502 18092 15642
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18156 14482 18184 34478
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20088 22778 20116 26930
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 17270 18552 17478
rect 18708 17338 18736 19382
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18984 18426 19012 18702
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19352 18222 19380 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19378 20024 20198
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 18340 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19524 18352 19576 18358
rect 19444 18312 19524 18340
rect 19524 18294 19576 18300
rect 19720 18222 19748 18362
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19996 18154 20024 19314
rect 20272 18834 20300 19654
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19168 17678 19196 17750
rect 19996 17678 20024 18090
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18432 16046 18460 17070
rect 18708 16590 18736 17274
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 19168 15994 19196 17614
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16114 19288 16526
rect 19352 16522 19380 17070
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 18604 15972 18656 15978
rect 19168 15966 19288 15994
rect 18604 15914 18656 15920
rect 18616 15858 18644 15914
rect 18432 15830 18644 15858
rect 18326 15056 18382 15065
rect 18326 14991 18382 15000
rect 18340 14958 18368 14991
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17972 13530 18000 14214
rect 18156 14006 18184 14418
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18340 13870 18368 14282
rect 18144 13864 18196 13870
rect 18328 13864 18380 13870
rect 18144 13806 18196 13812
rect 18248 13824 18328 13852
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18064 13394 18092 13738
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 17972 11694 18000 12854
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18064 11354 18092 13194
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18156 11234 18184 13806
rect 18248 12306 18276 13824
rect 18328 13806 18380 13812
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18064 11206 18184 11234
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17958 10160 18014 10169
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17696 8430 17724 9590
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17788 7954 17816 10134
rect 17958 10095 18014 10104
rect 17972 9994 18000 10095
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17880 9518 17908 9930
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17880 9110 17908 9454
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17972 9110 18000 9386
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17868 8560 17920 8566
rect 17920 8508 18000 8514
rect 17868 8502 18000 8508
rect 17880 8486 18000 8502
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 5846 17632 7346
rect 17788 7274 17816 7890
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17696 5846 17724 6190
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17604 4758 17632 5782
rect 17684 5092 17736 5098
rect 17684 5034 17736 5040
rect 17500 4752 17552 4758
rect 17314 4720 17370 4729
rect 17500 4694 17552 4700
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17314 4655 17316 4664
rect 17368 4655 17370 4664
rect 17316 4626 17368 4632
rect 17224 4480 17276 4486
rect 17316 4480 17368 4486
rect 17224 4422 17276 4428
rect 17314 4448 17316 4457
rect 17368 4448 17370 4457
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17236 3738 17264 4422
rect 17314 4383 17370 4392
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16868 2582 16896 3470
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17144 3126 17172 3334
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17512 2922 17540 4694
rect 17696 3738 17724 5034
rect 17788 4486 17816 7210
rect 17972 6866 18000 8486
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18064 6798 18092 11206
rect 18340 11150 18368 12378
rect 18328 11144 18380 11150
rect 18326 11112 18328 11121
rect 18380 11112 18382 11121
rect 18326 11047 18382 11056
rect 18144 10600 18196 10606
rect 18328 10600 18380 10606
rect 18144 10542 18196 10548
rect 18248 10560 18328 10588
rect 18156 9994 18184 10542
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18248 9382 18276 10560
rect 18328 10542 18380 10548
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18340 9654 18368 9862
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8906 18276 9318
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18156 7750 18184 8026
rect 18144 7744 18196 7750
rect 18248 7732 18276 8842
rect 18340 8673 18368 8842
rect 18326 8664 18382 8673
rect 18326 8599 18382 8608
rect 18432 7954 18460 15830
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 18524 15094 18552 15302
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18510 13832 18566 13841
rect 18510 13767 18566 13776
rect 18524 13190 18552 13767
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 10130 18552 13126
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18616 11626 18644 12378
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18616 11218 18644 11562
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18524 8809 18552 10066
rect 18616 9926 18644 10950
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18708 9194 18736 14554
rect 19168 14346 19196 15302
rect 19260 14958 19288 15966
rect 19248 14952 19300 14958
rect 19352 14940 19380 16458
rect 19444 15570 19472 17546
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20272 16998 20300 17138
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19432 14952 19484 14958
rect 19352 14912 19432 14940
rect 19248 14894 19300 14900
rect 19432 14894 19484 14900
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 14006 19196 14282
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18984 12918 19012 13194
rect 18972 12912 19024 12918
rect 18800 12872 18972 12900
rect 18800 9450 18828 12872
rect 18972 12854 19024 12860
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18984 12170 19012 12310
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18892 11150 18920 11494
rect 18984 11286 19012 11630
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18616 9166 18736 9194
rect 18510 8800 18566 8809
rect 18510 8735 18566 8744
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18248 7704 18460 7732
rect 18144 7686 18196 7692
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18432 6746 18460 7704
rect 18616 6866 18644 9166
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 17880 4729 17908 6734
rect 18432 6718 18644 6746
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18144 5840 18196 5846
rect 17972 5788 18144 5794
rect 17972 5782 18196 5788
rect 17972 5778 18184 5782
rect 17960 5772 18184 5778
rect 18012 5766 18184 5772
rect 17960 5714 18012 5720
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17866 4720 17922 4729
rect 17866 4655 17922 4664
rect 17972 4554 18000 5034
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17972 4049 18000 4150
rect 17958 4040 18014 4049
rect 17958 3975 18014 3984
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17972 3534 18000 3975
rect 18064 3942 18092 5238
rect 18156 4826 18184 5306
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18248 5030 18276 5102
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18236 4140 18288 4146
rect 18340 4128 18368 6326
rect 18432 4826 18460 6326
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18288 4100 18368 4128
rect 18236 4082 18288 4088
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18156 3602 18184 4014
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18248 3126 18276 3878
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17788 2650 17816 2858
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 18524 2446 18552 6598
rect 18616 3126 18644 6718
rect 18708 5302 18736 8978
rect 18800 7954 18828 9386
rect 18892 8265 18920 9590
rect 18878 8256 18934 8265
rect 18878 8191 18934 8200
rect 18878 8120 18934 8129
rect 19076 8090 19104 13942
rect 19260 13530 19288 14894
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 13938 19380 14758
rect 19536 14618 19564 15030
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19614 14648 19670 14657
rect 19524 14612 19576 14618
rect 19996 14618 20024 14826
rect 20088 14657 20116 16526
rect 20272 15586 20300 16934
rect 20180 15558 20300 15586
rect 20074 14648 20130 14657
rect 19614 14583 19670 14592
rect 19984 14612 20036 14618
rect 19524 14554 19576 14560
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19444 13394 19472 14418
rect 19628 14414 19656 14583
rect 20074 14583 20130 14592
rect 19984 14554 20036 14560
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19154 11928 19210 11937
rect 19154 11863 19210 11872
rect 19168 11830 19196 11863
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 19246 11792 19302 11801
rect 19246 11727 19302 11736
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 18878 8055 18934 8064
rect 19064 8084 19116 8090
rect 18892 8022 18920 8055
rect 19064 8026 19116 8032
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18800 6186 18828 7754
rect 19168 7698 19196 8298
rect 19260 8294 19288 11727
rect 19444 11694 19472 13330
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19524 12912 19576 12918
rect 19522 12880 19524 12889
rect 19576 12880 19578 12889
rect 19522 12815 19578 12824
rect 19996 12434 20024 14554
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20088 12850 20116 14486
rect 20180 13462 20208 15558
rect 20364 15162 20392 37198
rect 21180 36916 21232 36922
rect 21180 36858 21232 36864
rect 21088 35080 21140 35086
rect 21088 35022 21140 35028
rect 21100 32230 21128 35022
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 20720 29572 20772 29578
rect 20720 29514 20772 29520
rect 20732 29034 20760 29514
rect 20720 29028 20772 29034
rect 20720 28970 20772 28976
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20640 27130 20668 27814
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20732 26234 20760 28970
rect 20732 26206 20852 26234
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20548 22094 20576 25094
rect 20456 22066 20576 22094
rect 20456 16726 20484 22066
rect 20824 21690 20852 26206
rect 21100 25498 21128 32166
rect 21192 28762 21220 36858
rect 22296 36854 22324 37198
rect 22572 36922 22600 37198
rect 23216 37126 23244 39200
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22284 36848 22336 36854
rect 22284 36790 22336 36796
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22204 29170 22232 29786
rect 22296 29170 22324 36790
rect 23112 36780 23164 36786
rect 23112 36722 23164 36728
rect 23124 36582 23152 36722
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 23124 36378 23152 36518
rect 23112 36372 23164 36378
rect 23112 36314 23164 36320
rect 23124 29850 23152 36314
rect 23400 35290 23428 37198
rect 25148 37126 25176 39200
rect 27080 37126 27108 39200
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23112 29844 23164 29850
rect 23112 29786 23164 29792
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 23572 29028 23624 29034
rect 23572 28970 23624 28976
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21100 25294 21128 25434
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20916 19922 20944 22374
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20548 18426 20576 19382
rect 20732 18698 20760 19654
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20824 18970 20852 19382
rect 20916 19310 20944 19858
rect 21100 19854 21128 20402
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20916 18850 20944 19110
rect 20824 18822 20944 18850
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20824 18578 20852 18822
rect 21100 18766 21128 19790
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20732 18550 20852 18578
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20456 15570 20484 16662
rect 20640 16522 20668 16934
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 14346 20300 14418
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20272 12782 20300 14282
rect 20364 14006 20392 14486
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20456 13938 20484 14214
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20548 13734 20576 15302
rect 20640 14822 20668 16050
rect 20732 15978 20760 18550
rect 20916 17882 20944 18634
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20916 17270 20944 17818
rect 21088 17672 21140 17678
rect 21086 17640 21088 17649
rect 21140 17640 21142 17649
rect 20996 17604 21048 17610
rect 21086 17575 21142 17584
rect 20996 17546 21048 17552
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 21008 15570 21036 17546
rect 21100 17202 21128 17575
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 17270 21220 17478
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20628 14816 20680 14822
rect 21100 14770 21128 16662
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 20628 14758 20680 14764
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 19996 12406 20116 12434
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19522 11384 19578 11393
rect 19340 11348 19392 11354
rect 19522 11319 19578 11328
rect 19340 11290 19392 11296
rect 19352 10452 19380 11290
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10606 19472 11154
rect 19536 11150 19564 11319
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19616 10464 19668 10470
rect 19352 10424 19472 10452
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19352 8906 19380 9930
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19352 8362 19380 8502
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19338 8120 19394 8129
rect 19338 8055 19394 8064
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19076 7670 19196 7698
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18892 5710 18920 7210
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18788 5568 18840 5574
rect 18786 5536 18788 5545
rect 18840 5536 18842 5545
rect 18786 5471 18842 5480
rect 18984 5302 19012 6734
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 18786 5128 18842 5137
rect 18786 5063 18788 5072
rect 18840 5063 18842 5072
rect 18788 5034 18840 5040
rect 18696 5024 18748 5030
rect 18694 4992 18696 5001
rect 18748 4992 18750 5001
rect 18694 4927 18750 4936
rect 18694 4856 18750 4865
rect 18694 4791 18696 4800
rect 18748 4791 18750 4800
rect 18696 4762 18748 4768
rect 18708 3466 18736 4762
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 18786 3224 18842 3233
rect 18786 3159 18842 3168
rect 18800 3126 18828 3159
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18892 3058 18920 4422
rect 18984 4146 19012 4626
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19076 2938 19104 7670
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19168 6361 19196 7482
rect 19260 7274 19288 7822
rect 19352 7585 19380 8055
rect 19338 7576 19394 7585
rect 19338 7511 19394 7520
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19154 6352 19210 6361
rect 19154 6287 19210 6296
rect 19154 5944 19210 5953
rect 19154 5879 19210 5888
rect 19168 5778 19196 5879
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 19168 5409 19196 5578
rect 19154 5400 19210 5409
rect 19154 5335 19210 5344
rect 19260 5234 19288 6802
rect 19352 6730 19380 7414
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19260 4622 19288 5170
rect 19352 5001 19380 6394
rect 19444 6254 19472 10424
rect 19616 10406 19668 10412
rect 19628 10198 19656 10406
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19628 9994 19656 10134
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9110 20024 9930
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19720 8906 19748 9046
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 8090 19656 8366
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19616 7540 19668 7546
rect 19536 7500 19616 7528
rect 19536 7342 19564 7500
rect 19616 7482 19668 7488
rect 19614 7440 19670 7449
rect 19890 7440 19946 7449
rect 19614 7375 19670 7384
rect 19800 7404 19852 7410
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19628 7206 19656 7375
rect 19890 7375 19946 7384
rect 19800 7346 19852 7352
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19812 6730 19840 7346
rect 19904 7342 19932 7375
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19800 6724 19852 6730
rect 19800 6666 19852 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 7754
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 20088 6390 20116 12406
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 8430 20208 12038
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20272 10606 20300 11834
rect 20364 11830 20392 13466
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20456 12434 20484 13398
rect 20548 13394 20576 13670
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20548 12850 20576 13330
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20456 12406 20576 12434
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20364 11286 20392 11766
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20456 10606 20484 11222
rect 20548 10962 20576 12406
rect 20640 11801 20668 14758
rect 21008 14742 21128 14770
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 13462 20944 14282
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20810 13288 20866 13297
rect 20720 13252 20772 13258
rect 20810 13223 20866 13232
rect 20720 13194 20772 13200
rect 20626 11792 20682 11801
rect 20626 11727 20682 11736
rect 20732 11626 20760 13194
rect 20824 12782 20852 13223
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 21008 12434 21036 14742
rect 21192 13802 21220 16594
rect 21284 14822 21312 24074
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21376 17746 21404 18226
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21376 16658 21404 17682
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21454 15600 21510 15609
rect 21454 15535 21456 15544
rect 21508 15535 21510 15544
rect 21456 15506 21508 15512
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 13818 21312 14214
rect 21376 13938 21404 15438
rect 21560 14414 21588 18090
rect 21744 17814 21772 19314
rect 22112 18970 22140 19722
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22204 18850 22232 28970
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23400 27674 23428 28358
rect 23388 27668 23440 27674
rect 23388 27610 23440 27616
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19446 22508 20198
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 22204 18834 22324 18850
rect 22192 18828 22324 18834
rect 22244 18822 22324 18828
rect 22192 18770 22244 18776
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22204 18426 22232 18634
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22204 17814 22232 18226
rect 21732 17808 21784 17814
rect 21732 17750 21784 17756
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 21744 16522 21772 17750
rect 21822 17640 21878 17649
rect 22296 17626 22324 18822
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22388 18222 22416 18770
rect 22664 18630 22692 19722
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22296 17610 22416 17626
rect 22296 17604 22428 17610
rect 22296 17598 22376 17604
rect 21822 17575 21878 17584
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21652 13977 21680 15642
rect 21744 15434 21772 16458
rect 21732 15428 21784 15434
rect 21732 15370 21784 15376
rect 21836 15314 21864 17575
rect 22376 17546 22428 17552
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21928 16574 21956 16934
rect 22020 16726 22048 16934
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 21928 16546 22232 16574
rect 22204 16504 22232 16546
rect 22376 16516 22428 16522
rect 22204 16476 22376 16504
rect 22376 16458 22428 16464
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21928 15434 21956 16390
rect 22480 16182 22508 18022
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22192 16040 22244 16046
rect 22112 15988 22192 15994
rect 22112 15982 22244 15988
rect 22112 15966 22232 15982
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21836 15286 21956 15314
rect 21822 14784 21878 14793
rect 21822 14719 21878 14728
rect 21836 14414 21864 14719
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21638 13968 21694 13977
rect 21364 13932 21416 13938
rect 21638 13903 21694 13912
rect 21364 13874 21416 13880
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 21180 13796 21232 13802
rect 21284 13790 21588 13818
rect 21180 13738 21232 13744
rect 21100 12866 21128 13738
rect 21192 13297 21220 13738
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21178 13288 21234 13297
rect 21178 13223 21234 13232
rect 21100 12850 21220 12866
rect 21100 12844 21232 12850
rect 21100 12838 21180 12844
rect 21180 12786 21232 12792
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 12442 21128 12582
rect 20824 12406 21036 12434
rect 21088 12436 21140 12442
rect 20824 12345 20852 12406
rect 21088 12378 21140 12384
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20824 11150 20852 12271
rect 21192 12170 21220 12650
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 21086 11112 21142 11121
rect 20996 11076 21048 11082
rect 21086 11047 21142 11056
rect 20996 11018 21048 11024
rect 20548 10934 20760 10962
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20180 7478 20208 8026
rect 20168 7472 20220 7478
rect 20272 7449 20300 10542
rect 20456 10198 20484 10542
rect 20626 10432 20682 10441
rect 20626 10367 20682 10376
rect 20534 10296 20590 10305
rect 20640 10266 20668 10367
rect 20534 10231 20590 10240
rect 20628 10260 20680 10266
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20548 9994 20576 10231
rect 20628 10202 20680 10208
rect 20732 9994 20760 10934
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 20824 10266 20852 10678
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20916 10146 20944 10474
rect 20824 10118 20944 10146
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20824 9722 20852 10118
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20916 9722 20944 9998
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 21008 9330 21036 11018
rect 20824 9302 21036 9330
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20640 8498 20668 9114
rect 20824 8634 20852 9302
rect 21100 9194 21128 11047
rect 20916 9166 21128 9194
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20168 7414 20220 7420
rect 20258 7440 20314 7449
rect 20258 7375 20314 7384
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 20180 6089 20208 7278
rect 20364 7206 20392 8434
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20352 7200 20404 7206
rect 20272 7160 20352 7188
rect 20272 6225 20300 7160
rect 20352 7142 20404 7148
rect 20640 6914 20668 8230
rect 20732 8090 20760 8502
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20916 7750 20944 9166
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21008 8906 21036 9046
rect 21192 9042 21220 11630
rect 21284 10742 21312 13330
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11694 21404 12038
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21364 11552 21416 11558
rect 21362 11520 21364 11529
rect 21416 11520 21418 11529
rect 21362 11455 21418 11464
rect 21468 10742 21496 12786
rect 21560 12442 21588 13790
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21652 12322 21680 13398
rect 21836 12617 21864 14350
rect 21822 12608 21878 12617
rect 21822 12543 21878 12552
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21560 12306 21680 12322
rect 21548 12300 21680 12306
rect 21600 12294 21680 12300
rect 21548 12242 21600 12248
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11898 21588 12106
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21376 10441 21404 10610
rect 21362 10432 21418 10441
rect 21362 10367 21418 10376
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21100 8566 21128 8774
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20824 7562 20852 7686
rect 20824 7534 21036 7562
rect 20720 6928 20772 6934
rect 20640 6886 20720 6914
rect 20720 6870 20772 6876
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20258 6216 20314 6225
rect 20258 6151 20314 6160
rect 20166 6080 20222 6089
rect 20166 6015 20222 6024
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4010 19472 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4282 20024 5034
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19628 3738 19656 4082
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 18984 2910 19104 2938
rect 18984 2774 19012 2910
rect 18892 2746 19012 2774
rect 18892 2514 18920 2746
rect 19352 2650 19380 3402
rect 19444 2854 19472 3674
rect 19904 3398 19932 3674
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2848 19484 2854
rect 19430 2816 19432 2825
rect 19484 2816 19486 2825
rect 19430 2751 19486 2760
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 16212 1964 16264 1970
rect 16212 1906 16264 1912
rect 16776 800 16804 2246
rect 18708 800 18736 2246
rect 19444 2038 19472 2586
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19432 2032 19484 2038
rect 19432 1974 19484 1980
rect 19996 800 20024 3334
rect 20180 2378 20208 5850
rect 20272 4690 20300 6151
rect 20364 5914 20392 6258
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20456 5574 20484 6258
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20444 5160 20496 5166
rect 20548 5148 20576 5510
rect 20496 5120 20576 5148
rect 20444 5102 20496 5108
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20640 3890 20668 5782
rect 20732 4622 20760 6598
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20824 5846 20852 6190
rect 20916 6118 20944 6802
rect 21008 6662 21036 7534
rect 21100 7206 21128 8502
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21192 7274 21220 7822
rect 21284 7410 21312 9930
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 9042 21404 9318
rect 21560 9058 21588 11494
rect 21640 10736 21692 10742
rect 21640 10678 21692 10684
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 21468 9030 21588 9058
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21376 7206 21404 8978
rect 21468 8430 21496 9030
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21468 7954 21496 8230
rect 21560 8129 21588 8842
rect 21652 8634 21680 10678
rect 21744 9586 21772 12378
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21744 8566 21772 9522
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21546 8120 21602 8129
rect 21546 8055 21602 8064
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21454 7848 21510 7857
rect 21454 7783 21510 7792
rect 21468 7410 21496 7783
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20916 5642 20944 6054
rect 20996 5840 21048 5846
rect 20996 5782 21048 5788
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20812 5296 20864 5302
rect 20810 5264 20812 5273
rect 20904 5296 20956 5302
rect 20864 5264 20866 5273
rect 20904 5238 20956 5244
rect 20810 5199 20866 5208
rect 20916 4758 20944 5238
rect 20904 4752 20956 4758
rect 20904 4694 20956 4700
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20904 3936 20956 3942
rect 20640 3884 20904 3890
rect 20640 3878 20956 3884
rect 20548 3754 20576 3878
rect 20640 3862 20944 3878
rect 21008 3754 21036 5782
rect 20548 3726 21036 3754
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21008 3233 21036 3538
rect 20994 3224 21050 3233
rect 20994 3159 21050 3168
rect 21100 2530 21128 7142
rect 21376 6866 21404 7142
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21652 6730 21680 7686
rect 21744 6905 21772 8366
rect 21836 7732 21864 12543
rect 21928 8430 21956 15286
rect 22112 15162 22140 15966
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22572 15858 22600 18566
rect 22664 16726 22692 18566
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22756 17814 22784 18158
rect 22744 17808 22796 17814
rect 22744 17750 22796 17756
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22664 15978 22692 16662
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22204 15638 22232 15846
rect 22572 15830 22692 15858
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 22466 15600 22522 15609
rect 22466 15535 22522 15544
rect 22284 15360 22336 15366
rect 22336 15308 22416 15314
rect 22284 15302 22416 15308
rect 22296 15286 22416 15302
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22008 14272 22060 14278
rect 22060 14220 22324 14226
rect 22008 14214 22324 14220
rect 22020 14198 22324 14214
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 22020 13433 22048 13466
rect 22006 13424 22062 13433
rect 22006 13359 22062 13368
rect 22112 13258 22140 14010
rect 22204 13841 22232 14010
rect 22190 13832 22246 13841
rect 22190 13767 22246 13776
rect 22296 13512 22324 14198
rect 22388 14113 22416 15286
rect 22374 14104 22430 14113
rect 22374 14039 22430 14048
rect 22204 13484 22324 13512
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22204 12782 22232 13484
rect 22480 13376 22508 15535
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22296 13348 22508 13376
rect 22296 13258 22324 13348
rect 22572 13274 22600 13466
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22388 13246 22600 13274
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22020 11286 22048 12242
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22112 11121 22140 11766
rect 22190 11248 22246 11257
rect 22190 11183 22246 11192
rect 22098 11112 22154 11121
rect 22204 11082 22232 11183
rect 22098 11047 22154 11056
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22100 11008 22152 11014
rect 22098 10976 22100 10985
rect 22152 10976 22154 10985
rect 22098 10911 22154 10920
rect 22098 10840 22154 10849
rect 22098 10775 22100 10784
rect 22152 10775 22154 10784
rect 22100 10746 22152 10752
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22296 10554 22324 12854
rect 22388 12434 22416 13246
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22572 12986 22600 13126
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22388 12406 22508 12434
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21928 8090 21956 8366
rect 22020 8090 22048 9998
rect 22112 9466 22140 10542
rect 22296 10526 22416 10554
rect 22388 9738 22416 10526
rect 22480 10470 22508 12406
rect 22560 11280 22612 11286
rect 22664 11268 22692 15830
rect 22756 13394 22784 16730
rect 22848 15609 22876 21286
rect 23400 20602 23428 27610
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23204 20392 23256 20398
rect 23204 20334 23256 20340
rect 23216 19718 23244 20334
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23216 18154 23244 19654
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23204 18148 23256 18154
rect 23204 18090 23256 18096
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 22834 15600 22890 15609
rect 22834 15535 22890 15544
rect 22848 15434 22876 15535
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 23032 14482 23060 15982
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22926 14104 22982 14113
rect 22926 14039 22982 14048
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22756 12374 22784 12718
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 22848 12102 22876 13194
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22612 11240 22692 11268
rect 22560 11222 22612 11228
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22296 9710 22416 9738
rect 22466 9752 22522 9761
rect 22296 9654 22324 9710
rect 22466 9687 22468 9696
rect 22520 9687 22522 9696
rect 22468 9658 22520 9664
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22388 9466 22416 9590
rect 22112 9438 22416 9466
rect 22098 9208 22154 9217
rect 22098 9143 22100 9152
rect 22152 9143 22154 9152
rect 22100 9114 22152 9120
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21836 7721 22140 7732
rect 21836 7712 22154 7721
rect 21836 7704 22098 7712
rect 22098 7647 22154 7656
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22006 7168 22062 7177
rect 22006 7103 22062 7112
rect 22020 6914 22048 7103
rect 22112 6914 22140 7278
rect 21730 6896 21786 6905
rect 21730 6831 21786 6840
rect 21928 6886 22140 6914
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21560 6633 21588 6666
rect 21546 6624 21602 6633
rect 21546 6559 21602 6568
rect 21364 5840 21416 5846
rect 21416 5788 21588 5794
rect 21364 5782 21588 5788
rect 21376 5766 21588 5782
rect 21560 5642 21588 5766
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21192 5137 21220 5170
rect 21178 5128 21234 5137
rect 21178 5063 21234 5072
rect 21192 5030 21220 5063
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21284 4690 21312 5578
rect 21362 5400 21418 5409
rect 21362 5335 21418 5344
rect 21376 5234 21404 5335
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 21652 4758 21680 6666
rect 21744 6118 21772 6831
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21928 5642 21956 6886
rect 22204 6746 22232 8502
rect 22284 8492 22336 8498
rect 22336 8452 22416 8480
rect 22284 8434 22336 8440
rect 22112 6718 22232 6746
rect 22112 6390 22140 6718
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22100 6384 22152 6390
rect 22296 6361 22324 6394
rect 22100 6326 22152 6332
rect 22282 6352 22338 6361
rect 22282 6287 22338 6296
rect 22388 5642 22416 8452
rect 22480 7834 22508 9658
rect 22572 9450 22600 11222
rect 22650 11112 22706 11121
rect 22650 11047 22706 11056
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22664 9178 22692 11047
rect 22756 10577 22784 11766
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22742 10568 22798 10577
rect 22742 10503 22798 10512
rect 22848 10470 22876 10950
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22940 9674 22968 14039
rect 23032 13705 23060 14418
rect 23018 13696 23074 13705
rect 23018 13631 23074 13640
rect 23216 13512 23244 18090
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23308 17338 23336 17818
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23400 16522 23428 18566
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23492 15434 23520 17274
rect 23584 17134 23612 28970
rect 23768 19446 23796 29038
rect 26700 25152 26752 25158
rect 26700 25094 26752 25100
rect 25136 21412 25188 21418
rect 25136 21354 25188 21360
rect 25044 20324 25096 20330
rect 25044 20266 25096 20272
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23676 18154 23704 18702
rect 23768 18698 23796 19382
rect 24032 18896 24084 18902
rect 24032 18838 24084 18844
rect 23756 18692 23808 18698
rect 23756 18634 23808 18640
rect 23768 18358 23796 18634
rect 23756 18352 23808 18358
rect 23756 18294 23808 18300
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 23676 17678 23704 18090
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23768 17270 23796 18022
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23676 16046 23704 16594
rect 23848 16176 23900 16182
rect 23846 16144 23848 16153
rect 23900 16144 23902 16153
rect 23846 16079 23902 16088
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23032 13484 23244 13512
rect 23032 11665 23060 13484
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23018 11656 23074 11665
rect 23018 11591 23074 11600
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 10588 23060 11494
rect 23124 11098 23152 13330
rect 23308 12306 23336 14282
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 14006 23428 14214
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23400 13462 23428 13738
rect 23478 13560 23534 13569
rect 23478 13495 23534 13504
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23492 12646 23520 13495
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23584 12238 23612 15302
rect 23676 14958 23704 15982
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23860 14346 23888 14554
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23754 13968 23810 13977
rect 23754 13903 23810 13912
rect 23664 13796 23716 13802
rect 23664 13738 23716 13744
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23124 11082 23336 11098
rect 23124 11076 23348 11082
rect 23124 11070 23296 11076
rect 23296 11018 23348 11024
rect 23204 10600 23256 10606
rect 23032 10560 23204 10588
rect 23204 10542 23256 10548
rect 22940 9646 23060 9674
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22572 8362 22600 8842
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 22560 8356 22612 8362
rect 22560 8298 22612 8304
rect 22480 7806 22600 7834
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 21916 5636 21968 5642
rect 21916 5578 21968 5584
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 21914 4856 21970 4865
rect 21914 4791 21916 4800
rect 21968 4791 21970 4800
rect 21916 4762 21968 4768
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 22020 4690 22048 5102
rect 22098 4856 22154 4865
rect 22098 4791 22100 4800
rect 22152 4791 22154 4800
rect 22100 4762 22152 4768
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 21284 4010 21312 4626
rect 22098 4312 22154 4321
rect 22098 4247 22100 4256
rect 22152 4247 22154 4256
rect 22192 4276 22244 4282
rect 22100 4218 22152 4224
rect 22192 4218 22244 4224
rect 22204 4128 22232 4218
rect 22020 4100 22232 4128
rect 21454 4040 21510 4049
rect 21272 4004 21324 4010
rect 21454 3975 21510 3984
rect 21272 3946 21324 3952
rect 21284 3602 21312 3946
rect 21468 3942 21496 3975
rect 21456 3936 21508 3942
rect 21376 3896 21456 3924
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21284 3126 21312 3538
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21376 2854 21404 3896
rect 21456 3878 21508 3884
rect 21914 3768 21970 3777
rect 21914 3703 21916 3712
rect 21968 3703 21970 3712
rect 21916 3674 21968 3680
rect 21638 3632 21694 3641
rect 21638 3567 21640 3576
rect 21692 3567 21694 3576
rect 21916 3596 21968 3602
rect 21640 3538 21692 3544
rect 21916 3538 21968 3544
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21100 2502 21312 2530
rect 21468 2514 21496 2994
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 21100 1902 21128 2502
rect 21284 2378 21312 2502
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 21192 1970 21220 2314
rect 21928 2310 21956 3538
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22020 2122 22048 4100
rect 22112 4010 22324 4026
rect 22100 4004 22336 4010
rect 22152 3998 22284 4004
rect 22100 3946 22152 3952
rect 22284 3946 22336 3952
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22204 2825 22232 3674
rect 22296 2854 22324 3946
rect 22284 2848 22336 2854
rect 22190 2816 22246 2825
rect 22284 2790 22336 2796
rect 22190 2751 22246 2760
rect 22480 2310 22508 7210
rect 22572 4554 22600 7806
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22664 5574 22692 7754
rect 22744 7744 22796 7750
rect 22742 7712 22744 7721
rect 22796 7712 22798 7721
rect 22742 7647 22798 7656
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22756 2378 22784 4966
rect 22848 2990 22876 4966
rect 22940 3670 22968 8774
rect 23032 7818 23060 9646
rect 23216 9518 23244 10542
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 23202 9208 23258 9217
rect 23202 9143 23258 9152
rect 23216 9110 23244 9143
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23020 7812 23072 7818
rect 23020 7754 23072 7760
rect 23032 6254 23060 7754
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 23216 5642 23244 8774
rect 23308 8634 23336 11018
rect 23400 10441 23428 11766
rect 23584 11354 23612 12174
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23478 10840 23534 10849
rect 23478 10775 23480 10784
rect 23532 10775 23534 10784
rect 23480 10746 23532 10752
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23386 10432 23442 10441
rect 23386 10367 23442 10376
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23400 6934 23428 10367
rect 23584 10062 23612 10678
rect 23676 10266 23704 13738
rect 23768 12345 23796 13903
rect 23860 13870 23888 14282
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23952 13802 23980 17614
rect 24044 14890 24072 18838
rect 24136 18766 24164 19654
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 23940 13796 23992 13802
rect 23940 13738 23992 13744
rect 24044 13682 24072 14826
rect 23952 13654 24072 13682
rect 23754 12336 23810 12345
rect 23754 12271 23810 12280
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23492 7954 23520 8978
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23492 7478 23520 7890
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23204 5636 23256 5642
rect 23204 5578 23256 5584
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23124 3670 23152 4082
rect 22928 3664 22980 3670
rect 22928 3606 22980 3612
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 22940 3466 22968 3606
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 22744 2372 22796 2378
rect 22744 2314 22796 2320
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 21928 2094 22048 2122
rect 21180 1964 21232 1970
rect 21180 1906 21232 1912
rect 21088 1896 21140 1902
rect 21088 1838 21140 1844
rect 21928 800 21956 2094
rect 23216 1902 23244 5578
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 23308 3126 23336 5510
rect 23492 3641 23520 6190
rect 23584 3777 23612 9454
rect 23676 8566 23704 10202
rect 23768 9994 23796 12271
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23860 11898 23888 12106
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23860 11150 23888 11630
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23860 10810 23888 11086
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23860 10130 23888 10746
rect 23952 10305 23980 13654
rect 24136 13546 24164 18702
rect 24412 18290 24440 20198
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24412 18086 24440 18226
rect 24400 18080 24452 18086
rect 24400 18022 24452 18028
rect 24780 17814 24808 19246
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 24320 16794 24348 17614
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24044 13518 24164 13546
rect 24044 11880 24072 13518
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24136 12434 24164 12718
rect 24136 12406 24256 12434
rect 24044 11852 24164 11880
rect 24030 11792 24086 11801
rect 24030 11727 24086 11736
rect 24044 10810 24072 11727
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 23938 10296 23994 10305
rect 23938 10231 23994 10240
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23676 6934 23704 7278
rect 23664 6928 23716 6934
rect 23664 6870 23716 6876
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 23676 5778 23704 6326
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 23768 5370 23796 9930
rect 23860 8498 23888 10066
rect 24136 10010 24164 11852
rect 24228 10985 24256 12406
rect 24214 10976 24270 10985
rect 24214 10911 24270 10920
rect 24228 10606 24256 10911
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 23952 9982 24164 10010
rect 23952 9518 23980 9982
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 24044 9042 24072 9862
rect 24136 9654 24164 9862
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24320 8974 24348 16730
rect 24780 16658 24808 17750
rect 24872 17134 24900 18158
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 17270 24992 17478
rect 25056 17270 25084 20266
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 24860 17128 24912 17134
rect 25148 17082 25176 21354
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 24860 17070 24912 17076
rect 25056 17054 25176 17082
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24858 16552 24914 16561
rect 24858 16487 24914 16496
rect 24952 16516 25004 16522
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24780 15910 24808 15982
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24492 15428 24544 15434
rect 24544 15388 24808 15416
rect 24492 15370 24544 15376
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 24412 14618 24440 15030
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24582 14104 24638 14113
rect 24582 14039 24638 14048
rect 24596 13938 24624 14039
rect 24688 14006 24716 14214
rect 24780 14006 24808 15388
rect 24872 14226 24900 16487
rect 24952 16458 25004 16464
rect 24964 16046 24992 16458
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 25056 15026 25084 17054
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25148 16522 25176 16934
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 25240 15570 25268 16594
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 25240 15314 25268 15506
rect 25148 15286 25268 15314
rect 25148 15094 25176 15286
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25044 14544 25096 14550
rect 25148 14521 25176 14894
rect 25044 14486 25096 14492
rect 25134 14512 25190 14521
rect 24872 14198 24992 14226
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24412 11529 24440 11698
rect 24398 11520 24454 11529
rect 24398 11455 24454 11464
rect 24504 10130 24532 12718
rect 24596 12481 24624 13738
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24780 13258 24808 13670
rect 24964 13258 24992 14198
rect 25056 13938 25084 14486
rect 25134 14447 25190 14456
rect 25240 14278 25268 15098
rect 25332 14550 25360 20742
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25424 16561 25452 19246
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25516 18698 25544 18906
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25608 18358 25636 19654
rect 25872 19440 25924 19446
rect 25872 19382 25924 19388
rect 26056 19440 26108 19446
rect 26056 19382 26108 19388
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25700 18358 25728 18566
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25688 18352 25740 18358
rect 25688 18294 25740 18300
rect 25688 17264 25740 17270
rect 25688 17206 25740 17212
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25410 16552 25466 16561
rect 25410 16487 25466 16496
rect 25516 16250 25544 17070
rect 25608 16726 25636 17138
rect 25596 16720 25648 16726
rect 25596 16662 25648 16668
rect 25700 16522 25728 17206
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24582 12472 24638 12481
rect 24582 12407 24638 12416
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24596 11393 24624 11766
rect 24582 11384 24638 11393
rect 24582 11319 24638 11328
rect 24688 10985 24716 12582
rect 25134 12064 25190 12073
rect 25134 11999 25190 12008
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24674 10976 24730 10985
rect 24674 10911 24730 10920
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24308 8968 24360 8974
rect 24688 8922 24716 10911
rect 25056 10742 25084 11630
rect 25148 11082 25176 11999
rect 25240 11880 25268 14214
rect 25332 13870 25360 14214
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25424 12306 25452 15982
rect 25504 15972 25556 15978
rect 25504 15914 25556 15920
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 25240 11852 25452 11880
rect 25226 11792 25282 11801
rect 25226 11727 25282 11736
rect 25240 11082 25268 11727
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24858 10024 24914 10033
rect 24858 9959 24860 9968
rect 24912 9959 24914 9968
rect 24860 9930 24912 9936
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9722 24808 9862
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24308 8910 24360 8916
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 24320 8090 24348 8910
rect 24504 8894 24716 8922
rect 24858 8936 24914 8945
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24504 7970 24532 8894
rect 24858 8871 24860 8880
rect 24912 8871 24914 8880
rect 24860 8842 24912 8848
rect 24584 8832 24636 8838
rect 24636 8780 24716 8786
rect 24584 8774 24716 8780
rect 24596 8758 24716 8774
rect 24688 8430 24716 8758
rect 25044 8560 25096 8566
rect 25042 8528 25044 8537
rect 25096 8528 25098 8537
rect 25042 8463 25098 8472
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24320 7942 24532 7970
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23860 6322 23888 7414
rect 24044 6798 24072 7822
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23940 6724 23992 6730
rect 23940 6666 23992 6672
rect 23952 6633 23980 6666
rect 23938 6624 23994 6633
rect 23938 6559 23994 6568
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23860 5778 23888 6258
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23860 5137 23888 5306
rect 23846 5128 23902 5137
rect 23756 5092 23808 5098
rect 23846 5063 23902 5072
rect 23756 5034 23808 5040
rect 23570 3768 23626 3777
rect 23570 3703 23626 3712
rect 23478 3632 23534 3641
rect 23478 3567 23534 3576
rect 23768 3534 23796 5034
rect 23860 4622 23888 5063
rect 23952 4826 23980 6122
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24044 5710 24072 5850
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24044 5409 24072 5646
rect 24030 5400 24086 5409
rect 24030 5335 24086 5344
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23940 4480 23992 4486
rect 23940 4422 23992 4428
rect 23952 4214 23980 4422
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24044 3534 24072 3878
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23492 3346 23520 3402
rect 23400 3318 23520 3346
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23296 3120 23348 3126
rect 23296 3062 23348 3068
rect 23400 2582 23428 3318
rect 23388 2576 23440 2582
rect 23388 2518 23440 2524
rect 23204 1896 23256 1902
rect 23204 1838 23256 1844
rect 23860 800 23888 3334
rect 24320 3126 24348 7942
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 24490 7576 24546 7585
rect 24490 7511 24546 7520
rect 24504 7478 24532 7511
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24858 6760 24914 6769
rect 24858 6695 24914 6704
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 24400 5840 24452 5846
rect 24400 5782 24452 5788
rect 24412 5574 24440 5782
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24504 5234 24532 6598
rect 24872 6390 24900 6695
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24584 6248 24636 6254
rect 24582 6216 24584 6225
rect 24636 6216 24638 6225
rect 24582 6151 24638 6160
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24398 4992 24454 5001
rect 24398 4927 24454 4936
rect 24412 4214 24440 4927
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24412 3398 24440 4150
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24596 3126 24624 5102
rect 24688 4570 24716 6258
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24872 5778 24900 6054
rect 24964 5778 24992 6802
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 25056 5370 25084 7754
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 24964 5250 24992 5306
rect 25148 5250 25176 6734
rect 25318 5808 25374 5817
rect 25318 5743 25374 5752
rect 25332 5642 25360 5743
rect 25320 5636 25372 5642
rect 25320 5578 25372 5584
rect 24964 5222 25176 5250
rect 25148 5166 25176 5222
rect 25318 5264 25374 5273
rect 25318 5199 25374 5208
rect 25136 5160 25188 5166
rect 25136 5102 25188 5108
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24780 4729 24808 4762
rect 24766 4720 24822 4729
rect 24766 4655 24822 4664
rect 24952 4616 25004 4622
rect 24950 4584 24952 4593
rect 25004 4584 25006 4593
rect 24688 4542 24808 4570
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24688 2514 24716 4014
rect 24780 4010 24808 4542
rect 24950 4519 25006 4528
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 25056 4282 25084 4422
rect 25134 4312 25190 4321
rect 25044 4276 25096 4282
rect 25134 4247 25136 4256
rect 25044 4218 25096 4224
rect 25188 4247 25190 4256
rect 25136 4218 25188 4224
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24872 2106 24900 3062
rect 24964 2922 24992 3606
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 25056 2774 25084 4218
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 24964 2746 25084 2774
rect 24964 2378 24992 2746
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 24860 2100 24912 2106
rect 24860 2042 24912 2048
rect 25148 800 25176 4014
rect 25332 3466 25360 5199
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25424 2774 25452 11852
rect 25516 11098 25544 15914
rect 25792 15706 25820 18362
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 25780 15700 25832 15706
rect 25780 15642 25832 15648
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25608 15065 25636 15574
rect 25700 15366 25728 15642
rect 25780 15496 25832 15502
rect 25778 15464 25780 15473
rect 25832 15464 25834 15473
rect 25778 15399 25834 15408
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25594 15056 25650 15065
rect 25594 14991 25650 15000
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25608 13394 25636 14894
rect 25686 14648 25742 14657
rect 25686 14583 25742 14592
rect 25700 14414 25728 14583
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25688 14408 25740 14414
rect 25792 14385 25820 14418
rect 25688 14350 25740 14356
rect 25778 14376 25834 14385
rect 25778 14311 25834 14320
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25596 12912 25648 12918
rect 25594 12880 25596 12889
rect 25648 12880 25650 12889
rect 25594 12815 25650 12824
rect 25700 12434 25728 13330
rect 25700 12406 25820 12434
rect 25792 12170 25820 12406
rect 25780 12164 25832 12170
rect 25780 12106 25832 12112
rect 25516 11070 25728 11098
rect 25504 10736 25556 10742
rect 25504 10678 25556 10684
rect 25516 10198 25544 10678
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25700 9722 25728 11070
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25516 6866 25544 8774
rect 25608 8634 25636 9590
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25792 8294 25820 12106
rect 25884 9738 25912 19382
rect 26068 17882 26096 19382
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 25976 17202 26004 17818
rect 26056 17264 26108 17270
rect 26056 17206 26108 17212
rect 25964 17196 26016 17202
rect 25964 17138 26016 17144
rect 26068 16794 26096 17206
rect 26160 16794 26188 19790
rect 26712 19446 26740 25094
rect 27172 24682 27200 37198
rect 28368 37126 28396 39200
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 30300 37210 30328 39200
rect 30472 37256 30524 37262
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26700 19440 26752 19446
rect 26700 19382 26752 19388
rect 26712 18834 26740 19382
rect 26700 18828 26752 18834
rect 26700 18770 26752 18776
rect 26608 18148 26660 18154
rect 26608 18090 26660 18096
rect 26332 18080 26384 18086
rect 26332 18022 26384 18028
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26056 16788 26108 16794
rect 26056 16730 26108 16736
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 25964 15972 26016 15978
rect 25964 15914 26016 15920
rect 25976 13394 26004 15914
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 26068 15502 26096 15642
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26160 15065 26188 16730
rect 26252 16182 26280 17546
rect 26344 17542 26372 18022
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26424 17060 26476 17066
rect 26424 17002 26476 17008
rect 26332 16720 26384 16726
rect 26332 16662 26384 16668
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 26146 15056 26202 15065
rect 26146 14991 26202 15000
rect 26252 14634 26280 15982
rect 26344 14890 26372 16662
rect 26436 16182 26464 17002
rect 26528 16182 26556 17682
rect 26620 17678 26648 18090
rect 26608 17672 26660 17678
rect 26804 17660 26832 19722
rect 26896 19514 26924 19858
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 27172 18358 27200 18838
rect 27540 18358 27568 20266
rect 27816 18358 27844 27270
rect 28000 22094 28028 32370
rect 28000 22066 28120 22094
rect 27160 18352 27212 18358
rect 27160 18294 27212 18300
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27804 18352 27856 18358
rect 27804 18294 27856 18300
rect 27816 17814 27844 18294
rect 27804 17808 27856 17814
rect 27804 17750 27856 17756
rect 26884 17672 26936 17678
rect 26804 17632 26884 17660
rect 26608 17614 26660 17620
rect 26884 17614 26936 17620
rect 26608 16516 26660 16522
rect 26792 16516 26844 16522
rect 26660 16476 26792 16504
rect 26608 16458 26660 16464
rect 26792 16458 26844 16464
rect 26424 16176 26476 16182
rect 26424 16118 26476 16124
rect 26516 16176 26568 16182
rect 26516 16118 26568 16124
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26332 14884 26384 14890
rect 26332 14826 26384 14832
rect 26160 14606 26280 14634
rect 26056 14544 26108 14550
rect 26056 14486 26108 14492
rect 26068 14278 26096 14486
rect 26160 14482 26188 14606
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26252 14346 26280 14418
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 26160 14226 26188 14282
rect 26330 14240 26386 14249
rect 26160 14198 26280 14226
rect 26146 13968 26202 13977
rect 26146 13903 26202 13912
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25976 12434 26004 13194
rect 25976 12406 26096 12434
rect 25964 12368 26016 12374
rect 25964 12310 26016 12316
rect 25976 12209 26004 12310
rect 25962 12200 26018 12209
rect 25962 12135 26018 12144
rect 26068 11898 26096 12406
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 26056 11008 26108 11014
rect 26054 10976 26056 10985
rect 26108 10976 26110 10985
rect 26054 10911 26110 10920
rect 25884 9710 26004 9738
rect 25976 9654 26004 9710
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25884 7342 25912 8230
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 26160 7154 26188 13903
rect 26252 13818 26280 14198
rect 26330 14175 26386 14184
rect 26344 14006 26372 14175
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26436 13818 26464 13942
rect 26252 13790 26464 13818
rect 26528 13394 26556 14894
rect 26712 14414 26740 15302
rect 26700 14408 26752 14414
rect 26700 14350 26752 14356
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26436 12986 26464 13126
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26436 12306 26464 12922
rect 26528 12782 26556 13330
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26344 11218 26372 11834
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26252 10130 26280 11154
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26252 9586 26280 10066
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26252 8906 26280 9522
rect 26712 9518 26740 14350
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 26804 9994 26832 10202
rect 26792 9988 26844 9994
rect 26792 9930 26844 9936
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26712 9178 26740 9454
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 26620 8838 26648 9114
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26620 7970 26648 8774
rect 26896 8430 26924 17614
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27172 16998 27200 17138
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27080 16046 27108 16934
rect 27632 16522 27660 17478
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 26976 15904 27028 15910
rect 26976 15846 27028 15852
rect 26988 15434 27016 15846
rect 26976 15428 27028 15434
rect 26976 15370 27028 15376
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 27080 14890 27108 15030
rect 27068 14884 27120 14890
rect 27068 14826 27120 14832
rect 27172 14482 27200 16390
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27356 14618 27384 14894
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27068 14000 27120 14006
rect 27068 13942 27120 13948
rect 27080 12374 27108 13942
rect 27160 13796 27212 13802
rect 27160 13738 27212 13744
rect 27068 12368 27120 12374
rect 27068 12310 27120 12316
rect 27172 11830 27200 13738
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27080 11642 27108 11698
rect 27080 11614 27200 11642
rect 27264 11626 27292 14010
rect 27356 12306 27384 14282
rect 27528 13456 27580 13462
rect 27528 13398 27580 13404
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27448 12102 27476 13330
rect 27540 12986 27568 13398
rect 27632 13258 27660 15846
rect 27804 14884 27856 14890
rect 27804 14826 27856 14832
rect 27896 14884 27948 14890
rect 27896 14826 27948 14832
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27724 14006 27752 14758
rect 27816 14414 27844 14826
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27804 14272 27856 14278
rect 27804 14214 27856 14220
rect 27816 14006 27844 14214
rect 27712 14000 27764 14006
rect 27712 13942 27764 13948
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27816 13870 27844 13942
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 27712 13252 27764 13258
rect 27712 13194 27764 13200
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 27620 12708 27672 12714
rect 27724 12696 27752 13194
rect 27908 13190 27936 14826
rect 28000 14657 28028 17138
rect 28092 16046 28120 22066
rect 28460 20058 28488 37198
rect 30300 37182 30420 37210
rect 30472 37198 30524 37204
rect 30392 37126 30420 37182
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30484 35290 30512 37198
rect 32232 37126 32260 39200
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 29644 35080 29696 35086
rect 29644 35022 29696 35028
rect 30748 35080 30800 35086
rect 30748 35022 30800 35028
rect 29656 32366 29684 35022
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29656 25498 29684 32302
rect 30760 27470 30788 35022
rect 32600 32570 32628 37198
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37330 35480 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 35440 37324 35492 37330
rect 35440 37266 35492 37272
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33612 36922 33640 37198
rect 33600 36916 33652 36922
rect 33600 36858 33652 36864
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35820 36378 35848 37198
rect 36820 36780 36872 36786
rect 36820 36722 36872 36728
rect 36832 36582 36860 36722
rect 36820 36576 36872 36582
rect 36820 36518 36872 36524
rect 35808 36372 35860 36378
rect 35808 36314 35860 36320
rect 36728 36032 36780 36038
rect 36728 35974 36780 35980
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 32588 32564 32640 32570
rect 32588 32506 32640 32512
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 36740 29510 36768 35974
rect 36728 29504 36780 29510
rect 36728 29446 36780 29452
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 32036 25152 32088 25158
rect 32036 25094 32088 25100
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 28448 20052 28500 20058
rect 28448 19994 28500 20000
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 28908 18284 28960 18290
rect 28908 18226 28960 18232
rect 28356 17672 28408 17678
rect 28354 17640 28356 17649
rect 28408 17640 28410 17649
rect 28354 17575 28410 17584
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 28092 15434 28120 15982
rect 28080 15428 28132 15434
rect 28080 15370 28132 15376
rect 28092 14958 28120 15370
rect 28368 14958 28396 16594
rect 28460 15162 28488 17478
rect 28816 16652 28868 16658
rect 28816 16594 28868 16600
rect 28724 16176 28776 16182
rect 28724 16118 28776 16124
rect 28448 15156 28500 15162
rect 28448 15098 28500 15104
rect 28540 15088 28592 15094
rect 28540 15030 28592 15036
rect 28080 14952 28132 14958
rect 28080 14894 28132 14900
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 27986 14648 28042 14657
rect 27986 14583 28042 14592
rect 28368 14498 28396 14894
rect 28446 14512 28502 14521
rect 28080 14476 28132 14482
rect 28368 14470 28446 14498
rect 28446 14447 28502 14456
rect 28080 14418 28132 14424
rect 28092 14249 28120 14418
rect 28460 14414 28488 14447
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 28078 14240 28134 14249
rect 28078 14175 28134 14184
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27672 12668 27752 12696
rect 27620 12650 27672 12656
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27540 12170 27568 12582
rect 27618 12200 27674 12209
rect 27528 12164 27580 12170
rect 27618 12135 27620 12144
rect 27528 12106 27580 12112
rect 27672 12135 27674 12144
rect 27620 12106 27672 12112
rect 27436 12096 27488 12102
rect 27712 12096 27764 12102
rect 27436 12038 27488 12044
rect 27710 12064 27712 12073
rect 27764 12064 27766 12073
rect 27710 11999 27766 12008
rect 27816 11801 27844 12718
rect 27802 11792 27858 11801
rect 27802 11727 27858 11736
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27172 10130 27200 11614
rect 27252 11620 27304 11626
rect 27252 11562 27304 11568
rect 27710 11520 27766 11529
rect 27710 11455 27766 11464
rect 27724 11354 27752 11455
rect 27816 11354 27844 11630
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27804 11348 27856 11354
rect 27804 11290 27856 11296
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27436 10736 27488 10742
rect 27436 10678 27488 10684
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 10198 27292 10542
rect 27252 10192 27304 10198
rect 27252 10134 27304 10140
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 27356 9110 27384 9454
rect 27344 9104 27396 9110
rect 27344 9046 27396 9052
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26620 7942 26832 7970
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26332 7812 26384 7818
rect 26332 7754 26384 7760
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26252 7342 26280 7686
rect 26344 7546 26372 7754
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26608 7336 26660 7342
rect 26712 7324 26740 7822
rect 26804 7410 26832 7942
rect 26896 7546 26924 8366
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 26660 7296 26740 7324
rect 26608 7278 26660 7284
rect 25884 7126 26188 7154
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25884 4146 25912 7126
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 26068 6458 26096 6666
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 26252 6338 26280 6938
rect 26620 6866 26648 7278
rect 27172 6866 27200 7346
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26252 6310 26372 6338
rect 26240 6248 26292 6254
rect 26240 6190 26292 6196
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 25976 4010 26004 4626
rect 26252 4486 26280 6190
rect 26344 5846 26372 6310
rect 26332 5840 26384 5846
rect 26384 5788 26464 5794
rect 26332 5782 26464 5788
rect 26344 5766 26464 5782
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26344 5302 26372 5646
rect 26332 5296 26384 5302
rect 26332 5238 26384 5244
rect 26344 5166 26372 5238
rect 26332 5160 26384 5166
rect 26332 5102 26384 5108
rect 26344 4622 26372 5102
rect 26436 4690 26464 5766
rect 26528 5284 26556 6394
rect 26620 6254 26648 6802
rect 27264 6458 27292 7414
rect 27356 7154 27384 8434
rect 27448 7274 27476 10678
rect 27540 9654 27568 11018
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27632 10266 27660 10746
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 28000 9994 28028 10202
rect 28092 10130 28120 13806
rect 28264 13796 28316 13802
rect 28264 13738 28316 13744
rect 28276 13326 28304 13738
rect 28552 13569 28580 15030
rect 28630 14648 28686 14657
rect 28630 14583 28686 14592
rect 28538 13560 28594 13569
rect 28448 13524 28500 13530
rect 28644 13530 28672 14583
rect 28538 13495 28594 13504
rect 28632 13524 28684 13530
rect 28448 13466 28500 13472
rect 28632 13466 28684 13472
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28172 13184 28224 13190
rect 28172 13126 28224 13132
rect 28184 12782 28212 13126
rect 28460 12918 28488 13466
rect 28448 12912 28500 12918
rect 28448 12854 28500 12860
rect 28172 12776 28224 12782
rect 28172 12718 28224 12724
rect 28644 12434 28672 13466
rect 28552 12406 28672 12434
rect 28448 11688 28500 11694
rect 28354 11656 28410 11665
rect 28448 11630 28500 11636
rect 28354 11591 28410 11600
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28080 10124 28132 10130
rect 28080 10066 28132 10072
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 27528 9648 27580 9654
rect 27620 9648 27672 9654
rect 27528 9590 27580 9596
rect 27618 9616 27620 9625
rect 27672 9616 27674 9625
rect 27618 9551 27674 9560
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27724 8634 27752 9522
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27540 7954 27568 8366
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27436 7268 27488 7274
rect 27436 7210 27488 7216
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 27540 7154 27568 7210
rect 27356 7126 27568 7154
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 26620 5710 26648 6190
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 26608 5296 26660 5302
rect 26528 5256 26608 5284
rect 26608 5238 26660 5244
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26344 4214 26372 4558
rect 26620 4214 26648 5238
rect 27356 5234 27384 7126
rect 28000 6662 28028 9930
rect 28092 9926 28120 10066
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28092 5302 28120 9454
rect 28276 8786 28304 11494
rect 28368 8906 28396 11591
rect 28460 10810 28488 11630
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 28552 10606 28580 12406
rect 28736 12306 28764 16118
rect 28828 14113 28856 16594
rect 28814 14104 28870 14113
rect 28814 14039 28870 14048
rect 28920 13870 28948 18226
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 15910 29040 18022
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29012 14929 29040 14962
rect 28998 14920 29054 14929
rect 28998 14855 29054 14864
rect 29092 14544 29144 14550
rect 29092 14486 29144 14492
rect 29104 14385 29132 14486
rect 29090 14376 29146 14385
rect 29090 14311 29146 14320
rect 28908 13864 28960 13870
rect 28828 13812 28908 13818
rect 28828 13806 28960 13812
rect 28828 13790 28948 13806
rect 29196 13802 29224 19314
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29184 13796 29236 13802
rect 28828 12782 28856 13790
rect 29184 13738 29236 13744
rect 29092 13456 29144 13462
rect 29092 13398 29144 13404
rect 28908 13252 28960 13258
rect 28908 13194 28960 13200
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 28828 12374 28856 12718
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28724 12300 28776 12306
rect 28724 12242 28776 12248
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28736 10266 28764 10746
rect 28920 10266 28948 13194
rect 29104 12986 29132 13398
rect 29196 13326 29224 13738
rect 29184 13320 29236 13326
rect 29184 13262 29236 13268
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29012 11354 29040 12922
rect 29196 11830 29224 13262
rect 29184 11824 29236 11830
rect 29184 11766 29236 11772
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29104 10713 29132 11494
rect 29184 11280 29236 11286
rect 29184 11222 29236 11228
rect 29196 11082 29224 11222
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29090 10704 29146 10713
rect 29090 10639 29146 10648
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28460 9761 28488 9862
rect 28446 9752 28502 9761
rect 28446 9687 28502 9696
rect 28356 8900 28408 8906
rect 28356 8842 28408 8848
rect 28276 8758 28396 8786
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28276 6225 28304 8026
rect 28368 7546 28396 8758
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28460 6458 28488 9687
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28644 7818 28672 8230
rect 28632 7812 28684 7818
rect 28632 7754 28684 7760
rect 28538 7032 28594 7041
rect 28538 6967 28594 6976
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 28262 6216 28318 6225
rect 28262 6151 28318 6160
rect 28080 5296 28132 5302
rect 28080 5238 28132 5244
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 26332 4208 26384 4214
rect 26332 4150 26384 4156
rect 26608 4208 26660 4214
rect 26608 4150 26660 4156
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 25964 4004 26016 4010
rect 25964 3946 26016 3952
rect 25884 3890 25912 3946
rect 25884 3862 26188 3890
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25792 3233 25820 3402
rect 26160 3398 26188 3862
rect 26344 3602 26372 4150
rect 26620 4049 26648 4150
rect 27344 4072 27396 4078
rect 26606 4040 26662 4049
rect 27344 4014 27396 4020
rect 26606 3975 26662 3984
rect 26332 3596 26384 3602
rect 26332 3538 26384 3544
rect 26238 3496 26294 3505
rect 26238 3431 26294 3440
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 25778 3224 25834 3233
rect 25778 3159 25834 3168
rect 26252 2990 26280 3431
rect 26344 3126 26372 3538
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26700 2984 26752 2990
rect 26700 2926 26752 2932
rect 26712 2854 26740 2926
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 25424 2746 25912 2774
rect 25884 2106 25912 2746
rect 26896 2582 26924 3334
rect 27356 3126 27384 4014
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28460 3738 28488 3878
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 25964 2576 26016 2582
rect 25964 2518 26016 2524
rect 26884 2576 26936 2582
rect 26884 2518 26936 2524
rect 25976 2310 26004 2518
rect 27080 2446 27108 2994
rect 28552 2774 28580 6967
rect 28736 5642 28764 8230
rect 29000 7472 29052 7478
rect 29000 7414 29052 7420
rect 29012 7313 29040 7414
rect 28998 7304 29054 7313
rect 28998 7239 29054 7248
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 7002 29040 7142
rect 29104 7002 29132 9318
rect 29196 8906 29224 9318
rect 29184 8900 29236 8906
rect 29184 8842 29236 8848
rect 29288 8514 29316 16934
rect 29552 15972 29604 15978
rect 29552 15914 29604 15920
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29472 15162 29500 15846
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29380 10606 29408 14962
rect 29472 14770 29500 15098
rect 29564 14890 29592 15914
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29552 14884 29604 14890
rect 29552 14826 29604 14832
rect 29472 14742 29592 14770
rect 29460 12776 29512 12782
rect 29460 12718 29512 12724
rect 29472 11830 29500 12718
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29564 11676 29592 14742
rect 29748 14278 29776 15438
rect 29932 15162 29960 24550
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 30196 15428 30248 15434
rect 30196 15370 30248 15376
rect 29920 15156 29972 15162
rect 29920 15098 29972 15104
rect 29932 14414 29960 15098
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29736 14272 29788 14278
rect 29736 14214 29788 14220
rect 29748 13938 29776 14214
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29656 12442 29684 13806
rect 29736 13728 29788 13734
rect 29736 13670 29788 13676
rect 29748 12850 29776 13670
rect 29840 12918 29868 13806
rect 29828 12912 29880 12918
rect 29828 12854 29880 12860
rect 29736 12844 29788 12850
rect 29736 12786 29788 12792
rect 29932 12730 29960 13942
rect 29840 12702 29960 12730
rect 29644 12436 29696 12442
rect 29644 12378 29696 12384
rect 29734 12336 29790 12345
rect 29734 12271 29790 12280
rect 29748 12238 29776 12271
rect 29736 12232 29788 12238
rect 29736 12174 29788 12180
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 29656 11801 29684 12106
rect 29642 11792 29698 11801
rect 29642 11727 29698 11736
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29472 11648 29592 11676
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 29380 9178 29408 10542
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29196 8498 29408 8514
rect 29196 8492 29420 8498
rect 29196 8486 29368 8492
rect 29000 6996 29052 7002
rect 29000 6938 29052 6944
rect 29092 6996 29144 7002
rect 29092 6938 29144 6944
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28724 5636 28776 5642
rect 28724 5578 28776 5584
rect 28724 4276 28776 4282
rect 28724 4218 28776 4224
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 2990 28672 3878
rect 28736 3058 28764 4218
rect 28828 3126 28856 6394
rect 28906 6080 28962 6089
rect 28906 6015 28962 6024
rect 28920 5846 28948 6015
rect 28908 5840 28960 5846
rect 28908 5782 28960 5788
rect 28920 4554 28948 5782
rect 29196 5166 29224 8486
rect 29368 8434 29420 8440
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 29288 8294 29316 8366
rect 29276 8288 29328 8294
rect 29276 8230 29328 8236
rect 29472 7818 29500 11648
rect 29748 11234 29776 11698
rect 29564 11206 29776 11234
rect 29564 9926 29592 11206
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29656 9654 29684 9998
rect 29748 9926 29776 11086
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29644 8900 29696 8906
rect 29644 8842 29696 8848
rect 29550 8664 29606 8673
rect 29550 8599 29606 8608
rect 29564 8566 29592 8599
rect 29552 8560 29604 8566
rect 29552 8502 29604 8508
rect 29550 8392 29606 8401
rect 29550 8327 29552 8336
rect 29604 8327 29606 8336
rect 29552 8298 29604 8304
rect 29460 7812 29512 7818
rect 29460 7754 29512 7760
rect 29472 7562 29500 7754
rect 29472 7534 29592 7562
rect 29564 7478 29592 7534
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 29276 6112 29328 6118
rect 29276 6054 29328 6060
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 28908 4548 28960 4554
rect 28908 4490 28960 4496
rect 29012 4146 29040 4558
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28632 2984 28684 2990
rect 28632 2926 28684 2932
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28552 2746 28672 2774
rect 28644 2650 28672 2746
rect 28540 2644 28592 2650
rect 28540 2586 28592 2592
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 25964 2304 26016 2310
rect 25964 2246 26016 2252
rect 25872 2100 25924 2106
rect 25872 2042 25924 2048
rect 27080 800 27108 2382
rect 27620 2304 27672 2310
rect 27620 2246 27672 2252
rect 27632 2038 27660 2246
rect 27620 2032 27672 2038
rect 27620 1974 27672 1980
rect 28552 1970 28580 2586
rect 28920 2514 28948 2926
rect 29000 2916 29052 2922
rect 29000 2858 29052 2864
rect 28908 2508 28960 2514
rect 28908 2450 28960 2456
rect 28540 1964 28592 1970
rect 28540 1906 28592 1912
rect 29012 800 29040 2858
rect 29288 2310 29316 6054
rect 29380 4078 29408 6326
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29564 3126 29592 7414
rect 29552 3120 29604 3126
rect 29552 3062 29604 3068
rect 29656 2990 29684 8842
rect 29748 8294 29776 9862
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29748 6254 29776 6734
rect 29840 6390 29868 12702
rect 30024 12594 30052 14486
rect 29932 12566 30052 12594
rect 29932 11150 29960 12566
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 30024 10606 30052 11018
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 30024 10130 30052 10542
rect 30012 10124 30064 10130
rect 30012 10066 30064 10072
rect 30024 10010 30052 10066
rect 29932 9982 30052 10010
rect 29932 9518 29960 9982
rect 30012 9648 30064 9654
rect 30012 9590 30064 9596
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 29932 9042 29960 9454
rect 29920 9036 29972 9042
rect 29920 8978 29972 8984
rect 30024 6390 30052 9590
rect 29828 6384 29880 6390
rect 29828 6326 29880 6332
rect 30012 6384 30064 6390
rect 30012 6326 30064 6332
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 29748 5778 29776 6190
rect 29736 5772 29788 5778
rect 29736 5714 29788 5720
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 29748 4622 29776 5714
rect 30024 5370 30052 5714
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 30116 5234 30144 14962
rect 30208 14074 30236 15370
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30392 14958 30420 15302
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 30300 14346 30328 14758
rect 30288 14340 30340 14346
rect 30288 14282 30340 14288
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30196 13184 30248 13190
rect 30196 13126 30248 13132
rect 30208 12646 30236 13126
rect 30392 12986 30420 14214
rect 30470 14104 30526 14113
rect 30470 14039 30472 14048
rect 30524 14039 30526 14048
rect 30472 14010 30524 14016
rect 30748 13320 30800 13326
rect 30748 13262 30800 13268
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30380 12980 30432 12986
rect 30380 12922 30432 12928
rect 30196 12640 30248 12646
rect 30196 12582 30248 12588
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30208 11694 30236 12174
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30378 11384 30434 11393
rect 30378 11319 30434 11328
rect 30392 11150 30420 11319
rect 30484 11286 30512 13126
rect 30564 12164 30616 12170
rect 30564 12106 30616 12112
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 30196 10464 30248 10470
rect 30196 10406 30248 10412
rect 30208 10198 30236 10406
rect 30300 10266 30328 10950
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30300 8498 30328 8774
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30392 7954 30420 11086
rect 30472 11008 30524 11014
rect 30472 10950 30524 10956
rect 30484 9926 30512 10950
rect 30472 9920 30524 9926
rect 30472 9862 30524 9868
rect 30576 9654 30604 12106
rect 30564 9648 30616 9654
rect 30564 9590 30616 9596
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30668 9382 30696 9590
rect 30656 9376 30708 9382
rect 30656 9318 30708 9324
rect 30760 9194 30788 13262
rect 30944 12986 30972 18906
rect 32048 16153 32076 25094
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34060 22636 34112 22642
rect 34060 22578 34112 22584
rect 34072 19514 34100 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34060 19508 34112 19514
rect 34060 19450 34112 19456
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 32034 16144 32090 16153
rect 31392 16108 31444 16114
rect 32034 16079 32090 16088
rect 31392 16050 31444 16056
rect 31300 15360 31352 15366
rect 31300 15302 31352 15308
rect 31312 15162 31340 15302
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31208 14272 31260 14278
rect 31208 14214 31260 14220
rect 31114 13560 31170 13569
rect 31114 13495 31116 13504
rect 31168 13495 31170 13504
rect 31116 13466 31168 13472
rect 31220 13394 31248 14214
rect 31208 13388 31260 13394
rect 31208 13330 31260 13336
rect 30932 12980 30984 12986
rect 30932 12922 30984 12928
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 30930 11792 30986 11801
rect 30930 11727 30932 11736
rect 30984 11727 30986 11736
rect 30932 11698 30984 11704
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30944 10470 30972 10746
rect 30932 10464 30984 10470
rect 30932 10406 30984 10412
rect 30932 9376 30984 9382
rect 30932 9318 30984 9324
rect 30668 9166 30788 9194
rect 30564 8900 30616 8906
rect 30564 8842 30616 8848
rect 30576 8566 30604 8842
rect 30564 8560 30616 8566
rect 30564 8502 30616 8508
rect 30380 7948 30432 7954
rect 30380 7890 30432 7896
rect 30668 7546 30696 9166
rect 30944 9042 30972 9318
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30932 8832 30984 8838
rect 30932 8774 30984 8780
rect 30840 8356 30892 8362
rect 30840 8298 30892 8304
rect 30656 7540 30708 7546
rect 30656 7482 30708 7488
rect 30656 7268 30708 7274
rect 30656 7210 30708 7216
rect 30288 6724 30340 6730
rect 30288 6666 30340 6672
rect 30472 6724 30524 6730
rect 30472 6666 30524 6672
rect 30300 6322 30328 6666
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30300 6100 30328 6258
rect 30380 6112 30432 6118
rect 30300 6072 30380 6100
rect 30380 6054 30432 6060
rect 30484 5681 30512 6666
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30470 5672 30526 5681
rect 30470 5607 30526 5616
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 30576 5166 30604 6258
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30564 5160 30616 5166
rect 30564 5102 30616 5108
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 29748 3602 29776 4558
rect 29736 3596 29788 3602
rect 29736 3538 29788 3544
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 30392 2922 30420 5102
rect 30668 4826 30696 7210
rect 30852 7206 30880 8298
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 30656 4820 30708 4826
rect 30656 4762 30708 4768
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 29276 2304 29328 2310
rect 29276 2246 29328 2252
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30300 800 30328 2246
rect 30944 2038 30972 8774
rect 31036 5778 31064 12174
rect 31128 11898 31156 12174
rect 31220 12102 31248 12786
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31116 11688 31168 11694
rect 31116 11630 31168 11636
rect 31024 5772 31076 5778
rect 31024 5714 31076 5720
rect 31024 5568 31076 5574
rect 31024 5510 31076 5516
rect 31036 2394 31064 5510
rect 31128 3942 31156 11630
rect 31220 8022 31248 11698
rect 31312 8906 31340 12854
rect 31300 8900 31352 8906
rect 31300 8842 31352 8848
rect 31208 8016 31260 8022
rect 31208 7958 31260 7964
rect 31220 4434 31248 7958
rect 31300 7812 31352 7818
rect 31300 7754 31352 7760
rect 31312 4622 31340 7754
rect 31404 5846 31432 16050
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 36832 15706 36860 36518
rect 37200 36378 37228 38791
rect 37384 36922 37412 39200
rect 38290 37496 38346 37505
rect 38290 37431 38346 37440
rect 38304 37330 38332 37431
rect 38292 37324 38344 37330
rect 38292 37266 38344 37272
rect 37832 37256 37884 37262
rect 37832 37198 37884 37204
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 37464 35624 37516 35630
rect 37464 35566 37516 35572
rect 37740 35624 37792 35630
rect 37740 35566 37792 35572
rect 37476 35465 37504 35566
rect 37462 35456 37518 35465
rect 37462 35391 37518 35400
rect 37752 35086 37780 35566
rect 37740 35080 37792 35086
rect 37740 35022 37792 35028
rect 37844 29646 37872 37198
rect 38304 36922 38332 37266
rect 38292 36916 38344 36922
rect 38292 36858 38344 36864
rect 38672 36378 38700 39200
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 38028 35290 38056 36110
rect 38016 35284 38068 35290
rect 38016 35226 38068 35232
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38292 32360 38344 32366
rect 38292 32302 38344 32308
rect 38304 32065 38332 32302
rect 38290 32056 38346 32065
rect 38290 31991 38292 32000
rect 38344 31991 38346 32000
rect 38292 31962 38344 31968
rect 38016 30252 38068 30258
rect 38016 30194 38068 30200
rect 38028 29850 38056 30194
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38016 29844 38068 29850
rect 38016 29786 38068 29792
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 37844 25294 37872 29582
rect 38198 27976 38254 27985
rect 38198 27911 38200 27920
rect 38252 27911 38254 27920
rect 38200 27882 38252 27888
rect 38016 27668 38068 27674
rect 38016 27610 38068 27616
rect 38028 27062 38056 27610
rect 38016 27056 38068 27062
rect 38016 26998 38068 27004
rect 38200 26988 38252 26994
rect 38200 26930 38252 26936
rect 38212 26625 38240 26930
rect 38198 26616 38254 26625
rect 38198 26551 38254 26560
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 38016 24812 38068 24818
rect 38016 24754 38068 24760
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37476 21350 37504 21490
rect 37464 21344 37516 21350
rect 37464 21286 37516 21292
rect 37476 19922 37504 21286
rect 38028 20806 38056 24754
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38016 20800 38068 20806
rect 38016 20742 38068 20748
rect 37464 19916 37516 19922
rect 37464 19858 37516 19864
rect 38016 19372 38068 19378
rect 38016 19314 38068 19320
rect 38028 18426 38056 19314
rect 38200 19168 38252 19174
rect 38198 19136 38200 19145
rect 38252 19136 38254 19145
rect 38198 19071 38254 19080
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 38200 17196 38252 17202
rect 38200 17138 38252 17144
rect 38212 17105 38240 17138
rect 38198 17096 38254 17105
rect 38016 17060 38068 17066
rect 38198 17031 38254 17040
rect 38016 17002 38068 17008
rect 36820 15700 36872 15706
rect 36820 15642 36872 15648
rect 33968 15156 34020 15162
rect 33968 15098 34020 15104
rect 31576 13864 31628 13870
rect 31576 13806 31628 13812
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31496 7750 31524 12038
rect 31588 11898 31616 13806
rect 31668 12096 31720 12102
rect 31668 12038 31720 12044
rect 31576 11892 31628 11898
rect 31576 11834 31628 11840
rect 31680 11082 31708 12038
rect 32312 11824 32364 11830
rect 32312 11766 32364 11772
rect 32324 11558 32352 11766
rect 32312 11552 32364 11558
rect 32312 11494 32364 11500
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31680 10810 31708 11018
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 32036 10464 32088 10470
rect 32036 10406 32088 10412
rect 32048 10266 32076 10406
rect 32036 10260 32088 10266
rect 32036 10202 32088 10208
rect 32324 10198 32352 11494
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32312 10192 32364 10198
rect 32312 10134 32364 10140
rect 32416 9586 32444 11154
rect 33152 10742 33180 13806
rect 33232 12844 33284 12850
rect 33232 12786 33284 12792
rect 33140 10736 33192 10742
rect 33140 10678 33192 10684
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33152 10130 33180 10406
rect 33140 10124 33192 10130
rect 33140 10066 33192 10072
rect 32772 9648 32824 9654
rect 32772 9590 32824 9596
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32784 9110 32812 9590
rect 33152 9586 33180 10066
rect 33140 9580 33192 9586
rect 33140 9522 33192 9528
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 32772 9104 32824 9110
rect 32772 9046 32824 9052
rect 31576 9036 31628 9042
rect 31576 8978 31628 8984
rect 31588 8362 31616 8978
rect 32588 8900 32640 8906
rect 32588 8842 32640 8848
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 31576 8356 31628 8362
rect 31576 8298 31628 8304
rect 31484 7744 31536 7750
rect 31484 7686 31536 7692
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 31496 7002 31524 7686
rect 31956 7342 31984 7686
rect 31944 7336 31996 7342
rect 31944 7278 31996 7284
rect 31576 7268 31628 7274
rect 31576 7210 31628 7216
rect 32036 7268 32088 7274
rect 32036 7210 32088 7216
rect 31484 6996 31536 7002
rect 31484 6938 31536 6944
rect 31588 6866 31616 7210
rect 32048 7002 32076 7210
rect 32036 6996 32088 7002
rect 32036 6938 32088 6944
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 31576 6384 31628 6390
rect 31628 6332 31708 6338
rect 31576 6326 31708 6332
rect 31588 6310 31708 6326
rect 31576 6180 31628 6186
rect 31576 6122 31628 6128
rect 31588 5914 31616 6122
rect 31680 5914 31708 6310
rect 31944 6248 31996 6254
rect 31944 6190 31996 6196
rect 31576 5908 31628 5914
rect 31576 5850 31628 5856
rect 31668 5908 31720 5914
rect 31668 5850 31720 5856
rect 31392 5840 31444 5846
rect 31392 5782 31444 5788
rect 31956 5778 31984 6190
rect 31944 5772 31996 5778
rect 31944 5714 31996 5720
rect 31484 5228 31536 5234
rect 31484 5170 31536 5176
rect 31392 4684 31444 4690
rect 31392 4626 31444 4632
rect 31300 4616 31352 4622
rect 31300 4558 31352 4564
rect 31220 4406 31340 4434
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 31116 3664 31168 3670
rect 31116 3606 31168 3612
rect 31128 3126 31156 3606
rect 31220 3602 31248 4014
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31312 3126 31340 4406
rect 31404 3398 31432 4626
rect 31496 4146 31524 5170
rect 32140 5030 32168 8774
rect 32600 8362 32628 8842
rect 33060 8673 33088 9318
rect 33046 8664 33102 8673
rect 33046 8599 33102 8608
rect 32588 8356 32640 8362
rect 32588 8298 32640 8304
rect 33152 7478 33180 9522
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 32692 7041 32720 7142
rect 32218 7032 32274 7041
rect 32218 6967 32274 6976
rect 32678 7032 32734 7041
rect 32678 6967 32734 6976
rect 32128 5024 32180 5030
rect 32128 4966 32180 4972
rect 31576 4480 31628 4486
rect 31576 4422 31628 4428
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 31392 3392 31444 3398
rect 31496 3380 31524 3878
rect 31588 3738 31616 4422
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 31668 4004 31720 4010
rect 31668 3946 31720 3952
rect 31944 4004 31996 4010
rect 31944 3946 31996 3952
rect 31680 3738 31708 3946
rect 31576 3732 31628 3738
rect 31576 3674 31628 3680
rect 31668 3732 31720 3738
rect 31668 3674 31720 3680
rect 31760 3664 31812 3670
rect 31812 3624 31892 3652
rect 31760 3606 31812 3612
rect 31576 3392 31628 3398
rect 31496 3352 31576 3380
rect 31392 3334 31444 3340
rect 31576 3334 31628 3340
rect 31758 3224 31814 3233
rect 31758 3159 31760 3168
rect 31812 3159 31814 3168
rect 31760 3130 31812 3136
rect 31116 3120 31168 3126
rect 31116 3062 31168 3068
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 31300 2984 31352 2990
rect 31298 2952 31300 2961
rect 31352 2952 31354 2961
rect 31298 2887 31354 2896
rect 31758 2952 31814 2961
rect 31864 2922 31892 3624
rect 31956 3466 31984 3946
rect 31944 3460 31996 3466
rect 31944 3402 31996 3408
rect 31944 3188 31996 3194
rect 31944 3130 31996 3136
rect 31758 2887 31760 2896
rect 31812 2887 31814 2896
rect 31852 2916 31904 2922
rect 31760 2858 31812 2864
rect 31852 2858 31904 2864
rect 31772 2802 31800 2858
rect 31956 2802 31984 3130
rect 32140 2990 32168 4014
rect 32232 3466 32260 6967
rect 32496 6656 32548 6662
rect 32496 6598 32548 6604
rect 32508 6118 32536 6598
rect 33152 6186 33180 7414
rect 33140 6180 33192 6186
rect 33140 6122 33192 6128
rect 32496 6112 32548 6118
rect 32496 6054 32548 6060
rect 32508 5234 32536 6054
rect 32496 5228 32548 5234
rect 32496 5170 32548 5176
rect 32312 5092 32364 5098
rect 32312 5034 32364 5040
rect 32324 4622 32352 5034
rect 32772 5024 32824 5030
rect 32772 4966 32824 4972
rect 32864 5024 32916 5030
rect 32864 4966 32916 4972
rect 32680 4752 32732 4758
rect 32680 4694 32732 4700
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 32220 3460 32272 3466
rect 32220 3402 32272 3408
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 31772 2774 31984 2802
rect 32140 2514 32168 2926
rect 32324 2774 32352 4558
rect 32232 2746 32352 2774
rect 32128 2508 32180 2514
rect 32128 2450 32180 2456
rect 31036 2372 31432 2394
rect 31036 2366 31116 2372
rect 31168 2366 31432 2372
rect 31116 2314 31168 2320
rect 31404 2310 31432 2366
rect 31392 2304 31444 2310
rect 31392 2246 31444 2252
rect 30932 2032 30984 2038
rect 30932 1974 30984 1980
rect 32232 800 32260 2746
rect 32692 2582 32720 4694
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 32784 2378 32812 4966
rect 32876 4282 32904 4966
rect 33244 4826 33272 12786
rect 33508 11280 33560 11286
rect 33508 11222 33560 11228
rect 33416 11144 33468 11150
rect 33416 11086 33468 11092
rect 33428 10810 33456 11086
rect 33416 10804 33468 10810
rect 33416 10746 33468 10752
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33428 7274 33456 7686
rect 33416 7268 33468 7274
rect 33416 7210 33468 7216
rect 33428 6662 33456 7210
rect 33416 6656 33468 6662
rect 33416 6598 33468 6604
rect 33428 6186 33456 6598
rect 33416 6180 33468 6186
rect 33416 6122 33468 6128
rect 33232 4820 33284 4826
rect 33232 4762 33284 4768
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 33244 4146 33272 4762
rect 33324 4684 33376 4690
rect 33324 4626 33376 4632
rect 33232 4140 33284 4146
rect 33232 4082 33284 4088
rect 33232 3664 33284 3670
rect 33232 3606 33284 3612
rect 33244 3194 33272 3606
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 33336 2774 33364 4626
rect 33428 4554 33456 6122
rect 33416 4548 33468 4554
rect 33416 4490 33468 4496
rect 33428 4282 33456 4490
rect 33520 4486 33548 11222
rect 33600 9376 33652 9382
rect 33600 9318 33652 9324
rect 33612 8906 33640 9318
rect 33600 8900 33652 8906
rect 33600 8842 33652 8848
rect 33600 8288 33652 8294
rect 33600 8230 33652 8236
rect 33612 6458 33640 8230
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33600 6452 33652 6458
rect 33600 6394 33652 6400
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33508 3936 33560 3942
rect 33508 3878 33560 3884
rect 33520 2774 33548 3878
rect 33704 3670 33732 6598
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33888 3738 33916 3878
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 33980 3670 34008 15098
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 36820 14272 36872 14278
rect 36820 14214 36872 14220
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9716 34848 9722
rect 34796 9658 34848 9664
rect 34520 8356 34572 8362
rect 34520 8298 34572 8304
rect 34060 6316 34112 6322
rect 34060 6258 34112 6264
rect 34072 5778 34100 6258
rect 34532 6118 34560 8298
rect 34808 7546 34836 9658
rect 36084 9444 36136 9450
rect 36084 9386 36136 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 36096 8974 36124 9386
rect 36084 8968 36136 8974
rect 36084 8910 36136 8916
rect 35992 8900 36044 8906
rect 35992 8842 36044 8848
rect 36004 8401 36032 8842
rect 35990 8392 36046 8401
rect 35990 8327 36046 8336
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 36096 8090 36124 8910
rect 36832 8498 36860 14214
rect 37096 13388 37148 13394
rect 37096 13330 37148 13336
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36096 7886 36124 8026
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 36096 7546 36124 7822
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 36084 7540 36136 7546
rect 36084 7482 36136 7488
rect 34612 7336 34664 7342
rect 34612 7278 34664 7284
rect 34704 7336 34756 7342
rect 34704 7278 34756 7284
rect 34624 6866 34652 7278
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34520 6112 34572 6118
rect 34520 6054 34572 6060
rect 34532 5846 34560 6054
rect 34520 5840 34572 5846
rect 34520 5782 34572 5788
rect 34060 5772 34112 5778
rect 34060 5714 34112 5720
rect 34532 4622 34560 5782
rect 34624 5370 34652 6802
rect 34716 5642 34744 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35440 6860 35492 6866
rect 35440 6802 35492 6808
rect 35452 6322 35480 6802
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34704 5636 34756 5642
rect 34704 5578 34756 5584
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 34808 5030 34836 5510
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34072 4282 34100 4558
rect 34152 4480 34204 4486
rect 34808 4468 34836 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34888 4480 34940 4486
rect 34808 4440 34888 4468
rect 34152 4422 34204 4428
rect 34888 4422 34940 4428
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 33692 3664 33744 3670
rect 33692 3606 33744 3612
rect 33968 3664 34020 3670
rect 33968 3606 34020 3612
rect 34164 3466 34192 4422
rect 34336 4004 34388 4010
rect 34336 3946 34388 3952
rect 34152 3460 34204 3466
rect 34152 3402 34204 3408
rect 34244 3460 34296 3466
rect 34244 3402 34296 3408
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33612 3194 33640 3334
rect 33704 3233 33732 3334
rect 33690 3224 33746 3233
rect 33600 3188 33652 3194
rect 33690 3159 33746 3168
rect 33600 3130 33652 3136
rect 34152 2848 34204 2854
rect 34152 2790 34204 2796
rect 33336 2746 33456 2774
rect 33520 2746 33732 2774
rect 33428 2650 33456 2746
rect 33704 2650 33732 2746
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 32772 2372 32824 2378
rect 32772 2314 32824 2320
rect 34164 800 34192 2790
rect 34256 2582 34284 3402
rect 34244 2576 34296 2582
rect 34244 2518 34296 2524
rect 34348 2446 34376 3946
rect 34900 3942 34928 4422
rect 34888 3936 34940 3942
rect 34888 3878 34940 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35360 2990 35388 6054
rect 35544 3058 35572 7482
rect 35624 7268 35676 7274
rect 35624 7210 35676 7216
rect 35636 5914 35664 7210
rect 35716 7200 35768 7206
rect 35716 7142 35768 7148
rect 35624 5908 35676 5914
rect 35624 5850 35676 5856
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34428 2644 34480 2650
rect 34428 2586 34480 2592
rect 34336 2440 34388 2446
rect 34336 2382 34388 2388
rect 34440 2378 34468 2586
rect 35728 2446 35756 7142
rect 36096 7002 36124 7482
rect 36084 6996 36136 7002
rect 36084 6938 36136 6944
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35820 5846 35848 6598
rect 35808 5840 35860 5846
rect 35808 5782 35860 5788
rect 35820 5370 35848 5782
rect 35808 5364 35860 5370
rect 35808 5306 35860 5312
rect 36084 4548 36136 4554
rect 36084 4490 36136 4496
rect 36096 3942 36124 4490
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 36280 4214 36308 4422
rect 36268 4208 36320 4214
rect 36268 4150 36320 4156
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 36096 3466 36124 3878
rect 36084 3460 36136 3466
rect 36084 3402 36136 3408
rect 36096 3194 36124 3402
rect 36372 3398 36400 8298
rect 36634 7984 36690 7993
rect 36634 7919 36636 7928
rect 36688 7919 36690 7928
rect 36636 7890 36688 7896
rect 36636 6656 36688 6662
rect 36636 6598 36688 6604
rect 36648 5234 36676 6598
rect 37108 5914 37136 13330
rect 37924 13184 37976 13190
rect 37924 13126 37976 13132
rect 37556 9376 37608 9382
rect 37556 9318 37608 9324
rect 37568 8974 37596 9318
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37188 8424 37240 8430
rect 37188 8366 37240 8372
rect 37200 8265 37228 8366
rect 37186 8256 37242 8265
rect 37186 8191 37242 8200
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 37096 5908 37148 5914
rect 37096 5850 37148 5856
rect 36636 5228 36688 5234
rect 36636 5170 36688 5176
rect 36636 4004 36688 4010
rect 36636 3946 36688 3952
rect 36360 3392 36412 3398
rect 36360 3334 36412 3340
rect 36084 3188 36136 3194
rect 36084 3130 36136 3136
rect 36372 3058 36400 3334
rect 36648 3126 36676 3946
rect 36636 3120 36688 3126
rect 36636 3062 36688 3068
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 37108 2582 37136 5850
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 37384 3670 37412 4218
rect 37372 3664 37424 3670
rect 37372 3606 37424 3612
rect 37096 2576 37148 2582
rect 37096 2518 37148 2524
rect 37476 2446 37504 7686
rect 37568 7478 37596 8910
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37556 7472 37608 7478
rect 37556 7414 37608 7420
rect 37844 7002 37872 7822
rect 37832 6996 37884 7002
rect 37832 6938 37884 6944
rect 37844 4622 37872 6938
rect 37936 5302 37964 13126
rect 38028 12986 38056 17002
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38108 15904 38160 15910
rect 38108 15846 38160 15852
rect 38120 15570 38148 15846
rect 38212 15745 38240 16050
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38108 15564 38160 15570
rect 38108 15506 38160 15512
rect 38108 14816 38160 14822
rect 38108 14758 38160 14764
rect 38016 12980 38068 12986
rect 38016 12922 38068 12928
rect 38120 12866 38148 14758
rect 38292 13864 38344 13870
rect 38292 13806 38344 13812
rect 38304 13705 38332 13806
rect 38290 13696 38346 13705
rect 38290 13631 38346 13640
rect 38304 13530 38332 13631
rect 38292 13524 38344 13530
rect 38292 13466 38344 13472
rect 38028 12838 38148 12866
rect 38028 6390 38056 12838
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38212 11665 38240 11698
rect 38198 11656 38254 11665
rect 38198 11591 38254 11600
rect 38292 10668 38344 10674
rect 38292 10610 38344 10616
rect 38304 10305 38332 10610
rect 38290 10296 38346 10305
rect 38290 10231 38346 10240
rect 38292 9376 38344 9382
rect 38292 9318 38344 9324
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 38212 7002 38240 7346
rect 38200 6996 38252 7002
rect 38200 6938 38252 6944
rect 38212 6474 38240 6938
rect 38120 6446 38240 6474
rect 38016 6384 38068 6390
rect 38016 6326 38068 6332
rect 38120 5914 38148 6446
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38212 6225 38240 6258
rect 38198 6216 38254 6225
rect 38198 6151 38254 6160
rect 38108 5908 38160 5914
rect 38108 5850 38160 5856
rect 37924 5296 37976 5302
rect 37924 5238 37976 5244
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37844 4146 37872 4558
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37556 4072 37608 4078
rect 37556 4014 37608 4020
rect 37568 3534 37596 4014
rect 37556 3528 37608 3534
rect 37556 3470 37608 3476
rect 37556 3392 37608 3398
rect 37556 3334 37608 3340
rect 37568 2854 37596 3334
rect 37556 2848 37608 2854
rect 37556 2790 37608 2796
rect 37568 2650 37596 2790
rect 37936 2774 37964 5238
rect 38120 4078 38148 5850
rect 38200 5228 38252 5234
rect 38200 5170 38252 5176
rect 38212 4865 38240 5170
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38108 4072 38160 4078
rect 38108 4014 38160 4020
rect 38200 3936 38252 3942
rect 38200 3878 38252 3884
rect 37936 2746 38056 2774
rect 37556 2644 37608 2650
rect 37556 2586 37608 2592
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35716 2440 35768 2446
rect 35716 2382 35768 2388
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 34428 2372 34480 2378
rect 34428 2314 34480 2320
rect 35452 800 35480 2382
rect 35716 2304 35768 2310
rect 35716 2246 35768 2252
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 35728 2106 35756 2246
rect 35716 2100 35768 2106
rect 35716 2042 35768 2048
rect 37200 1465 37228 2246
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37384 800 37412 2246
rect 38028 1970 38056 2746
rect 38212 2650 38240 3878
rect 38304 3534 38332 9318
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 38292 2848 38344 2854
rect 38290 2816 38292 2825
rect 38344 2816 38346 2825
rect 38290 2751 38346 2760
rect 38200 2644 38252 2650
rect 38200 2586 38252 2592
rect 38016 1964 38068 1970
rect 38016 1906 38068 1912
rect 39316 800 39344 3470
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21914 200 21970 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
rect 39302 200 39358 800
<< via2 >>
rect 2962 39480 3018 39536
rect 2870 37440 2926 37496
rect 1674 36080 1730 36136
rect 1674 34040 1730 34096
rect 1582 32020 1638 32056
rect 1582 32000 1584 32020
rect 1584 32000 1636 32020
rect 1636 32000 1638 32020
rect 1674 30660 1730 30696
rect 1674 30640 1676 30660
rect 1676 30640 1728 30660
rect 1728 30640 1730 30660
rect 1582 28636 1584 28656
rect 1584 28636 1636 28656
rect 1636 28636 1638 28656
rect 1582 28600 1638 28636
rect 1674 26560 1730 26616
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1674 23160 1730 23216
rect 1674 21120 1730 21176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1674 19760 1730 19816
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 1674 15680 1730 15736
rect 1674 14320 1730 14376
rect 1674 12280 1730 12336
rect 1582 10260 1638 10296
rect 1582 10240 1584 10260
rect 1584 10240 1636 10260
rect 1636 10240 1638 10260
rect 1582 8916 1584 8936
rect 1584 8916 1636 8936
rect 1636 8916 1638 8936
rect 1582 8880 1638 8916
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1582 6840 1638 6896
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1674 4800 1730 4856
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1582 3476 1584 3496
rect 1584 3476 1636 3496
rect 1636 3476 1638 3496
rect 1582 3440 1638 3476
rect 1766 3440 1822 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 13174 13796 13230 13832
rect 13174 13776 13176 13796
rect 13176 13776 13228 13796
rect 13228 13776 13230 13796
rect 12898 12416 12954 12472
rect 10414 4392 10470 4448
rect 13174 5888 13230 5944
rect 14278 13948 14280 13968
rect 14280 13948 14332 13968
rect 14332 13948 14334 13968
rect 14278 13912 14334 13948
rect 13818 8880 13874 8936
rect 13634 8064 13690 8120
rect 13910 8200 13966 8256
rect 13818 6976 13874 7032
rect 14278 8472 14334 8528
rect 15566 14068 15622 14104
rect 15566 14048 15568 14068
rect 15568 14048 15620 14068
rect 15620 14048 15622 14068
rect 16578 15020 16634 15056
rect 16578 15000 16580 15020
rect 16580 15000 16632 15020
rect 16632 15000 16634 15020
rect 16302 13812 16304 13832
rect 16304 13812 16356 13832
rect 16356 13812 16358 13832
rect 16302 13776 16358 13812
rect 16394 13368 16450 13424
rect 15566 11192 15622 11248
rect 14094 3984 14150 4040
rect 15382 10124 15438 10160
rect 15382 10104 15384 10124
rect 15384 10104 15436 10124
rect 15436 10104 15438 10124
rect 15382 9560 15438 9616
rect 15290 7928 15346 7984
rect 14830 7112 14886 7168
rect 15198 5752 15254 5808
rect 14922 5516 14924 5536
rect 14924 5516 14976 5536
rect 14976 5516 14978 5536
rect 14922 5480 14978 5516
rect 15750 9152 15806 9208
rect 16302 11872 16358 11928
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 16854 14048 16910 14104
rect 16854 13524 16910 13560
rect 16854 13504 16856 13524
rect 16856 13504 16908 13524
rect 16908 13504 16910 13524
rect 16210 9968 16266 10024
rect 16578 10512 16634 10568
rect 16578 8780 16580 8800
rect 16580 8780 16632 8800
rect 16632 8780 16634 8800
rect 16578 8744 16634 8780
rect 16026 5072 16082 5128
rect 16210 5636 16266 5672
rect 16210 5616 16212 5636
rect 16212 5616 16264 5636
rect 16264 5616 16266 5636
rect 16118 4800 16174 4856
rect 15934 4528 15990 4584
rect 16302 4392 16358 4448
rect 15750 3168 15806 3224
rect 1674 1400 1730 1456
rect 16578 7248 16634 7304
rect 17866 16496 17922 16552
rect 17038 13932 17094 13968
rect 17038 13912 17040 13932
rect 17040 13912 17092 13932
rect 17092 13912 17094 13932
rect 17038 12144 17094 12200
rect 17590 13640 17646 13696
rect 17682 12552 17738 12608
rect 17314 12280 17370 12336
rect 17406 11772 17408 11792
rect 17408 11772 17460 11792
rect 17460 11772 17462 11792
rect 17406 11736 17462 11772
rect 17314 9152 17370 9208
rect 17222 8628 17278 8664
rect 17222 8608 17224 8628
rect 17224 8608 17276 8628
rect 17276 8608 17278 8628
rect 17406 7792 17462 7848
rect 17038 6724 17094 6760
rect 17038 6704 17040 6724
rect 17040 6704 17092 6724
rect 17092 6704 17094 6724
rect 16578 4936 16634 4992
rect 16946 5364 17002 5400
rect 16946 5344 16948 5364
rect 16948 5344 17000 5364
rect 17000 5344 17002 5364
rect 17222 6840 17278 6896
rect 16854 4684 16910 4720
rect 16854 4664 16856 4684
rect 16856 4664 16908 4684
rect 16908 4664 16910 4684
rect 17774 10668 17830 10704
rect 17774 10648 17776 10668
rect 17776 10648 17828 10668
rect 17828 10648 17830 10668
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18326 15000 18382 15056
rect 17958 10104 18014 10160
rect 17314 4684 17370 4720
rect 17314 4664 17316 4684
rect 17316 4664 17368 4684
rect 17368 4664 17370 4684
rect 17314 4428 17316 4448
rect 17316 4428 17368 4448
rect 17368 4428 17370 4448
rect 17314 4392 17370 4428
rect 18326 11092 18328 11112
rect 18328 11092 18380 11112
rect 18380 11092 18382 11112
rect 18326 11056 18382 11092
rect 18326 8608 18382 8664
rect 18510 13776 18566 13832
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 18510 8744 18566 8800
rect 17866 4664 17922 4720
rect 17958 3984 18014 4040
rect 18878 8200 18934 8256
rect 18878 8064 18934 8120
rect 19614 14592 19670 14648
rect 20074 14592 20130 14648
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19154 11872 19210 11928
rect 19246 11736 19302 11792
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19522 12860 19524 12880
rect 19524 12860 19576 12880
rect 19576 12860 19578 12880
rect 19522 12824 19578 12860
rect 21086 17620 21088 17640
rect 21088 17620 21140 17640
rect 21140 17620 21142 17640
rect 21086 17584 21142 17620
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19522 11328 19578 11384
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19338 8064 19394 8120
rect 18786 5516 18788 5536
rect 18788 5516 18840 5536
rect 18840 5516 18842 5536
rect 18786 5480 18842 5516
rect 18786 5092 18842 5128
rect 18786 5072 18788 5092
rect 18788 5072 18840 5092
rect 18840 5072 18842 5092
rect 18694 4972 18696 4992
rect 18696 4972 18748 4992
rect 18748 4972 18750 4992
rect 18694 4936 18750 4972
rect 18694 4820 18750 4856
rect 18694 4800 18696 4820
rect 18696 4800 18748 4820
rect 18748 4800 18750 4820
rect 18786 3168 18842 3224
rect 19338 7520 19394 7576
rect 19154 6296 19210 6352
rect 19154 5888 19210 5944
rect 19154 5344 19210 5400
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19614 7384 19670 7440
rect 19890 7384 19946 7440
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20810 13232 20866 13288
rect 20626 11736 20682 11792
rect 21454 15564 21510 15600
rect 21454 15544 21456 15564
rect 21456 15544 21508 15564
rect 21508 15544 21510 15564
rect 21822 17584 21878 17640
rect 21822 14728 21878 14784
rect 21638 13912 21694 13968
rect 21178 13232 21234 13288
rect 20810 12280 20866 12336
rect 21086 11056 21142 11112
rect 20626 10376 20682 10432
rect 20534 10240 20590 10296
rect 20258 7384 20314 7440
rect 21362 11500 21364 11520
rect 21364 11500 21416 11520
rect 21416 11500 21418 11520
rect 21362 11464 21418 11500
rect 21822 12552 21878 12608
rect 21362 10376 21418 10432
rect 20258 6160 20314 6216
rect 20166 6024 20222 6080
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19338 4936 19394 4992
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19430 2796 19432 2816
rect 19432 2796 19484 2816
rect 19484 2796 19486 2816
rect 19430 2760 19486 2796
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21546 8064 21602 8120
rect 21454 7792 21510 7848
rect 20810 5244 20812 5264
rect 20812 5244 20864 5264
rect 20864 5244 20866 5264
rect 20810 5208 20866 5244
rect 20994 3168 21050 3224
rect 22466 15544 22522 15600
rect 22006 13368 22062 13424
rect 22190 13776 22246 13832
rect 22374 14048 22430 14104
rect 22190 11192 22246 11248
rect 22098 11056 22154 11112
rect 22098 10956 22100 10976
rect 22100 10956 22152 10976
rect 22152 10956 22154 10976
rect 22098 10920 22154 10956
rect 22098 10804 22154 10840
rect 22098 10784 22100 10804
rect 22100 10784 22152 10804
rect 22152 10784 22154 10804
rect 22834 15544 22890 15600
rect 22926 14048 22982 14104
rect 22466 9716 22522 9752
rect 22466 9696 22468 9716
rect 22468 9696 22520 9716
rect 22520 9696 22522 9716
rect 22098 9172 22154 9208
rect 22098 9152 22100 9172
rect 22100 9152 22152 9172
rect 22152 9152 22154 9172
rect 22098 7656 22154 7712
rect 22006 7112 22062 7168
rect 21730 6840 21786 6896
rect 21546 6568 21602 6624
rect 21178 5072 21234 5128
rect 21362 5344 21418 5400
rect 22282 6296 22338 6352
rect 22650 11056 22706 11112
rect 22742 10512 22798 10568
rect 23018 13640 23074 13696
rect 23846 16124 23848 16144
rect 23848 16124 23900 16144
rect 23900 16124 23902 16144
rect 23846 16088 23902 16124
rect 23018 11600 23074 11656
rect 23478 13504 23534 13560
rect 23754 13912 23810 13968
rect 21914 4820 21970 4856
rect 21914 4800 21916 4820
rect 21916 4800 21968 4820
rect 21968 4800 21970 4820
rect 22098 4820 22154 4856
rect 22098 4800 22100 4820
rect 22100 4800 22152 4820
rect 22152 4800 22154 4820
rect 22098 4276 22154 4312
rect 22098 4256 22100 4276
rect 22100 4256 22152 4276
rect 22152 4256 22154 4276
rect 21454 3984 21510 4040
rect 21914 3732 21970 3768
rect 21914 3712 21916 3732
rect 21916 3712 21968 3732
rect 21968 3712 21970 3732
rect 21638 3596 21694 3632
rect 21638 3576 21640 3596
rect 21640 3576 21692 3596
rect 21692 3576 21694 3596
rect 22190 2760 22246 2816
rect 22742 7692 22744 7712
rect 22744 7692 22796 7712
rect 22796 7692 22798 7712
rect 22742 7656 22798 7692
rect 23202 9152 23258 9208
rect 23478 10804 23534 10840
rect 23478 10784 23480 10804
rect 23480 10784 23532 10804
rect 23532 10784 23534 10804
rect 23386 10376 23442 10432
rect 23754 12280 23810 12336
rect 24030 11736 24086 11792
rect 23938 10240 23994 10296
rect 24214 10920 24270 10976
rect 24858 16496 24914 16552
rect 24582 14048 24638 14104
rect 24398 11464 24454 11520
rect 25134 14456 25190 14512
rect 25410 16496 25466 16552
rect 24582 12416 24638 12472
rect 24582 11328 24638 11384
rect 25134 12008 25190 12064
rect 24674 10920 24730 10976
rect 25226 11736 25282 11792
rect 24858 9988 24914 10024
rect 24858 9968 24860 9988
rect 24860 9968 24912 9988
rect 24912 9968 24914 9988
rect 24858 8900 24914 8936
rect 24858 8880 24860 8900
rect 24860 8880 24912 8900
rect 24912 8880 24914 8900
rect 25042 8508 25044 8528
rect 25044 8508 25096 8528
rect 25096 8508 25098 8528
rect 25042 8472 25098 8508
rect 23938 6568 23994 6624
rect 23846 5072 23902 5128
rect 23570 3712 23626 3768
rect 23478 3576 23534 3632
rect 24030 5344 24086 5400
rect 24490 7520 24546 7576
rect 24858 6704 24914 6760
rect 24582 6196 24584 6216
rect 24584 6196 24636 6216
rect 24636 6196 24638 6216
rect 24582 6160 24638 6196
rect 24398 4936 24454 4992
rect 25318 5752 25374 5808
rect 25318 5208 25374 5264
rect 24766 4664 24822 4720
rect 24950 4564 24952 4584
rect 24952 4564 25004 4584
rect 25004 4564 25006 4584
rect 24950 4528 25006 4564
rect 25134 4276 25190 4312
rect 25134 4256 25136 4276
rect 25136 4256 25188 4276
rect 25188 4256 25190 4276
rect 25778 15444 25780 15464
rect 25780 15444 25832 15464
rect 25832 15444 25834 15464
rect 25778 15408 25834 15444
rect 25594 15000 25650 15056
rect 25686 14592 25742 14648
rect 25778 14320 25834 14376
rect 25594 12860 25596 12880
rect 25596 12860 25648 12880
rect 25648 12860 25650 12880
rect 25594 12824 25650 12860
rect 26146 15000 26202 15056
rect 26146 13912 26202 13968
rect 25962 12144 26018 12200
rect 26054 10956 26056 10976
rect 26056 10956 26108 10976
rect 26108 10956 26110 10976
rect 26054 10920 26110 10956
rect 26330 14184 26386 14240
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38800 37242 38856
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 28354 17620 28356 17640
rect 28356 17620 28408 17640
rect 28408 17620 28410 17640
rect 28354 17584 28410 17620
rect 27986 14592 28042 14648
rect 28446 14456 28502 14512
rect 28078 14184 28134 14240
rect 27618 12164 27674 12200
rect 27618 12144 27620 12164
rect 27620 12144 27672 12164
rect 27672 12144 27674 12164
rect 27710 12044 27712 12064
rect 27712 12044 27764 12064
rect 27764 12044 27766 12064
rect 27710 12008 27766 12044
rect 27802 11736 27858 11792
rect 27710 11464 27766 11520
rect 28630 14592 28686 14648
rect 28538 13504 28594 13560
rect 28354 11600 28410 11656
rect 27618 9596 27620 9616
rect 27620 9596 27672 9616
rect 27672 9596 27674 9616
rect 27618 9560 27674 9596
rect 28814 14048 28870 14104
rect 28998 14864 29054 14920
rect 29090 14320 29146 14376
rect 29090 10648 29146 10704
rect 28446 9696 28502 9752
rect 28538 6976 28594 7032
rect 28262 6160 28318 6216
rect 26606 3984 26662 4040
rect 26238 3440 26294 3496
rect 25778 3168 25834 3224
rect 28998 7248 29054 7304
rect 29734 12280 29790 12336
rect 29642 11736 29698 11792
rect 28906 6024 28962 6080
rect 29550 8608 29606 8664
rect 29550 8356 29606 8392
rect 29550 8336 29552 8356
rect 29552 8336 29604 8356
rect 29604 8336 29606 8356
rect 30470 14068 30526 14104
rect 30470 14048 30472 14068
rect 30472 14048 30524 14068
rect 30524 14048 30526 14068
rect 30378 11328 30434 11384
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 32034 16088 32090 16144
rect 31114 13524 31170 13560
rect 31114 13504 31116 13524
rect 31116 13504 31168 13524
rect 31168 13504 31170 13524
rect 30930 11756 30986 11792
rect 30930 11736 30932 11756
rect 30932 11736 30984 11756
rect 30984 11736 30986 11756
rect 30470 5616 30526 5672
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38290 37440 38346 37496
rect 37462 35400 37518 35456
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38290 32020 38346 32056
rect 38290 32000 38292 32020
rect 38292 32000 38344 32020
rect 38344 32000 38346 32020
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38198 27940 38254 27976
rect 38198 27920 38200 27940
rect 38200 27920 38252 27940
rect 38252 27920 38254 27940
rect 38198 26560 38254 26616
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21120 38254 21176
rect 38198 19116 38200 19136
rect 38200 19116 38252 19136
rect 38252 19116 38254 19136
rect 38198 19080 38254 19116
rect 38198 17040 38254 17096
rect 33046 8608 33102 8664
rect 32218 6976 32274 7032
rect 32678 6976 32734 7032
rect 31758 3188 31814 3224
rect 31758 3168 31760 3188
rect 31760 3168 31812 3188
rect 31812 3168 31814 3188
rect 31298 2932 31300 2952
rect 31300 2932 31352 2952
rect 31352 2932 31354 2952
rect 31298 2896 31354 2932
rect 31758 2916 31814 2952
rect 31758 2896 31760 2916
rect 31760 2896 31812 2916
rect 31812 2896 31814 2916
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35990 8336 36046 8392
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 33690 3168 33746 3224
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36634 7948 36690 7984
rect 36634 7928 36636 7948
rect 36636 7928 36688 7948
rect 36688 7928 36690 7948
rect 37186 8200 37242 8256
rect 38198 15680 38254 15736
rect 38290 13640 38346 13696
rect 38198 11600 38254 11656
rect 38290 10240 38346 10296
rect 38198 6160 38254 6216
rect 38198 4800 38254 4856
rect 37186 1400 37242 1456
rect 38290 2796 38292 2816
rect 38292 2796 38344 2816
rect 38344 2796 38346 2816
rect 38290 2760 38346 2796
<< metal3 >>
rect 200 39538 800 39568
rect 2957 39538 3023 39541
rect 200 39536 3023 39538
rect 200 39480 2962 39536
rect 3018 39480 3023 39536
rect 200 39478 3023 39480
rect 200 39448 800 39478
rect 2957 39475 3023 39478
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 2865 37498 2931 37501
rect 200 37496 2931 37498
rect 200 37440 2870 37496
rect 2926 37440 2931 37496
rect 200 37438 2931 37440
rect 200 37408 800 37438
rect 2865 37435 2931 37438
rect 38285 37498 38351 37501
rect 39200 37498 39800 37528
rect 38285 37496 39800 37498
rect 38285 37440 38290 37496
rect 38346 37440 39800 37496
rect 38285 37438 39800 37440
rect 38285 37435 38351 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 36048 800 36078
rect 1669 36075 1735 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 37457 35458 37523 35461
rect 39200 35458 39800 35488
rect 37457 35456 39800 35458
rect 37457 35400 37462 35456
rect 37518 35400 39800 35456
rect 37457 35398 39800 35400
rect 37457 35395 37523 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1669 34098 1735 34101
rect 200 34096 1735 34098
rect 200 34040 1674 34096
rect 1730 34040 1735 34096
rect 200 34038 1735 34040
rect 200 34008 800 34038
rect 1669 34035 1735 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31968 800 31998
rect 1577 31995 1643 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1577 28658 1643 28661
rect 200 28656 1643 28658
rect 200 28600 1582 28656
rect 1638 28600 1643 28656
rect 200 28598 1643 28600
rect 200 28568 800 28598
rect 1577 28595 1643 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 38193 27978 38259 27981
rect 39200 27978 39800 28008
rect 38193 27976 39800 27978
rect 38193 27920 38198 27976
rect 38254 27920 39800 27976
rect 38193 27918 39800 27920
rect 38193 27915 38259 27918
rect 39200 27888 39800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 38193 26618 38259 26621
rect 39200 26618 39800 26648
rect 38193 26616 39800 26618
rect 38193 26560 38198 26616
rect 38254 26560 39800 26616
rect 38193 26558 39800 26560
rect 38193 26555 38259 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25168 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1669 23218 1735 23221
rect 200 23216 1735 23218
rect 200 23160 1674 23216
rect 1730 23160 1735 23216
rect 200 23158 1735 23160
rect 200 23128 800 23158
rect 1669 23155 1735 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1669 19818 1735 19821
rect 200 19816 1735 19818
rect 200 19760 1674 19816
rect 1730 19760 1735 19816
rect 200 19758 1735 19760
rect 200 19728 800 19758
rect 1669 19755 1735 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1577 17778 1643 17781
rect 200 17776 1643 17778
rect 200 17720 1582 17776
rect 1638 17720 1643 17776
rect 200 17718 1643 17720
rect 200 17688 800 17718
rect 1577 17715 1643 17718
rect 21081 17642 21147 17645
rect 21817 17642 21883 17645
rect 28349 17642 28415 17645
rect 21081 17640 28415 17642
rect 21081 17584 21086 17640
rect 21142 17584 21822 17640
rect 21878 17584 28354 17640
rect 28410 17584 28415 17640
rect 21081 17582 28415 17584
rect 21081 17579 21147 17582
rect 21817 17579 21883 17582
rect 28349 17579 28415 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 17861 16554 17927 16557
rect 24853 16554 24919 16557
rect 25405 16554 25471 16557
rect 17861 16552 25471 16554
rect 17861 16496 17866 16552
rect 17922 16496 24858 16552
rect 24914 16496 25410 16552
rect 25466 16496 25471 16552
rect 17861 16494 25471 16496
rect 17861 16491 17927 16494
rect 24853 16491 24919 16494
rect 25405 16491 25471 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 23841 16146 23907 16149
rect 32029 16146 32095 16149
rect 23841 16144 32095 16146
rect 23841 16088 23846 16144
rect 23902 16088 32034 16144
rect 32090 16088 32095 16144
rect 23841 16086 32095 16088
rect 23841 16083 23907 16086
rect 32029 16083 32095 16086
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 21449 15602 21515 15605
rect 22461 15602 22527 15605
rect 22829 15602 22895 15605
rect 21449 15600 22895 15602
rect 21449 15544 21454 15600
rect 21510 15544 22466 15600
rect 22522 15544 22834 15600
rect 22890 15544 22895 15600
rect 21449 15542 22895 15544
rect 21449 15539 21515 15542
rect 22461 15539 22527 15542
rect 22829 15539 22895 15542
rect 24710 15404 24716 15468
rect 24780 15466 24786 15468
rect 25773 15466 25839 15469
rect 24780 15464 25839 15466
rect 24780 15408 25778 15464
rect 25834 15408 25839 15464
rect 24780 15406 25839 15408
rect 24780 15404 24786 15406
rect 25773 15403 25839 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 16573 15058 16639 15061
rect 18321 15058 18387 15061
rect 25589 15058 25655 15061
rect 16573 15056 18387 15058
rect 16573 15000 16578 15056
rect 16634 15000 18326 15056
rect 18382 15000 18387 15056
rect 16573 14998 18387 15000
rect 16573 14995 16639 14998
rect 18321 14995 18387 14998
rect 22050 15056 25655 15058
rect 22050 15000 25594 15056
rect 25650 15000 25655 15056
rect 22050 14998 25655 15000
rect 21817 14786 21883 14789
rect 22050 14786 22110 14998
rect 25589 14995 25655 14998
rect 26141 15060 26207 15061
rect 26141 15056 26188 15060
rect 26252 15058 26258 15060
rect 26141 15000 26146 15056
rect 26141 14996 26188 15000
rect 26252 14998 26298 15058
rect 26252 14996 26258 14998
rect 26141 14995 26207 14996
rect 28993 14922 29059 14925
rect 28950 14920 29059 14922
rect 28950 14864 28998 14920
rect 29054 14864 29059 14920
rect 28950 14859 29059 14864
rect 28950 14786 29010 14859
rect 21817 14784 22110 14786
rect 21817 14728 21822 14784
rect 21878 14728 22110 14784
rect 21817 14726 22110 14728
rect 22188 14726 29010 14786
rect 21817 14723 21883 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 19609 14650 19675 14653
rect 20069 14650 20135 14653
rect 22188 14650 22248 14726
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19609 14648 22248 14650
rect 19609 14592 19614 14648
rect 19670 14592 20074 14648
rect 20130 14592 22248 14648
rect 19609 14590 22248 14592
rect 25681 14650 25747 14653
rect 27981 14650 28047 14653
rect 28625 14650 28691 14653
rect 25681 14648 28691 14650
rect 25681 14592 25686 14648
rect 25742 14592 27986 14648
rect 28042 14592 28630 14648
rect 28686 14592 28691 14648
rect 25681 14590 28691 14592
rect 19609 14587 19675 14590
rect 20069 14587 20135 14590
rect 25681 14587 25747 14590
rect 27981 14587 28047 14590
rect 28625 14587 28691 14590
rect 25129 14514 25195 14517
rect 28441 14514 28507 14517
rect 25129 14512 28507 14514
rect 25129 14456 25134 14512
rect 25190 14456 28446 14512
rect 28502 14456 28507 14512
rect 25129 14454 28507 14456
rect 25129 14451 25195 14454
rect 28441 14451 28507 14454
rect 200 14378 800 14408
rect 1669 14378 1735 14381
rect 200 14376 1735 14378
rect 200 14320 1674 14376
rect 1730 14320 1735 14376
rect 200 14318 1735 14320
rect 200 14288 800 14318
rect 1669 14315 1735 14318
rect 25773 14378 25839 14381
rect 29085 14378 29151 14381
rect 25773 14376 29151 14378
rect 25773 14320 25778 14376
rect 25834 14320 29090 14376
rect 29146 14320 29151 14376
rect 25773 14318 29151 14320
rect 25773 14315 25839 14318
rect 29085 14315 29151 14318
rect 26325 14242 26391 14245
rect 28073 14242 28139 14245
rect 26325 14240 28139 14242
rect 26325 14184 26330 14240
rect 26386 14184 28078 14240
rect 28134 14184 28139 14240
rect 26325 14182 28139 14184
rect 26325 14179 26391 14182
rect 28073 14179 28139 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 15561 14106 15627 14109
rect 16849 14106 16915 14109
rect 15561 14104 16915 14106
rect 15561 14048 15566 14104
rect 15622 14048 16854 14104
rect 16910 14048 16915 14104
rect 15561 14046 16915 14048
rect 15561 14043 15627 14046
rect 16849 14043 16915 14046
rect 22369 14106 22435 14109
rect 22921 14106 22987 14109
rect 24577 14106 24643 14109
rect 28809 14106 28875 14109
rect 30465 14106 30531 14109
rect 22369 14104 30531 14106
rect 22369 14048 22374 14104
rect 22430 14048 22926 14104
rect 22982 14048 24582 14104
rect 24638 14048 28814 14104
rect 28870 14048 30470 14104
rect 30526 14048 30531 14104
rect 22369 14046 30531 14048
rect 22369 14043 22435 14046
rect 22921 14043 22987 14046
rect 24577 14043 24643 14046
rect 28809 14043 28875 14046
rect 30465 14043 30531 14046
rect 14273 13970 14339 13973
rect 17033 13970 17099 13973
rect 14273 13968 17099 13970
rect 14273 13912 14278 13968
rect 14334 13912 17038 13968
rect 17094 13912 17099 13968
rect 14273 13910 17099 13912
rect 14273 13907 14339 13910
rect 17033 13907 17099 13910
rect 21633 13970 21699 13973
rect 23749 13970 23815 13973
rect 26141 13972 26207 13973
rect 26141 13970 26188 13972
rect 21633 13968 23815 13970
rect 21633 13912 21638 13968
rect 21694 13912 23754 13968
rect 23810 13912 23815 13968
rect 21633 13910 23815 13912
rect 26096 13968 26188 13970
rect 26096 13912 26146 13968
rect 26096 13910 26188 13912
rect 21633 13907 21699 13910
rect 23749 13907 23815 13910
rect 26141 13908 26188 13910
rect 26252 13908 26258 13972
rect 26141 13907 26207 13908
rect 13169 13834 13235 13837
rect 16297 13834 16363 13837
rect 13169 13832 16363 13834
rect 13169 13776 13174 13832
rect 13230 13776 16302 13832
rect 16358 13776 16363 13832
rect 13169 13774 16363 13776
rect 13169 13771 13235 13774
rect 16297 13771 16363 13774
rect 18505 13834 18571 13837
rect 22185 13834 22251 13837
rect 18505 13832 22251 13834
rect 18505 13776 18510 13832
rect 18566 13776 22190 13832
rect 22246 13776 22251 13832
rect 18505 13774 22251 13776
rect 18505 13771 18571 13774
rect 22185 13771 22251 13774
rect 17585 13698 17651 13701
rect 23013 13698 23079 13701
rect 17585 13696 23079 13698
rect 17585 13640 17590 13696
rect 17646 13640 23018 13696
rect 23074 13640 23079 13696
rect 17585 13638 23079 13640
rect 17585 13635 17651 13638
rect 23013 13635 23079 13638
rect 38285 13698 38351 13701
rect 39200 13698 39800 13728
rect 38285 13696 39800 13698
rect 38285 13640 38290 13696
rect 38346 13640 39800 13696
rect 38285 13638 39800 13640
rect 38285 13635 38351 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 16849 13562 16915 13565
rect 23473 13562 23539 13565
rect 16849 13560 23539 13562
rect 16849 13504 16854 13560
rect 16910 13504 23478 13560
rect 23534 13504 23539 13560
rect 16849 13502 23539 13504
rect 16849 13499 16915 13502
rect 23473 13499 23539 13502
rect 28533 13562 28599 13565
rect 31109 13562 31175 13565
rect 28533 13560 31175 13562
rect 28533 13504 28538 13560
rect 28594 13504 31114 13560
rect 31170 13504 31175 13560
rect 28533 13502 31175 13504
rect 28533 13499 28599 13502
rect 31109 13499 31175 13502
rect 16389 13426 16455 13429
rect 22001 13426 22067 13429
rect 16389 13424 22067 13426
rect 16389 13368 16394 13424
rect 16450 13368 22006 13424
rect 22062 13368 22067 13424
rect 16389 13366 22067 13368
rect 16389 13363 16455 13366
rect 22001 13363 22067 13366
rect 20805 13290 20871 13293
rect 21173 13290 21239 13293
rect 20805 13288 21239 13290
rect 20805 13232 20810 13288
rect 20866 13232 21178 13288
rect 21234 13232 21239 13288
rect 20805 13230 21239 13232
rect 20805 13227 20871 13230
rect 21173 13227 21239 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 19517 12882 19583 12885
rect 25589 12882 25655 12885
rect 19517 12880 25655 12882
rect 19517 12824 19522 12880
rect 19578 12824 25594 12880
rect 25650 12824 25655 12880
rect 19517 12822 25655 12824
rect 19517 12819 19583 12822
rect 25589 12819 25655 12822
rect 17677 12610 17743 12613
rect 21817 12610 21883 12613
rect 17677 12608 21883 12610
rect 17677 12552 17682 12608
rect 17738 12552 21822 12608
rect 21878 12552 21883 12608
rect 17677 12550 21883 12552
rect 17677 12547 17743 12550
rect 21817 12547 21883 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 12893 12474 12959 12477
rect 24577 12474 24643 12477
rect 12893 12472 24643 12474
rect 12893 12416 12898 12472
rect 12954 12416 24582 12472
rect 24638 12416 24643 12472
rect 12893 12414 24643 12416
rect 12893 12411 12959 12414
rect 24577 12411 24643 12414
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 17309 12338 17375 12341
rect 20805 12338 20871 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 17174 12336 20871 12338
rect 17174 12280 17314 12336
rect 17370 12280 20810 12336
rect 20866 12280 20871 12336
rect 17174 12278 20871 12280
rect 17033 12202 17099 12205
rect 17174 12202 17234 12278
rect 17309 12275 17375 12278
rect 20805 12275 20871 12278
rect 23749 12338 23815 12341
rect 29729 12338 29795 12341
rect 23749 12336 29795 12338
rect 23749 12280 23754 12336
rect 23810 12280 29734 12336
rect 29790 12280 29795 12336
rect 23749 12278 29795 12280
rect 23749 12275 23815 12278
rect 29729 12275 29795 12278
rect 17033 12200 17234 12202
rect 17033 12144 17038 12200
rect 17094 12144 17234 12200
rect 17033 12142 17234 12144
rect 25957 12202 26023 12205
rect 27613 12202 27679 12205
rect 25957 12200 27679 12202
rect 25957 12144 25962 12200
rect 26018 12144 27618 12200
rect 27674 12144 27679 12200
rect 25957 12142 27679 12144
rect 17033 12139 17099 12142
rect 25957 12139 26023 12142
rect 27613 12139 27679 12142
rect 25129 12066 25195 12069
rect 27705 12066 27771 12069
rect 25129 12064 27771 12066
rect 25129 12008 25134 12064
rect 25190 12008 27710 12064
rect 27766 12008 27771 12064
rect 25129 12006 27771 12008
rect 25129 12003 25195 12006
rect 27705 12003 27771 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 16297 11930 16363 11933
rect 19149 11930 19215 11933
rect 16297 11928 19215 11930
rect 16297 11872 16302 11928
rect 16358 11872 19154 11928
rect 19210 11872 19215 11928
rect 16297 11870 19215 11872
rect 16297 11867 16363 11870
rect 19149 11867 19215 11870
rect 17401 11794 17467 11797
rect 19241 11794 19307 11797
rect 17401 11792 19307 11794
rect 17401 11736 17406 11792
rect 17462 11736 19246 11792
rect 19302 11736 19307 11792
rect 17401 11734 19307 11736
rect 17401 11731 17467 11734
rect 19241 11731 19307 11734
rect 20621 11794 20687 11797
rect 24025 11794 24091 11797
rect 20621 11792 24091 11794
rect 20621 11736 20626 11792
rect 20682 11736 24030 11792
rect 24086 11736 24091 11792
rect 20621 11734 24091 11736
rect 20621 11731 20687 11734
rect 24025 11731 24091 11734
rect 25221 11794 25287 11797
rect 27797 11794 27863 11797
rect 25221 11792 27863 11794
rect 25221 11736 25226 11792
rect 25282 11736 27802 11792
rect 27858 11736 27863 11792
rect 25221 11734 27863 11736
rect 25221 11731 25287 11734
rect 27797 11731 27863 11734
rect 29637 11794 29703 11797
rect 30925 11794 30991 11797
rect 29637 11792 30991 11794
rect 29637 11736 29642 11792
rect 29698 11736 30930 11792
rect 30986 11736 30991 11792
rect 29637 11734 30991 11736
rect 29637 11731 29703 11734
rect 30925 11731 30991 11734
rect 23013 11658 23079 11661
rect 28349 11658 28415 11661
rect 23013 11656 28415 11658
rect 23013 11600 23018 11656
rect 23074 11600 28354 11656
rect 28410 11600 28415 11656
rect 23013 11598 28415 11600
rect 23013 11595 23079 11598
rect 28349 11595 28415 11598
rect 38193 11658 38259 11661
rect 39200 11658 39800 11688
rect 38193 11656 39800 11658
rect 38193 11600 38198 11656
rect 38254 11600 39800 11656
rect 38193 11598 39800 11600
rect 38193 11595 38259 11598
rect 39200 11568 39800 11598
rect 21357 11522 21423 11525
rect 24393 11522 24459 11525
rect 27705 11522 27771 11525
rect 21357 11520 29010 11522
rect 21357 11464 21362 11520
rect 21418 11464 24398 11520
rect 24454 11464 27710 11520
rect 27766 11464 29010 11520
rect 21357 11462 29010 11464
rect 21357 11459 21423 11462
rect 24393 11459 24459 11462
rect 27705 11459 27771 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 19517 11386 19583 11389
rect 24577 11386 24643 11389
rect 19517 11384 24643 11386
rect 19517 11328 19522 11384
rect 19578 11328 24582 11384
rect 24638 11328 24643 11384
rect 19517 11326 24643 11328
rect 28950 11386 29010 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 30373 11386 30439 11389
rect 28950 11384 30439 11386
rect 28950 11328 30378 11384
rect 30434 11328 30439 11384
rect 28950 11326 30439 11328
rect 19517 11323 19583 11326
rect 24577 11323 24643 11326
rect 30373 11323 30439 11326
rect 15561 11250 15627 11253
rect 22185 11250 22251 11253
rect 15561 11248 22251 11250
rect 15561 11192 15566 11248
rect 15622 11192 22190 11248
rect 22246 11192 22251 11248
rect 15561 11190 22251 11192
rect 15561 11187 15627 11190
rect 22185 11187 22251 11190
rect 18321 11114 18387 11117
rect 21081 11114 21147 11117
rect 18321 11112 21147 11114
rect 18321 11056 18326 11112
rect 18382 11056 21086 11112
rect 21142 11056 21147 11112
rect 18321 11054 21147 11056
rect 18321 11051 18387 11054
rect 21081 11051 21147 11054
rect 22093 11114 22159 11117
rect 22645 11114 22711 11117
rect 22093 11112 22711 11114
rect 22093 11056 22098 11112
rect 22154 11056 22650 11112
rect 22706 11056 22711 11112
rect 22093 11054 22711 11056
rect 22093 11051 22159 11054
rect 22645 11051 22711 11054
rect 22093 10978 22159 10981
rect 24209 10978 24275 10981
rect 22093 10976 24275 10978
rect 22093 10920 22098 10976
rect 22154 10920 24214 10976
rect 24270 10920 24275 10976
rect 22093 10918 24275 10920
rect 22093 10915 22159 10918
rect 24209 10915 24275 10918
rect 24669 10978 24735 10981
rect 26049 10978 26115 10981
rect 24669 10976 26115 10978
rect 24669 10920 24674 10976
rect 24730 10920 26054 10976
rect 26110 10920 26115 10976
rect 24669 10918 26115 10920
rect 24669 10915 24735 10918
rect 26049 10915 26115 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 22093 10842 22159 10845
rect 23473 10842 23539 10845
rect 22093 10840 23539 10842
rect 22093 10784 22098 10840
rect 22154 10784 23478 10840
rect 23534 10784 23539 10840
rect 22093 10782 23539 10784
rect 22093 10779 22159 10782
rect 23473 10779 23539 10782
rect 17769 10706 17835 10709
rect 29085 10706 29151 10709
rect 17769 10704 29151 10706
rect 17769 10648 17774 10704
rect 17830 10648 29090 10704
rect 29146 10648 29151 10704
rect 17769 10646 29151 10648
rect 17769 10643 17835 10646
rect 29085 10643 29151 10646
rect 16573 10570 16639 10573
rect 22737 10570 22803 10573
rect 16573 10568 22803 10570
rect 16573 10512 16578 10568
rect 16634 10512 22742 10568
rect 22798 10512 22803 10568
rect 16573 10510 22803 10512
rect 16573 10507 16639 10510
rect 22737 10507 22803 10510
rect 20621 10434 20687 10437
rect 21357 10434 21423 10437
rect 23381 10434 23447 10437
rect 20621 10432 23447 10434
rect 20621 10376 20626 10432
rect 20682 10376 21362 10432
rect 21418 10376 23386 10432
rect 23442 10376 23447 10432
rect 20621 10374 23447 10376
rect 20621 10371 20687 10374
rect 21357 10371 21423 10374
rect 23381 10371 23447 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1577 10298 1643 10301
rect 200 10296 1643 10298
rect 200 10240 1582 10296
rect 1638 10240 1643 10296
rect 200 10238 1643 10240
rect 200 10208 800 10238
rect 1577 10235 1643 10238
rect 20529 10298 20595 10301
rect 23933 10298 23999 10301
rect 20529 10296 23999 10298
rect 20529 10240 20534 10296
rect 20590 10240 23938 10296
rect 23994 10240 23999 10296
rect 20529 10238 23999 10240
rect 20529 10235 20595 10238
rect 23933 10235 23999 10238
rect 38285 10298 38351 10301
rect 39200 10298 39800 10328
rect 38285 10296 39800 10298
rect 38285 10240 38290 10296
rect 38346 10240 39800 10296
rect 38285 10238 39800 10240
rect 38285 10235 38351 10238
rect 39200 10208 39800 10238
rect 15377 10162 15443 10165
rect 17953 10162 18019 10165
rect 15377 10160 18019 10162
rect 15377 10104 15382 10160
rect 15438 10104 17958 10160
rect 18014 10104 18019 10160
rect 15377 10102 18019 10104
rect 15377 10099 15443 10102
rect 17953 10099 18019 10102
rect 16205 10026 16271 10029
rect 24853 10026 24919 10029
rect 16205 10024 24919 10026
rect 16205 9968 16210 10024
rect 16266 9968 24858 10024
rect 24914 9968 24919 10024
rect 16205 9966 24919 9968
rect 16205 9963 16271 9966
rect 24853 9963 24919 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 22461 9754 22527 9757
rect 28441 9754 28507 9757
rect 22461 9752 28507 9754
rect 22461 9696 22466 9752
rect 22522 9696 28446 9752
rect 28502 9696 28507 9752
rect 22461 9694 28507 9696
rect 22461 9691 22527 9694
rect 28441 9691 28507 9694
rect 15377 9618 15443 9621
rect 27613 9618 27679 9621
rect 15377 9616 27679 9618
rect 15377 9560 15382 9616
rect 15438 9560 27618 9616
rect 27674 9560 27679 9616
rect 15377 9558 27679 9560
rect 15377 9555 15443 9558
rect 27613 9555 27679 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 15745 9210 15811 9213
rect 17309 9210 17375 9213
rect 15745 9208 17375 9210
rect 15745 9152 15750 9208
rect 15806 9152 17314 9208
rect 17370 9152 17375 9208
rect 15745 9150 17375 9152
rect 15745 9147 15811 9150
rect 17309 9147 17375 9150
rect 22093 9210 22159 9213
rect 23197 9210 23263 9213
rect 22093 9208 23263 9210
rect 22093 9152 22098 9208
rect 22154 9152 23202 9208
rect 23258 9152 23263 9208
rect 22093 9150 23263 9152
rect 22093 9147 22159 9150
rect 23197 9147 23263 9150
rect 200 8938 800 8968
rect 1577 8938 1643 8941
rect 200 8936 1643 8938
rect 200 8880 1582 8936
rect 1638 8880 1643 8936
rect 200 8878 1643 8880
rect 200 8848 800 8878
rect 1577 8875 1643 8878
rect 13813 8938 13879 8941
rect 24853 8938 24919 8941
rect 13813 8936 24919 8938
rect 13813 8880 13818 8936
rect 13874 8880 24858 8936
rect 24914 8880 24919 8936
rect 13813 8878 24919 8880
rect 13813 8875 13879 8878
rect 24853 8875 24919 8878
rect 16573 8802 16639 8805
rect 18505 8802 18571 8805
rect 16573 8800 18571 8802
rect 16573 8744 16578 8800
rect 16634 8744 18510 8800
rect 18566 8744 18571 8800
rect 16573 8742 18571 8744
rect 16573 8739 16639 8742
rect 18505 8739 18571 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 17217 8666 17283 8669
rect 18321 8666 18387 8669
rect 17217 8664 18387 8666
rect 17217 8608 17222 8664
rect 17278 8608 18326 8664
rect 18382 8608 18387 8664
rect 17217 8606 18387 8608
rect 17217 8603 17283 8606
rect 18321 8603 18387 8606
rect 29545 8666 29611 8669
rect 33041 8666 33107 8669
rect 29545 8664 33107 8666
rect 29545 8608 29550 8664
rect 29606 8608 33046 8664
rect 33102 8608 33107 8664
rect 29545 8606 33107 8608
rect 29545 8603 29611 8606
rect 33041 8603 33107 8606
rect 14273 8530 14339 8533
rect 25037 8530 25103 8533
rect 14273 8528 25103 8530
rect 14273 8472 14278 8528
rect 14334 8472 25042 8528
rect 25098 8472 25103 8528
rect 14273 8470 25103 8472
rect 14273 8467 14339 8470
rect 25037 8467 25103 8470
rect 29545 8394 29611 8397
rect 35985 8394 36051 8397
rect 29545 8392 36051 8394
rect 29545 8336 29550 8392
rect 29606 8336 35990 8392
rect 36046 8336 36051 8392
rect 29545 8334 36051 8336
rect 29545 8331 29611 8334
rect 35985 8331 36051 8334
rect 13905 8258 13971 8261
rect 18873 8258 18939 8261
rect 13905 8256 18939 8258
rect 13905 8200 13910 8256
rect 13966 8200 18878 8256
rect 18934 8200 18939 8256
rect 13905 8198 18939 8200
rect 13905 8195 13971 8198
rect 18873 8195 18939 8198
rect 37181 8258 37247 8261
rect 39200 8258 39800 8288
rect 37181 8256 39800 8258
rect 37181 8200 37186 8256
rect 37242 8200 39800 8256
rect 37181 8198 39800 8200
rect 37181 8195 37247 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 13629 8122 13695 8125
rect 18873 8122 18939 8125
rect 13629 8120 18939 8122
rect 13629 8064 13634 8120
rect 13690 8064 18878 8120
rect 18934 8064 18939 8120
rect 13629 8062 18939 8064
rect 13629 8059 13695 8062
rect 18873 8059 18939 8062
rect 19333 8122 19399 8125
rect 21541 8122 21607 8125
rect 19333 8120 21607 8122
rect 19333 8064 19338 8120
rect 19394 8064 21546 8120
rect 21602 8064 21607 8120
rect 19333 8062 21607 8064
rect 19333 8059 19399 8062
rect 21541 8059 21607 8062
rect 15285 7986 15351 7989
rect 36629 7986 36695 7989
rect 15285 7984 36695 7986
rect 15285 7928 15290 7984
rect 15346 7928 36634 7984
rect 36690 7928 36695 7984
rect 15285 7926 36695 7928
rect 15285 7923 15351 7926
rect 36629 7923 36695 7926
rect 17401 7850 17467 7853
rect 21449 7850 21515 7853
rect 17401 7848 21515 7850
rect 17401 7792 17406 7848
rect 17462 7792 21454 7848
rect 21510 7792 21515 7848
rect 17401 7790 21515 7792
rect 17401 7787 17467 7790
rect 21449 7787 21515 7790
rect 22093 7714 22159 7717
rect 22737 7714 22803 7717
rect 22093 7712 22803 7714
rect 22093 7656 22098 7712
rect 22154 7656 22742 7712
rect 22798 7656 22803 7712
rect 22093 7654 22803 7656
rect 22093 7651 22159 7654
rect 22737 7651 22803 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 19333 7578 19399 7581
rect 24485 7578 24551 7581
rect 24710 7578 24716 7580
rect 19333 7576 19442 7578
rect 19333 7520 19338 7576
rect 19394 7520 19442 7576
rect 19333 7515 19442 7520
rect 24485 7576 24716 7578
rect 24485 7520 24490 7576
rect 24546 7520 24716 7576
rect 24485 7518 24716 7520
rect 24485 7515 24551 7518
rect 24710 7516 24716 7518
rect 24780 7516 24786 7580
rect 19382 7442 19442 7515
rect 19609 7442 19675 7445
rect 19382 7440 19675 7442
rect 19382 7384 19614 7440
rect 19670 7384 19675 7440
rect 19382 7382 19675 7384
rect 19609 7379 19675 7382
rect 19885 7442 19951 7445
rect 20253 7442 20319 7445
rect 19885 7440 20319 7442
rect 19885 7384 19890 7440
rect 19946 7384 20258 7440
rect 20314 7384 20319 7440
rect 19885 7382 20319 7384
rect 19885 7379 19951 7382
rect 20253 7379 20319 7382
rect 16573 7306 16639 7309
rect 28993 7306 29059 7309
rect 16573 7304 29059 7306
rect 16573 7248 16578 7304
rect 16634 7248 28998 7304
rect 29054 7248 29059 7304
rect 16573 7246 29059 7248
rect 16573 7243 16639 7246
rect 28993 7243 29059 7246
rect 14825 7170 14891 7173
rect 22001 7170 22067 7173
rect 14825 7168 22067 7170
rect 14825 7112 14830 7168
rect 14886 7112 22006 7168
rect 22062 7112 22067 7168
rect 14825 7110 22067 7112
rect 14825 7107 14891 7110
rect 22001 7107 22067 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 13813 7034 13879 7037
rect 28533 7034 28599 7037
rect 32213 7034 32279 7037
rect 32673 7034 32739 7037
rect 13813 7032 32739 7034
rect 13813 6976 13818 7032
rect 13874 6976 28538 7032
rect 28594 6976 32218 7032
rect 32274 6976 32678 7032
rect 32734 6976 32739 7032
rect 13813 6974 32739 6976
rect 13813 6971 13879 6974
rect 28533 6971 28599 6974
rect 32213 6971 32279 6974
rect 32673 6971 32739 6974
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 17217 6898 17283 6901
rect 21725 6898 21791 6901
rect 17217 6896 21791 6898
rect 17217 6840 17222 6896
rect 17278 6840 21730 6896
rect 21786 6840 21791 6896
rect 17217 6838 21791 6840
rect 17217 6835 17283 6838
rect 21725 6835 21791 6838
rect 17033 6762 17099 6765
rect 24853 6762 24919 6765
rect 17033 6760 24919 6762
rect 17033 6704 17038 6760
rect 17094 6704 24858 6760
rect 24914 6704 24919 6760
rect 17033 6702 24919 6704
rect 17033 6699 17099 6702
rect 24853 6699 24919 6702
rect 21541 6626 21607 6629
rect 23933 6626 23999 6629
rect 21541 6624 23999 6626
rect 21541 6568 21546 6624
rect 21602 6568 23938 6624
rect 23994 6568 23999 6624
rect 21541 6566 23999 6568
rect 21541 6563 21607 6566
rect 23933 6563 23999 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 19149 6354 19215 6357
rect 22277 6354 22343 6357
rect 19149 6352 22343 6354
rect 19149 6296 19154 6352
rect 19210 6296 22282 6352
rect 22338 6296 22343 6352
rect 19149 6294 22343 6296
rect 19149 6291 19215 6294
rect 22277 6291 22343 6294
rect 20253 6218 20319 6221
rect 24577 6218 24643 6221
rect 28257 6218 28323 6221
rect 20253 6216 28323 6218
rect 20253 6160 20258 6216
rect 20314 6160 24582 6216
rect 24638 6160 28262 6216
rect 28318 6160 28323 6216
rect 20253 6158 28323 6160
rect 20253 6155 20319 6158
rect 24577 6155 24643 6158
rect 28257 6155 28323 6158
rect 38193 6218 38259 6221
rect 39200 6218 39800 6248
rect 38193 6216 39800 6218
rect 38193 6160 38198 6216
rect 38254 6160 39800 6216
rect 38193 6158 39800 6160
rect 38193 6155 38259 6158
rect 39200 6128 39800 6158
rect 20161 6082 20227 6085
rect 28901 6082 28967 6085
rect 20161 6080 28967 6082
rect 20161 6024 20166 6080
rect 20222 6024 28906 6080
rect 28962 6024 28967 6080
rect 20161 6022 28967 6024
rect 20161 6019 20227 6022
rect 28901 6019 28967 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 13169 5946 13235 5949
rect 19149 5946 19215 5949
rect 13169 5944 19215 5946
rect 13169 5888 13174 5944
rect 13230 5888 19154 5944
rect 19210 5888 19215 5944
rect 13169 5886 19215 5888
rect 13169 5883 13235 5886
rect 19149 5883 19215 5886
rect 15193 5810 15259 5813
rect 25313 5810 25379 5813
rect 15193 5808 25379 5810
rect 15193 5752 15198 5808
rect 15254 5752 25318 5808
rect 25374 5752 25379 5808
rect 15193 5750 25379 5752
rect 15193 5747 15259 5750
rect 25313 5747 25379 5750
rect 16205 5674 16271 5677
rect 30465 5674 30531 5677
rect 16205 5672 30531 5674
rect 16205 5616 16210 5672
rect 16266 5616 30470 5672
rect 30526 5616 30531 5672
rect 16205 5614 30531 5616
rect 16205 5611 16271 5614
rect 30465 5611 30531 5614
rect 14917 5538 14983 5541
rect 18781 5538 18847 5541
rect 14917 5536 18847 5538
rect 14917 5480 14922 5536
rect 14978 5480 18786 5536
rect 18842 5480 18847 5536
rect 14917 5478 18847 5480
rect 14917 5475 14983 5478
rect 18781 5475 18847 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 16941 5402 17007 5405
rect 19149 5402 19215 5405
rect 16941 5400 19215 5402
rect 16941 5344 16946 5400
rect 17002 5344 19154 5400
rect 19210 5344 19215 5400
rect 16941 5342 19215 5344
rect 16941 5339 17007 5342
rect 19149 5339 19215 5342
rect 21357 5402 21423 5405
rect 24025 5402 24091 5405
rect 21357 5400 24091 5402
rect 21357 5344 21362 5400
rect 21418 5344 24030 5400
rect 24086 5344 24091 5400
rect 21357 5342 24091 5344
rect 21357 5339 21423 5342
rect 24025 5339 24091 5342
rect 20805 5266 20871 5269
rect 25313 5266 25379 5269
rect 20805 5264 25379 5266
rect 20805 5208 20810 5264
rect 20866 5208 25318 5264
rect 25374 5208 25379 5264
rect 20805 5206 25379 5208
rect 20805 5203 20871 5206
rect 25313 5203 25379 5206
rect 16021 5130 16087 5133
rect 18781 5130 18847 5133
rect 16021 5128 18847 5130
rect 16021 5072 16026 5128
rect 16082 5072 18786 5128
rect 18842 5072 18847 5128
rect 16021 5070 18847 5072
rect 16021 5067 16087 5070
rect 18781 5067 18847 5070
rect 21173 5130 21239 5133
rect 23841 5130 23907 5133
rect 21173 5128 23907 5130
rect 21173 5072 21178 5128
rect 21234 5072 23846 5128
rect 23902 5072 23907 5128
rect 21173 5070 23907 5072
rect 21173 5067 21239 5070
rect 23841 5067 23907 5070
rect 16573 4994 16639 4997
rect 18689 4994 18755 4997
rect 16573 4992 18755 4994
rect 16573 4936 16578 4992
rect 16634 4936 18694 4992
rect 18750 4936 18755 4992
rect 16573 4934 18755 4936
rect 16573 4931 16639 4934
rect 18689 4931 18755 4934
rect 19333 4994 19399 4997
rect 24393 4994 24459 4997
rect 19333 4992 24459 4994
rect 19333 4936 19338 4992
rect 19394 4936 24398 4992
rect 24454 4936 24459 4992
rect 19333 4934 24459 4936
rect 19333 4931 19399 4934
rect 24393 4931 24459 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 200 4856 1735 4858
rect 200 4800 1674 4856
rect 1730 4800 1735 4856
rect 200 4798 1735 4800
rect 200 4768 800 4798
rect 1669 4795 1735 4798
rect 16113 4858 16179 4861
rect 18689 4858 18755 4861
rect 16113 4856 18755 4858
rect 16113 4800 16118 4856
rect 16174 4800 18694 4856
rect 18750 4800 18755 4856
rect 16113 4798 18755 4800
rect 16113 4795 16179 4798
rect 18689 4795 18755 4798
rect 21909 4858 21975 4861
rect 22093 4858 22159 4861
rect 21909 4856 22159 4858
rect 21909 4800 21914 4856
rect 21970 4800 22098 4856
rect 22154 4800 22159 4856
rect 21909 4798 22159 4800
rect 21909 4795 21975 4798
rect 22093 4795 22159 4798
rect 38193 4858 38259 4861
rect 39200 4858 39800 4888
rect 38193 4856 39800 4858
rect 38193 4800 38198 4856
rect 38254 4800 39800 4856
rect 38193 4798 39800 4800
rect 38193 4795 38259 4798
rect 39200 4768 39800 4798
rect 16849 4722 16915 4725
rect 17309 4722 17375 4725
rect 16849 4720 17375 4722
rect 16849 4664 16854 4720
rect 16910 4664 17314 4720
rect 17370 4664 17375 4720
rect 16849 4662 17375 4664
rect 16849 4659 16915 4662
rect 17309 4659 17375 4662
rect 17861 4722 17927 4725
rect 24761 4722 24827 4725
rect 17861 4720 24827 4722
rect 17861 4664 17866 4720
rect 17922 4664 24766 4720
rect 24822 4664 24827 4720
rect 17861 4662 24827 4664
rect 17861 4659 17927 4662
rect 24761 4659 24827 4662
rect 15929 4586 15995 4589
rect 24945 4586 25011 4589
rect 15929 4584 25011 4586
rect 15929 4528 15934 4584
rect 15990 4528 24950 4584
rect 25006 4528 25011 4584
rect 15929 4526 25011 4528
rect 15929 4523 15995 4526
rect 24945 4523 25011 4526
rect 10409 4450 10475 4453
rect 16297 4450 16363 4453
rect 17309 4450 17375 4453
rect 10409 4448 17375 4450
rect 10409 4392 10414 4448
rect 10470 4392 16302 4448
rect 16358 4392 17314 4448
rect 17370 4392 17375 4448
rect 10409 4390 17375 4392
rect 10409 4387 10475 4390
rect 16297 4387 16363 4390
rect 17309 4387 17375 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 22093 4314 22159 4317
rect 25129 4314 25195 4317
rect 22093 4312 25195 4314
rect 22093 4256 22098 4312
rect 22154 4256 25134 4312
rect 25190 4256 25195 4312
rect 22093 4254 25195 4256
rect 22093 4251 22159 4254
rect 25129 4251 25195 4254
rect 14089 4042 14155 4045
rect 17953 4042 18019 4045
rect 14089 4040 18019 4042
rect 14089 3984 14094 4040
rect 14150 3984 17958 4040
rect 18014 3984 18019 4040
rect 14089 3982 18019 3984
rect 14089 3979 14155 3982
rect 17953 3979 18019 3982
rect 21449 4042 21515 4045
rect 26601 4042 26667 4045
rect 21449 4040 26667 4042
rect 21449 3984 21454 4040
rect 21510 3984 26606 4040
rect 26662 3984 26667 4040
rect 21449 3982 26667 3984
rect 21449 3979 21515 3982
rect 26601 3979 26667 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 21909 3770 21975 3773
rect 23565 3770 23631 3773
rect 21909 3768 23631 3770
rect 21909 3712 21914 3768
rect 21970 3712 23570 3768
rect 23626 3712 23631 3768
rect 21909 3710 23631 3712
rect 21909 3707 21975 3710
rect 23565 3707 23631 3710
rect 21633 3634 21699 3637
rect 23473 3634 23539 3637
rect 21633 3632 23539 3634
rect 21633 3576 21638 3632
rect 21694 3576 23478 3632
rect 23534 3576 23539 3632
rect 21633 3574 23539 3576
rect 21633 3571 21699 3574
rect 23473 3571 23539 3574
rect 200 3498 800 3528
rect 1577 3498 1643 3501
rect 200 3496 1643 3498
rect 200 3440 1582 3496
rect 1638 3440 1643 3496
rect 200 3438 1643 3440
rect 200 3408 800 3438
rect 1577 3435 1643 3438
rect 1761 3498 1827 3501
rect 26233 3498 26299 3501
rect 1761 3496 26299 3498
rect 1761 3440 1766 3496
rect 1822 3440 26238 3496
rect 26294 3440 26299 3496
rect 1761 3438 26299 3440
rect 1761 3435 1827 3438
rect 26233 3435 26299 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 15745 3226 15811 3229
rect 18781 3226 18847 3229
rect 15745 3224 18847 3226
rect 15745 3168 15750 3224
rect 15806 3168 18786 3224
rect 18842 3168 18847 3224
rect 15745 3166 18847 3168
rect 15745 3163 15811 3166
rect 18781 3163 18847 3166
rect 20989 3226 21055 3229
rect 25773 3226 25839 3229
rect 20989 3224 25839 3226
rect 20989 3168 20994 3224
rect 21050 3168 25778 3224
rect 25834 3168 25839 3224
rect 20989 3166 25839 3168
rect 20989 3163 21055 3166
rect 25773 3163 25839 3166
rect 31753 3226 31819 3229
rect 33685 3226 33751 3229
rect 31753 3224 33751 3226
rect 31753 3168 31758 3224
rect 31814 3168 33690 3224
rect 33746 3168 33751 3224
rect 31753 3166 33751 3168
rect 31753 3163 31819 3166
rect 33685 3163 33751 3166
rect 31293 2954 31359 2957
rect 31753 2954 31819 2957
rect 31293 2952 31819 2954
rect 31293 2896 31298 2952
rect 31354 2896 31758 2952
rect 31814 2896 31819 2952
rect 31293 2894 31819 2896
rect 31293 2891 31359 2894
rect 31753 2891 31819 2894
rect 19425 2818 19491 2821
rect 22185 2818 22251 2821
rect 19425 2816 22251 2818
rect 19425 2760 19430 2816
rect 19486 2760 22190 2816
rect 22246 2760 22251 2816
rect 19425 2758 22251 2760
rect 19425 2755 19491 2758
rect 22185 2755 22251 2758
rect 38285 2818 38351 2821
rect 39200 2818 39800 2848
rect 38285 2816 39800 2818
rect 38285 2760 38290 2816
rect 38346 2760 39800 2816
rect 38285 2758 39800 2760
rect 38285 2755 38351 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 37181 1458 37247 1461
rect 37181 1456 39314 1458
rect 37181 1400 37186 1456
rect 37242 1400 39314 1456
rect 37181 1398 39314 1400
rect 37181 1395 37247 1398
rect 39254 1050 39314 1398
rect 39070 990 39314 1050
rect 39070 778 39130 990
rect 39200 778 39800 808
rect 39070 718 39800 778
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 24716 15404 24780 15468
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 26188 15056 26252 15060
rect 26188 15000 26202 15056
rect 26202 15000 26252 15056
rect 26188 14996 26252 15000
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 26188 13968 26252 13972
rect 26188 13912 26202 13968
rect 26202 13912 26252 13968
rect 26188 13908 26252 13912
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 24716 7516 24780 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 24715 15468 24781 15469
rect 24715 15404 24716 15468
rect 24780 15404 24781 15468
rect 24715 15403 24781 15404
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 24718 7581 24778 15403
rect 26187 15060 26253 15061
rect 26187 14996 26188 15060
rect 26252 14996 26253 15060
rect 26187 14995 26253 14996
rect 26190 13973 26250 14995
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 26187 13972 26253 13973
rect 26187 13908 26188 13972
rect 26252 13908 26253 13972
rect 26187 13907 26253 13908
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 24715 7580 24781 7581
rect 24715 7516 24716 7580
rect 24780 7516 24781 7580
rect 24715 7515 24781 7516
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1667941163
transform -1 0 31648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform -1 0 28980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 16008 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1667941163
transform -1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1667941163
transform -1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1667941163
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1667941163
transform 1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1667941163
transform 1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform -1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1667941163
transform -1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1667941163
transform -1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1667941163
transform -1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1667941163
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1667941163
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1667941163
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform -1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1667941163
transform -1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform 1 0 28336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform -1 0 31648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1667941163
transform -1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform -1 0 24656 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1667941163
transform -1 0 14904 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform 1 0 29348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1667941163
transform -1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform 1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform 1 0 25852 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1667941163
transform -1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1667941163
transform -1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1667941163
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1667941163
transform -1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1667941163
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform 1 0 28980 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1667941163
transform 1 0 31648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 1667941163
transform -1 0 11960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1667941163
transform -1 0 32200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform -1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform -1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1667941163
transform -1 0 12604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1667941163
transform -1 0 32384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1667941163
transform -1 0 15824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1667941163
transform -1 0 17112 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform 1 0 21160 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1667941163
transform 1 0 2944 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1667941163
transform -1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1667941163
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform -1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform -1 0 13248 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1667941163
transform 1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform 1 0 13248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform -1 0 32476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1667941163
transform -1 0 10028 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 31556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform 1 0 18308 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform -1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform -1 0 20424 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform -1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform 1 0 17480 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform 1 0 28244 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform -1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1667941163
transform -1 0 32384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform -1 0 23736 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform -1 0 33304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1667941163
transform 1 0 12328 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1667941163
transform 1 0 31188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform 1 0 31464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1667941163
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1667941163
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1667941163
transform 1 0 35880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform 1 0 36524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1667941163
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform 1 0 26496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1667941163
transform 1 0 26496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform -1 0 12328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1667941163
transform 1 0 37076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1667941163
transform 1 0 36248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1667941163
transform 1 0 37628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1667941163
transform 1 0 34132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1667941163
transform -1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1667941163
transform 1 0 33028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1667941163
transform 1 0 35972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1667941163
transform -1 0 37812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1667941163
transform 1 0 36064 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1667941163
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform 1 0 34500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1667941163
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1667941163
transform 1 0 35972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1667941163
transform 1 0 34408 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1667941163
transform 1 0 31924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1667941163
transform 1 0 31280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1667941163
transform -1 0 36708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1667941163
transform 1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1667941163
transform 1 0 20056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1667941163
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1667941163
transform -1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 14904 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1667941163
transform 1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1667941163
transform -1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1667941163
transform 1 0 36800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1667941163
transform -1 0 33580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1667941163
transform 1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1667941163
transform -1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1667941163
transform 1 0 20608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1667941163
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1667941163
transform 1 0 13064 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1667941163
transform 1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__CLK
timestamp 1667941163
transform 1 0 35512 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__CLK
timestamp 1667941163
transform 1 0 34132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__CLK
timestamp 1667941163
transform 1 0 20792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__CLK
timestamp 1667941163
transform 1 0 30912 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__D
timestamp 1667941163
transform 1 0 30360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__CLK
timestamp 1667941163
transform 1 0 28980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__D
timestamp 1667941163
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__CLK
timestamp 1667941163
transform 1 0 35788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__D
timestamp 1667941163
transform -1 0 35420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1667941163
transform 1 0 36524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1667941163
transform 1 0 33580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1667941163
transform 1 0 32108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__D
timestamp 1667941163
transform 1 0 31096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1667941163
transform 1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__D
timestamp 1667941163
transform -1 0 32660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1667941163
transform 1 0 34408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1667941163
transform 1 0 38180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1667941163
transform 1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1667941163
transform -1 0 37260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1667941163
transform 1 0 32844 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1667941163
transform 1 0 33396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1667941163
transform 1 0 34960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1667941163
transform 1 0 38180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__D
timestamp 1667941163
transform -1 0 34132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1667941163
transform 1 0 35972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1667941163
transform 1 0 33304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__D
timestamp 1667941163
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1667941163
transform 1 0 31464 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1667941163
transform 1 0 33672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__D
timestamp 1667941163
transform -1 0 33304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1667941163
transform 1 0 35420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1667941163
transform 1 0 32936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1667941163
transform 1 0 34868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1667941163
transform 1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__D
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1667941163
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__D
timestamp 1667941163
transform -1 0 20976 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1667941163
transform 1 0 30728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__D
timestamp 1667941163
transform 1 0 30176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__D
timestamp 1667941163
transform -1 0 35052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1667941163
transform 1 0 34132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1667941163
transform 1 0 34868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1667941163
transform 1 0 34960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__D
timestamp 1667941163
transform -1 0 34132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1667941163
transform 1 0 32844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1667941163
transform 1 0 33120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__D
timestamp 1667941163
transform -1 0 33856 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1667941163
transform 1 0 34132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1667941163
transform 1 0 35512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1667941163
transform 1 0 36708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1667941163
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__D
timestamp 1667941163
transform -1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1667941163
transform 1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1667941163
transform 1 0 32568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__D
timestamp 1667941163
transform -1 0 32200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1667941163
transform 1 0 33580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1667941163
transform 1 0 36524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1667941163
transform 1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1667941163
transform 1 0 33488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__D
timestamp 1667941163
transform -1 0 34040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1667941163
transform 1 0 32476 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__CLK
timestamp 1667941163
transform 1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__D
timestamp 1667941163
transform -1 0 33212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__CLK
timestamp 1667941163
transform 1 0 32292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__CLK
timestamp 1667941163
transform 1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__CLK
timestamp 1667941163
transform 1 0 31648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__CLK
timestamp 1667941163
transform 1 0 32844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__CLK
timestamp 1667941163
transform 1 0 32292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__CLK
timestamp 1667941163
transform 1 0 20240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__D
timestamp 1667941163
transform -1 0 20976 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__CLK
timestamp 1667941163
transform 1 0 30820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__CLK
timestamp 1667941163
transform 1 0 31924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__CLK
timestamp 1667941163
transform 1 0 33396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__CLK
timestamp 1667941163
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__CLK
timestamp 1667941163
transform 1 0 31556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__CLK
timestamp 1667941163
transform 1 0 30912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__CLK
timestamp 1667941163
transform 1 0 32568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__CLK
timestamp 1667941163
transform 1 0 34868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__CLK
timestamp 1667941163
transform 1 0 32844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__CLK
timestamp 1667941163
transform 1 0 31004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__CLK
timestamp 1667941163
transform 1 0 19688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__CLK
timestamp 1667941163
transform 1 0 19504 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__CLK
timestamp 1667941163
transform 1 0 33396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1667941163
transform 1 0 25208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1667941163
transform -1 0 21988 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1667941163
transform -1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1667941163
transform -1 0 20148 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1667941163
transform -1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1667941163
transform -1 0 30544 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1667941163
transform -1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1667941163
transform 1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1667941163
transform -1 0 28244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1667941163
transform -1 0 4140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1667941163
transform 1 0 5336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1667941163
transform -1 0 22264 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1667941163
transform 1 0 36616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1667941163
transform 1 0 20056 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1667941163
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1667941163
transform -1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1667941163
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A
timestamp 1667941163
transform 1 0 26404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1667941163
transform -1 0 7912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1667941163
transform 1 0 23000 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1667941163
transform 1 0 30636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1667941163
transform -1 0 9476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1667941163
transform -1 0 19228 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__A
timestamp 1667941163
transform -1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__A
timestamp 1667941163
transform -1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__A
timestamp 1667941163
transform -1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 35788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 37628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 37628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 36708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 1748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 37628 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 1748 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 37628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 1748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 7452 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 36800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 37628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 34040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 37720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 35604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1667941163
transform 1 0 36800 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1667941163
transform 1 0 37444 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1667941163
transform 1 0 1932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1667941163
transform -1 0 28060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1667941163
transform -1 0 35236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1667941163
transform -1 0 20976 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform 1 0 37444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1667941163
transform -1 0 12604 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1667941163
transform 1 0 13340 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1667941163
transform -1 0 36892 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1667941163
transform -1 0 5520 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1667941163
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1667941163
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1667941163
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_147
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156
timestamp 1667941163
transform 1 0 15456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186
timestamp 1667941163
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1667941163
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1667941163
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1667941163
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1667941163
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_42
timestamp 1667941163
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_80
timestamp 1667941163
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_92
timestamp 1667941163
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1667941163
transform 1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1667941163
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_122
timestamp 1667941163
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1667941163
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1667941163
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1667941163
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_160
timestamp 1667941163
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1667941163
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_186
timestamp 1667941163
transform 1 0 18216 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1667941163
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_201
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1667941163
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1667941163
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1667941163
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1667941163
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1667941163
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1667941163
transform 1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_379
timestamp 1667941163
transform 1 0 35972 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1667941163
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1667941163
transform 1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_14
timestamp 1667941163
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1667941163
transform 1 0 11868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_129
timestamp 1667941163
transform 1 0 12972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_132
timestamp 1667941163
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_156
timestamp 1667941163
transform 1 0 15456 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1667941163
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_210
timestamp 1667941163
transform 1 0 20424 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_218
timestamp 1667941163
transform 1 0 21160 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_239
timestamp 1667941163
transform 1 0 23092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1667941163
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_299
timestamp 1667941163
transform 1 0 28612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1667941163
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1667941163
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_355
timestamp 1667941163
transform 1 0 33764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1667941163
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1667941163
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_375
timestamp 1667941163
transform 1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_381
timestamp 1667941163
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_387
timestamp 1667941163
transform 1 0 36708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_393
timestamp 1667941163
transform 1 0 37260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1667941163
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1667941163
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1667941163
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1667941163
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1667941163
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1667941163
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_195
timestamp 1667941163
transform 1 0 19044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_201
timestamp 1667941163
transform 1 0 19596 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1667941163
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_210
timestamp 1667941163
transform 1 0 20424 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_216
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_231
timestamp 1667941163
transform 1 0 22356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1667941163
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1667941163
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_303
timestamp 1667941163
transform 1 0 28980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_327
timestamp 1667941163
transform 1 0 31188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1667941163
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_346
timestamp 1667941163
transform 1 0 32936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_352
timestamp 1667941163
transform 1 0 33488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_358
timestamp 1667941163
transform 1 0 34040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_364
timestamp 1667941163
transform 1 0 34592 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_370
timestamp 1667941163
transform 1 0 35144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_376
timestamp 1667941163
transform 1 0 35696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_382
timestamp 1667941163
transform 1 0 36248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_386
timestamp 1667941163
transform 1 0 36616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1667941163
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_399
timestamp 1667941163
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_102
timestamp 1667941163
transform 1 0 10488 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_114
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_126
timestamp 1667941163
transform 1 0 12696 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1667941163
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1667941163
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1667941163
transform 1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1667941163
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_168
timestamp 1667941163
transform 1 0 16560 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1667941163
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_188
timestamp 1667941163
transform 1 0 18400 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1667941163
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1667941163
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1667941163
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_238
timestamp 1667941163
transform 1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_246
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1667941163
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_281
timestamp 1667941163
transform 1 0 26956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1667941163
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_331
timestamp 1667941163
transform 1 0 31556 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_342
timestamp 1667941163
transform 1 0 32568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_348
timestamp 1667941163
transform 1 0 33120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_354
timestamp 1667941163
transform 1 0 33672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1667941163
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_369
timestamp 1667941163
transform 1 0 35052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_376
timestamp 1667941163
transform 1 0 35696 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_383
timestamp 1667941163
transform 1 0 36340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_400
timestamp 1667941163
transform 1 0 37904 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1667941163
transform 1 0 38456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_124
timestamp 1667941163
transform 1 0 12512 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_132
timestamp 1667941163
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1667941163
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1667941163
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_148
timestamp 1667941163
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_155
timestamp 1667941163
transform 1 0 15364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1667941163
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_174
timestamp 1667941163
transform 1 0 17112 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1667941163
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_197
timestamp 1667941163
transform 1 0 19228 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1667941163
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1667941163
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_248
timestamp 1667941163
transform 1 0 23920 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_272
timestamp 1667941163
transform 1 0 26128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1667941163
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_286
timestamp 1667941163
transform 1 0 27416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_294
timestamp 1667941163
transform 1 0 28152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1667941163
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_344
timestamp 1667941163
transform 1 0 32752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_348
timestamp 1667941163
transform 1 0 33120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_352
timestamp 1667941163
transform 1 0 33488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_358
timestamp 1667941163
transform 1 0 34040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_364
timestamp 1667941163
transform 1 0 34592 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_370
timestamp 1667941163
transform 1 0 35144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_376
timestamp 1667941163
transform 1 0 35696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_382
timestamp 1667941163
transform 1 0 36248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1667941163
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_397
timestamp 1667941163
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1667941163
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_122
timestamp 1667941163
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp 1667941163
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1667941163
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_152
timestamp 1667941163
transform 1 0 15088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1667941163
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_166
timestamp 1667941163
transform 1 0 16376 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1667941163
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1667941163
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1667941163
transform 1 0 19596 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_204
timestamp 1667941163
transform 1 0 19872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1667941163
transform 1 0 20424 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_216
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_243
timestamp 1667941163
transform 1 0 23460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1667941163
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_275
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1667941163
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1667941163
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_355
timestamp 1667941163
transform 1 0 33764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1667941163
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_369
timestamp 1667941163
transform 1 0 35052 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1667941163
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_381
timestamp 1667941163
transform 1 0 36156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_387
timestamp 1667941163
transform 1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1667941163
transform 1 0 37260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_399
timestamp 1667941163
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1667941163
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1667941163
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1667941163
transform 1 0 13892 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1667941163
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_173
timestamp 1667941163
transform 1 0 17020 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_177
timestamp 1667941163
transform 1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_190
timestamp 1667941163
transform 1 0 18584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_203
timestamp 1667941163
transform 1 0 19780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1667941163
transform 1 0 20424 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_216
timestamp 1667941163
transform 1 0 20976 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_248
timestamp 1667941163
transform 1 0 23920 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_254
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_290
timestamp 1667941163
transform 1 0 27784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_312
timestamp 1667941163
transform 1 0 29808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_319
timestamp 1667941163
transform 1 0 30452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_325
timestamp 1667941163
transform 1 0 31004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 1667941163
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_341
timestamp 1667941163
transform 1 0 32476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_347
timestamp 1667941163
transform 1 0 33028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_353
timestamp 1667941163
transform 1 0 33580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_359
timestamp 1667941163
transform 1 0 34132 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_365
timestamp 1667941163
transform 1 0 34684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_374
timestamp 1667941163
transform 1 0 35512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_381
timestamp 1667941163
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1667941163
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_397
timestamp 1667941163
transform 1 0 37628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_124
timestamp 1667941163
transform 1 0 12512 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1667941163
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1667941163
transform 1 0 14720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_155
timestamp 1667941163
transform 1 0 15364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 1667941163
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1667941163
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_176
timestamp 1667941163
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_183
timestamp 1667941163
transform 1 0 17940 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1667941163
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1667941163
transform 1 0 21252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_258
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_267
timestamp 1667941163
transform 1 0 25668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1667941163
transform 1 0 28152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1667941163
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_337
timestamp 1667941163
transform 1 0 32108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_343
timestamp 1667941163
transform 1 0 32660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_349
timestamp 1667941163
transform 1 0 33212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_355
timestamp 1667941163
transform 1 0 33764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1667941163
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_369
timestamp 1667941163
transform 1 0 35052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_375
timestamp 1667941163
transform 1 0 35604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_381
timestamp 1667941163
transform 1 0 36156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_387
timestamp 1667941163
transform 1 0 36708 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_393
timestamp 1667941163
transform 1 0 37260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_399
timestamp 1667941163
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1667941163
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_121
timestamp 1667941163
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_128
timestamp 1667941163
transform 1 0 12880 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_134
timestamp 1667941163
transform 1 0 13432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1667941163
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1667941163
transform 1 0 14444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1667941163
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_159
timestamp 1667941163
transform 1 0 15732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_180
timestamp 1667941163
transform 1 0 17664 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_186
timestamp 1667941163
transform 1 0 18216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_190
timestamp 1667941163
transform 1 0 18584 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_203
timestamp 1667941163
transform 1 0 19780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_207
timestamp 1667941163
transform 1 0 20148 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_210
timestamp 1667941163
transform 1 0 20424 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_216
timestamp 1667941163
transform 1 0 20976 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_250
timestamp 1667941163
transform 1 0 24104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_312
timestamp 1667941163
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_318
timestamp 1667941163
transform 1 0 30360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_324
timestamp 1667941163
transform 1 0 30912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_330
timestamp 1667941163
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1667941163
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_347
timestamp 1667941163
transform 1 0 33028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_353
timestamp 1667941163
transform 1 0 33580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1667941163
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1667941163
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_371
timestamp 1667941163
transform 1 0 35236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_377
timestamp 1667941163
transform 1 0 35788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_381
timestamp 1667941163
transform 1 0 36156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_384
timestamp 1667941163
transform 1 0 36432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1667941163
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_398
timestamp 1667941163
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1667941163
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1667941163
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1667941163
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_156
timestamp 1667941163
transform 1 0 15456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_160
timestamp 1667941163
transform 1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1667941163
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_208
timestamp 1667941163
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_215
timestamp 1667941163
transform 1 0 20884 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_279
timestamp 1667941163
transform 1 0 26772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1667941163
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_337
timestamp 1667941163
transform 1 0 32108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_343
timestamp 1667941163
transform 1 0 32660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_349
timestamp 1667941163
transform 1 0 33212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1667941163
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_374
timestamp 1667941163
transform 1 0 35512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_380
timestamp 1667941163
transform 1 0 36064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_388
timestamp 1667941163
transform 1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1667941163
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_402
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1667941163
transform 1 0 38456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1667941163
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1667941163
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1667941163
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_146
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1667941163
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1667941163
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_173
timestamp 1667941163
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_177
timestamp 1667941163
transform 1 0 17388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_190
timestamp 1667941163
transform 1 0 18584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_194
timestamp 1667941163
transform 1 0 18952 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1667941163
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_211
timestamp 1667941163
transform 1 0 20516 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1667941163
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1667941163
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_320
timestamp 1667941163
transform 1 0 30544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_326
timestamp 1667941163
transform 1 0 31096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1667941163
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_341
timestamp 1667941163
transform 1 0 32476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_347
timestamp 1667941163
transform 1 0 33028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_353
timestamp 1667941163
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_359
timestamp 1667941163
transform 1 0 34132 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_371
timestamp 1667941163
transform 1 0 35236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_379
timestamp 1667941163
transform 1 0 35972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_384
timestamp 1667941163
transform 1 0 36432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1667941163
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1667941163
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_129
timestamp 1667941163
transform 1 0 12972 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1667941163
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1667941163
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1667941163
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1667941163
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_240
timestamp 1667941163
transform 1 0 23184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_247
timestamp 1667941163
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_332
timestamp 1667941163
transform 1 0 31648 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_344
timestamp 1667941163
transform 1 0 32752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_350
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_356
timestamp 1667941163
transform 1 0 33856 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_381
timestamp 1667941163
transform 1 0 36156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_387
timestamp 1667941163
transform 1 0 36708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_393
timestamp 1667941163
transform 1 0 37260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_397
timestamp 1667941163
transform 1 0 37628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1667941163
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1667941163
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_91
timestamp 1667941163
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1667941163
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_121
timestamp 1667941163
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 1667941163
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1667941163
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1667941163
transform 1 0 13892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1667941163
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1667941163
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_194
timestamp 1667941163
transform 1 0 18952 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1667941163
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_243
timestamp 1667941163
transform 1 0 23460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_270
timestamp 1667941163
transform 1 0 25944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1667941163
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_290
timestamp 1667941163
transform 1 0 27784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1667941163
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_320
timestamp 1667941163
transform 1 0 30544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_326
timestamp 1667941163
transform 1 0 31096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1667941163
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_342
timestamp 1667941163
transform 1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_355
timestamp 1667941163
transform 1 0 33764 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_397
timestamp 1667941163
transform 1 0 37628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_7
timestamp 1667941163
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1667941163
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 10764 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_129
timestamp 1667941163
transform 1 0 12972 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_132
timestamp 1667941163
transform 1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_150
timestamp 1667941163
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_157
timestamp 1667941163
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1667941163
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1667941163
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_208
timestamp 1667941163
transform 1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_212
timestamp 1667941163
transform 1 0 20608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1667941163
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_243
timestamp 1667941163
transform 1 0 23460 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_262
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1667941163
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_297
timestamp 1667941163
transform 1 0 28428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1667941163
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_332
timestamp 1667941163
transform 1 0 31648 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1667941163
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_344
timestamp 1667941163
transform 1 0 32752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_350
timestamp 1667941163
transform 1 0 33304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_356
timestamp 1667941163
transform 1 0 33856 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_369
timestamp 1667941163
transform 1 0 35052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_373
timestamp 1667941163
transform 1 0 35420 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_379
timestamp 1667941163
transform 1 0 35972 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_391
timestamp 1667941163
transform 1 0 37076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1667941163
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 1667941163
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_91
timestamp 1667941163
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_97
timestamp 1667941163
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1667941163
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1667941163
transform 1 0 12420 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1667941163
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1667941163
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_142
timestamp 1667941163
transform 1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1667941163
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_173
timestamp 1667941163
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1667941163
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1667941163
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_200
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1667941163
transform 1 0 20700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1667941163
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_248
timestamp 1667941163
transform 1 0 23920 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_256
timestamp 1667941163
transform 1 0 24656 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1667941163
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_315
timestamp 1667941163
transform 1 0 30084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_322
timestamp 1667941163
transform 1 0 30728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_328
timestamp 1667941163
transform 1 0 31280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_341
timestamp 1667941163
transform 1 0 32476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_347
timestamp 1667941163
transform 1 0 33028 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_353
timestamp 1667941163
transform 1 0 33580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_365
timestamp 1667941163
transform 1 0 34684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_377
timestamp 1667941163
transform 1 0 35788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1667941163
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_398
timestamp 1667941163
transform 1 0 37720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_117
timestamp 1667941163
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1667941163
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_129
timestamp 1667941163
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1667941163
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_178
timestamp 1667941163
transform 1 0 17480 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1667941163
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1667941163
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_264
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1667941163
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1667941163
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_327
timestamp 1667941163
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_339
timestamp 1667941163
transform 1 0 32292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_347
timestamp 1667941163
transform 1 0 33028 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_352
timestamp 1667941163
transform 1 0 33488 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_119
timestamp 1667941163
transform 1 0 12052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1667941163
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1667941163
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_254
timestamp 1667941163
transform 1 0 24472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1667941163
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_312
timestamp 1667941163
transform 1 0 29808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_319
timestamp 1667941163
transform 1 0 30452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_326
timestamp 1667941163
transform 1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1667941163
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_341
timestamp 1667941163
transform 1 0 32476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_353
timestamp 1667941163
transform 1 0 33580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_365
timestamp 1667941163
transform 1 0 34684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_377
timestamp 1667941163
transform 1 0 35788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1667941163
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_397
timestamp 1667941163
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1667941163
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1667941163
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1667941163
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_176
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_184
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1667941163
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_238
timestamp 1667941163
transform 1 0 23000 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1667941163
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1667941163
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1667941163
transform 1 0 29992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_328
timestamp 1667941163
transform 1 0 31280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_334
timestamp 1667941163
transform 1 0 31832 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_340
timestamp 1667941163
transform 1 0 32384 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_352
timestamp 1667941163
transform 1 0 33488 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1667941163
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1667941163
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1667941163
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1667941163
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1667941163
transform 1 0 15088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1667941163
transform 1 0 15732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1667941163
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1667941163
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1667941163
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_212
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1667941163
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_262
timestamp 1667941163
transform 1 0 25208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1667941163
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_292
timestamp 1667941163
transform 1 0 27968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_312
timestamp 1667941163
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_319
timestamp 1667941163
transform 1 0 30452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_326
timestamp 1667941163
transform 1 0 31096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1667941163
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_352
timestamp 1667941163
transform 1 0 33488 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_364
timestamp 1667941163
transform 1 0 34592 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_376
timestamp 1667941163
transform 1 0 35696 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1667941163
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1667941163
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_105
timestamp 1667941163
transform 1 0 10764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_120
timestamp 1667941163
transform 1 0 12144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1667941163
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1667941163
transform 1 0 13248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_152
timestamp 1667941163
transform 1 0 15088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1667941163
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1667941163
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_174
timestamp 1667941163
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1667941163
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_217
timestamp 1667941163
transform 1 0 21068 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_232
timestamp 1667941163
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1667941163
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_283
timestamp 1667941163
transform 1 0 27140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_293
timestamp 1667941163
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_314
timestamp 1667941163
transform 1 0 29992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_328
timestamp 1667941163
transform 1 0 31280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_334
timestamp 1667941163
transform 1 0 31832 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_340
timestamp 1667941163
transform 1 0 32384 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_352
timestamp 1667941163
transform 1 0 33488 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_121
timestamp 1667941163
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1667941163
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1667941163
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1667941163
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1667941163
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1667941163
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_179
timestamp 1667941163
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_207
timestamp 1667941163
transform 1 0 20148 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1667941163
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_235
timestamp 1667941163
transform 1 0 22724 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_241
timestamp 1667941163
transform 1 0 23276 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_264
timestamp 1667941163
transform 1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_292
timestamp 1667941163
transform 1 0 27968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_312
timestamp 1667941163
transform 1 0 29808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_319
timestamp 1667941163
transform 1 0 30452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_326
timestamp 1667941163
transform 1 0 31096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1667941163
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1667941163
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_73
timestamp 1667941163
transform 1 0 7820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1667941163
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_89
timestamp 1667941163
transform 1 0 9292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_101
timestamp 1667941163
transform 1 0 10396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1667941163
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1667941163
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_129
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_132
timestamp 1667941163
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1667941163
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1667941163
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_206
timestamp 1667941163
transform 1 0 20056 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_216
timestamp 1667941163
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1667941163
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1667941163
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_243
timestamp 1667941163
transform 1 0 23460 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1667941163
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_284
timestamp 1667941163
transform 1 0 27232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1667941163
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1667941163
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1667941163
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1667941163
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_143
timestamp 1667941163
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_150
timestamp 1667941163
transform 1 0 14904 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_156
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1667941163
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1667941163
transform 1 0 20700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1667941163
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_234
timestamp 1667941163
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_239
timestamp 1667941163
transform 1 0 23092 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1667941163
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1667941163
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_268
timestamp 1667941163
transform 1 0 25760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1667941163
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_303
timestamp 1667941163
transform 1 0 28980 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_310
timestamp 1667941163
transform 1 0 29624 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1667941163
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1667941163
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_110
timestamp 1667941163
transform 1 0 11224 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_122
timestamp 1667941163
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1667941163
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_147
timestamp 1667941163
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_150
timestamp 1667941163
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_156
timestamp 1667941163
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1667941163
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_176
timestamp 1667941163
transform 1 0 17296 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1667941163
transform 1 0 18308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1667941163
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_264
timestamp 1667941163
transform 1 0 25392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_271
timestamp 1667941163
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_279
timestamp 1667941163
transform 1 0 26772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1667941163
transform 1 0 28060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_300
timestamp 1667941163
transform 1 0 28704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1667941163
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_313
timestamp 1667941163
transform 1 0 29900 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_319
timestamp 1667941163
transform 1 0 30452 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_331
timestamp 1667941163
transform 1 0 31556 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_343
timestamp 1667941163
transform 1 0 32660 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_355
timestamp 1667941163
transform 1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1667941163
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_160
timestamp 1667941163
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_182
timestamp 1667941163
transform 1 0 17848 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_188
timestamp 1667941163
transform 1 0 18400 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1667941163
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1667941163
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1667941163
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1667941163
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_262
timestamp 1667941163
transform 1 0 25208 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_268
timestamp 1667941163
transform 1 0 25760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_303
timestamp 1667941163
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_309
timestamp 1667941163
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_321
timestamp 1667941163
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1667941163
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_397
timestamp 1667941163
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1667941163
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_33
timestamp 1667941163
transform 1 0 4140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_45
timestamp 1667941163
transform 1 0 5244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_57
timestamp 1667941163
transform 1 0 6348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_69
timestamp 1667941163
transform 1 0 7452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1667941163
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_132
timestamp 1667941163
transform 1 0 13248 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1667941163
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_171
timestamp 1667941163
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1667941163
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1667941163
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1667941163
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1667941163
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_206
timestamp 1667941163
transform 1 0 20056 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_264
timestamp 1667941163
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1667941163
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1667941163
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_297
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1667941163
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_186
timestamp 1667941163
transform 1 0 18216 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1667941163
transform 1 0 19136 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_211
timestamp 1667941163
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1667941163
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1667941163
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1667941163
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp 1667941163
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1667941163
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_299
timestamp 1667941163
transform 1 0 28612 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_397
timestamp 1667941163
transform 1 0 37628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1667941163
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1667941163
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_186
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1667941163
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_210
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_216
timestamp 1667941163
transform 1 0 20976 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp 1667941163
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_226
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_239
timestamp 1667941163
transform 1 0 23092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1667941163
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1667941163
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1667941163
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1667941163
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_292
timestamp 1667941163
transform 1 0 27968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_299
timestamp 1667941163
transform 1 0 28612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1667941163
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1667941163
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1667941163
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1667941163
transform 1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1667941163
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1667941163
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1667941163
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_254
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_269
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1667941163
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_298
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_310
timestamp 1667941163
transform 1 0 29624 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_322
timestamp 1667941163
transform 1 0 30728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1667941163
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_398
timestamp 1667941163
transform 1 0 37720 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1667941163
transform 1 0 38456 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp 1667941163
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1667941163
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_48
timestamp 1667941163
transform 1 0 5520 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_60
timestamp 1667941163
transform 1 0 6624 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_72
timestamp 1667941163
transform 1 0 7728 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_187
timestamp 1667941163
transform 1 0 18308 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1667941163
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_216
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_223
timestamp 1667941163
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_236
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_243
timestamp 1667941163
transform 1 0 23460 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_281
timestamp 1667941163
transform 1 0 26956 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_288
timestamp 1667941163
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1667941163
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_189
timestamp 1667941163
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1667941163
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1667941163
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1667941163
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_239
timestamp 1667941163
transform 1 0 23092 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_247
timestamp 1667941163
transform 1 0 23828 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1667941163
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_360
timestamp 1667941163
transform 1 0 34224 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_372
timestamp 1667941163
transform 1 0 35328 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1667941163
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_9
timestamp 1667941163
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1667941163
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1667941163
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_211
timestamp 1667941163
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_218
timestamp 1667941163
transform 1 0 21160 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_235
timestamp 1667941163
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_241
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_260
timestamp 1667941163
transform 1 0 25024 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_269
timestamp 1667941163
transform 1 0 25852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_281
timestamp 1667941163
transform 1 0 26956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_293
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1667941163
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1667941163
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_236
timestamp 1667941163
transform 1 0 22816 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_246
timestamp 1667941163
transform 1 0 23736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_256
timestamp 1667941163
transform 1 0 24656 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1667941163
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1667941163
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_10
timestamp 1667941163
transform 1 0 2024 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1667941163
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_68
timestamp 1667941163
transform 1 0 7360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_74
timestamp 1667941163
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1667941163
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1667941163
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_211
timestamp 1667941163
transform 1 0 20516 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_214
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1667941163
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_397
timestamp 1667941163
transform 1 0 37628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1667941163
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_210
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_9
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_21
timestamp 1667941163
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_33
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_45
timestamp 1667941163
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1667941163
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1667941163
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1667941163
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_267
timestamp 1667941163
transform 1 0 25668 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_271
timestamp 1667941163
transform 1 0 26036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1667941163
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1667941163
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_220
timestamp 1667941163
transform 1 0 21344 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_232
timestamp 1667941163
transform 1 0 22448 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1667941163
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_285
timestamp 1667941163
transform 1 0 27324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_291
timestamp 1667941163
transform 1 0 27876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1667941163
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1667941163
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_338
timestamp 1667941163
transform 1 0 32200 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_350
timestamp 1667941163
transform 1 0 33304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_10
timestamp 1667941163
transform 1 0 2024 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_16
timestamp 1667941163
transform 1 0 2576 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_28
timestamp 1667941163
transform 1 0 3680 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_40
timestamp 1667941163
transform 1 0 4784 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1667941163
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1667941163
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1667941163
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1667941163
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1667941163
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_208
timestamp 1667941163
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1667941163
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_397
timestamp 1667941163
transform 1 0 37628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 1667941163
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_323
timestamp 1667941163
transform 1 0 30820 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_335
timestamp 1667941163
transform 1 0 31924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_347
timestamp 1667941163
transform 1 0 33028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1667941163
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1667941163
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_397
timestamp 1667941163
transform 1 0 37628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1667941163
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_227
timestamp 1667941163
transform 1 0 21988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_239
timestamp 1667941163
transform 1 0 23092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1667941163
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1667941163
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_207
timestamp 1667941163
transform 1 0 20148 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_215
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_227
timestamp 1667941163
transform 1 0 21988 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_232
timestamp 1667941163
transform 1 0 22448 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_244
timestamp 1667941163
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_397
timestamp 1667941163
transform 1 0 37628 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_402
timestamp 1667941163
transform 1 0 38088 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1667941163
transform 1 0 38456 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_7
timestamp 1667941163
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1667941163
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1667941163
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1667941163
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1667941163
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_124
timestamp 1667941163
transform 1 0 12512 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_136
timestamp 1667941163
transform 1 0 13616 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_148
timestamp 1667941163
transform 1 0 14720 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1667941163
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1667941163
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1667941163
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_344
timestamp 1667941163
transform 1 0 32752 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_350
timestamp 1667941163
transform 1 0 33304 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_362
timestamp 1667941163
transform 1 0 34408 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1667941163
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1667941163
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_397
timestamp 1667941163
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_11
timestamp 1667941163
transform 1 0 2116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1667941163
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_16
timestamp 1667941163
transform 1 0 2576 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_22
timestamp 1667941163
transform 1 0 3128 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_34
timestamp 1667941163
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_46
timestamp 1667941163
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1667941163
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1667941163
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_230
timestamp 1667941163
transform 1 0 22264 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1667941163
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1667941163
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1667941163
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_320
timestamp 1667941163
transform 1 0 30544 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_332
timestamp 1667941163
transform 1 0 31648 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_344
timestamp 1667941163
transform 1 0 32752 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_356
timestamp 1667941163
transform 1 0 33856 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_397
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_402
timestamp 1667941163
transform 1 0 38088 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1667941163
transform 1 0 38456 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_385
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_17
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_101
timestamp 1667941163
transform 1 0 10396 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_135
timestamp 1667941163
transform 1 0 13524 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_147
timestamp 1667941163
transform 1 0 14628 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_159
timestamp 1667941163
transform 1 0 15732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_234
timestamp 1667941163
transform 1 0 22632 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_240
timestamp 1667941163
transform 1 0 23184 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_252
timestamp 1667941163
transform 1 0 24288 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_264
timestamp 1667941163
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1667941163
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_292
timestamp 1667941163
transform 1 0 27968 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_304
timestamp 1667941163
transform 1 0 29072 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_316
timestamp 1667941163
transform 1 0 30176 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 1667941163
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1667941163
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 1667941163
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_160
timestamp 1667941163
transform 1 0 15824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_261
timestamp 1667941163
transform 1 0 25116 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_317
timestamp 1667941163
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _213_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1667941163
transform -1 0 20976 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform 1 0 21160 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform -1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform -1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform 1 0 29532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform -1 0 16192 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform -1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform -1 0 26036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform -1 0 23736 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform -1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform -1 0 31096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform -1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform 1 0 31004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 24564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform -1 0 27968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform 1 0 28336 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform 1 0 30360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 27876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 25024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform 1 0 21068 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform 1 0 30176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 18952 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform -1 0 27324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 21160 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform -1 0 16376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform 1 0 14628 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform -1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform -1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform -1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 20240 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform 1 0 19872 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 14628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform -1 0 13248 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform 1 0 12880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 13248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform -1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform 1 0 31004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform -1 0 30452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 26496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 29072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform -1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform -1 0 28980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform -1 0 24104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform -1 0 26680 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform 1 0 27140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform -1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform -1 0 24472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform 1 0 14260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform -1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 28980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform 1 0 15272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 14628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform -1 0 17296 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform 1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform -1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform -1 0 29808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform -1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform -1 0 29624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform -1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform -1 0 30452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform -1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform -1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform -1 0 28704 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform -1 0 29992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform 1 0 19780 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform -1 0 31096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform 1 0 20976 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform 1 0 16100 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform -1 0 24472 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform 1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform 1 0 14168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform -1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform -1 0 18952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform -1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform -1 0 24840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform 1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform 1 0 30360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform -1 0 17204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 14168 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform -1 0 29992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform -1 0 16376 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform 1 0 17940 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform 1 0 18032 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform 1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform -1 0 20792 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform -1 0 2576 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform -1 0 21620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform 1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform 1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform 1 0 37444 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 30728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform -1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform -1 0 27416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform 1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform -1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform -1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform -1 0 30268 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform 1 0 20148 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform 1 0 26956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform 1 0 12972 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform -1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform -1 0 22264 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform 1 0 19596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform -1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform -1 0 27876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform 1 0 10396 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform -1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform 1 0 22632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 28520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform -1 0 30636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 33948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform 1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform -1 0 10488 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _380_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16652 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1667941163
transform -1 0 32200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform -1 0 32752 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform -1 0 11960 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform -1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform -1 0 29992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform -1 0 29808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform 1 0 14720 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _391_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _392_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform -1 0 35512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 36156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform -1 0 24104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform -1 0 24104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1667941163
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform -1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform -1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform 1 0 37812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform -1 0 32568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _403_
timestamp 1667941163
transform -1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform -1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform -1 0 33488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform -1 0 36340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform 1 0 32476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 30452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform -1 0 35696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _414_
timestamp 1667941163
transform -1 0 14996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform -1 0 27416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform 1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 36156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform -1 0 24104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1667941163
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform 1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform 1 0 17112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform -1 0 35512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _425_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14444 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform -1 0 37720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1667941163
transform -1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform -1 0 33212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform -1 0 35420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform -1 0 24104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform -1 0 37628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 36984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _436_
timestamp 1667941163
transform -1 0 18032 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform 1 0 15088 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform 1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform 1 0 14444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _447_
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform 1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform 1 0 14444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform 1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform 1 0 13616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform -1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform 1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _464_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1667941163
transform 1 0 27140 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _467_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23460 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _468_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _469_
timestamp 1667941163
transform -1 0 26680 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1667941163
transform -1 0 31188 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1667941163
transform 1 0 29716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _473_
timestamp 1667941163
transform 1 0 25944 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1667941163
transform -1 0 23920 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _475_
timestamp 1667941163
transform 1 0 26220 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1667941163
transform -1 0 28980 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1667941163
transform -1 0 31556 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1667941163
transform -1 0 34132 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _479_
timestamp 1667941163
transform -1 0 30084 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _480_
timestamp 1667941163
transform -1 0 31648 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _481_
timestamp 1667941163
transform 1 0 24656 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1667941163
transform 1 0 21252 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _485_
timestamp 1667941163
transform -1 0 25944 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _486_
timestamp 1667941163
transform -1 0 28796 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _487_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1667941163
transform -1 0 24748 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1667941163
transform -1 0 26404 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1667941163
transform -1 0 21528 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _491_
timestamp 1667941163
transform 1 0 21344 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _492_
timestamp 1667941163
transform -1 0 24104 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _493_
timestamp 1667941163
transform -1 0 31740 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1667941163
transform 1 0 31924 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1667941163
transform 1 0 28244 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _497_
timestamp 1667941163
transform 1 0 27784 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1667941163
transform -1 0 31648 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _499_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1667941163
transform -1 0 28888 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1667941163
transform 1 0 29716 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _503_
timestamp 1667941163
transform -1 0 23184 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1667941163
transform -1 0 26496 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _505_
timestamp 1667941163
transform -1 0 29992 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1667941163
transform -1 0 28612 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1667941163
transform -1 0 21528 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1667941163
transform -1 0 26128 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _509_
timestamp 1667941163
transform -1 0 26772 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _510_
timestamp 1667941163
transform -1 0 29256 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _511_
timestamp 1667941163
transform -1 0 26680 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1667941163
transform -1 0 26680 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1667941163
transform 1 0 27968 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _515_
timestamp 1667941163
transform 1 0 24288 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _516_
timestamp 1667941163
transform -1 0 23460 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _517_
timestamp 1667941163
transform -1 0 23920 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _518_
timestamp 1667941163
transform -1 0 26588 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1667941163
transform 1 0 19688 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _521_
timestamp 1667941163
transform -1 0 23920 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _522_
timestamp 1667941163
transform -1 0 23920 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _523_
timestamp 1667941163
transform -1 0 27232 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform -1 0 26404 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1667941163
transform -1 0 23828 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp 1667941163
transform 1 0 21620 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1667941163
transform -1 0 23000 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _529_
timestamp 1667941163
transform -1 0 29808 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10488 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _542_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21436 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1667941163
transform -1 0 20240 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _544_
timestamp 1667941163
transform -1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1667941163
transform -1 0 36984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _546_
timestamp 1667941163
transform 1 0 20516 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1667941163
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1667941163
transform -1 0 29992 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1667941163
transform -1 0 38088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _550_
timestamp 1667941163
transform 1 0 12696 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1667941163
transform 1 0 11500 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1667941163
transform -1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1667941163
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1667941163
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1667941163
transform -1 0 38088 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1667941163
transform 1 0 1748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _559_
timestamp 1667941163
transform -1 0 21712 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1667941163
transform -1 0 37444 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1667941163
transform -1 0 19688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1667941163
transform -1 0 31832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1667941163
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform 1 0 33212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _565_
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _566_
timestamp 1667941163
transform -1 0 23092 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _567_
timestamp 1667941163
transform 1 0 19136 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1667941163
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform -1 0 26036 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _570_
timestamp 1667941163
transform -1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform -1 0 27968 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1667941163
transform -1 0 22632 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _575_
timestamp 1667941163
transform -1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1667941163
transform -1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1667941163
transform -1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21252 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _580_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _581_
timestamp 1667941163
transform -1 0 20148 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _582_
timestamp 1667941163
transform 1 0 17848 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _583__91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 15088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _583_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _584_
timestamp 1667941163
transform -1 0 25392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18768 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _586_
timestamp 1667941163
transform -1 0 19320 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _587_
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _588_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1667941163
transform 1 0 16652 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _590_
timestamp 1667941163
transform -1 0 21068 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _591_
timestamp 1667941163
transform 1 0 28336 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _592_
timestamp 1667941163
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _592__92
timestamp 1667941163
transform -1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _593_
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1667941163
transform 1 0 28336 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _595_
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _596_
timestamp 1667941163
transform 1 0 19780 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _597_
timestamp 1667941163
transform -1 0 28428 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _598_
timestamp 1667941163
transform 1 0 18676 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _599_
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _600_
timestamp 1667941163
transform 1 0 15272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _601_
timestamp 1667941163
transform -1 0 23460 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _602_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _603_
timestamp 1667941163
transform -1 0 18584 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _604_
timestamp 1667941163
transform -1 0 19780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _605_
timestamp 1667941163
transform 1 0 19320 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _606__93
timestamp 1667941163
transform 1 0 27600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _606_
timestamp 1667941163
transform -1 0 24196 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _607_
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _608_
timestamp 1667941163
transform -1 0 25392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _609_
timestamp 1667941163
transform -1 0 26772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _610_
timestamp 1667941163
transform -1 0 26680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _611_
timestamp 1667941163
transform -1 0 20240 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _612_
timestamp 1667941163
transform -1 0 27784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _613_
timestamp 1667941163
transform -1 0 25392 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _614_
timestamp 1667941163
transform -1 0 26588 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _615_
timestamp 1667941163
transform -1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _616_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _617_
timestamp 1667941163
transform 1 0 17020 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _618__94
timestamp 1667941163
transform 1 0 19596 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _618_
timestamp 1667941163
transform 1 0 19412 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _619_
timestamp 1667941163
transform -1 0 21436 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _620_
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _621_
timestamp 1667941163
transform -1 0 24656 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _622_
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _623_
timestamp 1667941163
transform -1 0 20240 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _624_
timestamp 1667941163
transform 1 0 21988 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _625_
timestamp 1667941163
transform 1 0 18768 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _626_
timestamp 1667941163
transform -1 0 27968 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _627_
timestamp 1667941163
transform 1 0 16560 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _628_
timestamp 1667941163
transform 1 0 15364 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _629_
timestamp 1667941163
transform 1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _630__95
timestamp 1667941163
transform 1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _630_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _631_
timestamp 1667941163
transform 1 0 15548 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _632_
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform -1 0 17664 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform -1 0 29072 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _635_
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform -1 0 24012 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform -1 0 27968 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _638_
timestamp 1667941163
transform -1 0 26312 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _639_
timestamp 1667941163
transform 1 0 27232 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform -1 0 27968 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _642__96
timestamp 1667941163
transform -1 0 24104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _643_
timestamp 1667941163
transform 1 0 20516 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _644_
timestamp 1667941163
transform 1 0 20424 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform -1 0 26588 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _647_
timestamp 1667941163
transform 1 0 28336 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _649_
timestamp 1667941163
transform 1 0 18676 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform -1 0 27968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _651_
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _652_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _653_
timestamp 1667941163
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _654_
timestamp 1667941163
transform 1 0 14536 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _654__97
timestamp 1667941163
transform -1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _655_
timestamp 1667941163
transform 1 0 16928 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _656_
timestamp 1667941163
transform -1 0 24012 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform 1 0 18124 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform -1 0 22448 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _659_
timestamp 1667941163
transform -1 0 19872 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _660_
timestamp 1667941163
transform 1 0 15548 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _661_
timestamp 1667941163
transform 1 0 17572 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _662_
timestamp 1667941163
transform 1 0 20148 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform 1 0 16928 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _665_
timestamp 1667941163
transform -1 0 24012 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform -1 0 23460 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _666__98
timestamp 1667941163
transform 1 0 23368 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _667_
timestamp 1667941163
transform -1 0 25208 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _668_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _669_
timestamp 1667941163
transform -1 0 21528 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform 1 0 18124 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform -1 0 18676 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform 1 0 17020 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _673_
timestamp 1667941163
transform -1 0 21620 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _675_
timestamp 1667941163
transform 1 0 26864 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _676_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _678__99
timestamp 1667941163
transform 1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform -1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _679_
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _680_
timestamp 1667941163
transform -1 0 25208 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _681_
timestamp 1667941163
transform -1 0 26680 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _683_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform -1 0 26588 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _685_
timestamp 1667941163
transform 1 0 18124 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _687_
timestamp 1667941163
transform -1 0 25760 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _688_
timestamp 1667941163
transform 1 0 22632 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform 1 0 18308 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _690__100
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 20148 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform 1 0 21896 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform -1 0 25392 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _695_
timestamp 1667941163
transform -1 0 25116 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform -1 0 23644 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform -1 0 26036 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform -1 0 17020 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _700__101
timestamp 1667941163
transform -1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform 1 0 17480 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform 1 0 18124 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform 1 0 20976 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _704_
timestamp 1667941163
transform -1 0 23644 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _705_
timestamp 1667941163
transform -1 0 19780 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform -1 0 26404 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform -1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform -1 0 35972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform -1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform 1 0 37444 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 35512 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform -1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform -1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform -1 0 38364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform 1 0 37444 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1667941163
transform -1 0 38364 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform -1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform -1 0 38364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform -1 0 38364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1667941163
transform -1 0 38364 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform -1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform -1 0 26128 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform -1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 38088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 30452 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1667941163
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform -1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 25208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform -1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform -1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform -1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 24104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform -1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 6900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 13340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform -1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform -1 0 3036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 12 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 13 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 14 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 15 nsew signal input
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 16 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 17 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 18 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 19 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 20 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 21 nsew signal tristate
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 22 nsew signal tristate
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 23 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 24 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 26 nsew signal tristate
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_bottom_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 28 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_bottom_out[17]
port 29 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 30 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 31 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 32 nsew signal tristate
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 33 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 34 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 35 nsew signal tristate
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 36 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 37 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 38 nsew signal tristate
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
port 78 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
port 79 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
port 80 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
port 81 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_
port 82 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_
port 83 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_
port 84 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_
port 85 nsew signal tristate
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 pReset
port 86 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 prog_clk
port 87 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 88 nsew signal tristate
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 89 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 90 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 31241 4590 31241 4590 0 _000_
rlabel metal1 28711 5610 28711 5610 0 _001_
rlabel metal1 21259 6698 21259 6698 0 _002_
rlabel metal2 22034 9044 22034 9044 0 _003_
rlabel metal1 24610 6630 24610 6630 0 _004_
rlabel metal2 15318 2176 15318 2176 0 _005_
rlabel metal2 36294 4318 36294 4318 0 _006_
rlabel metal1 37168 3978 37168 3978 0 _007_
rlabel metal1 34822 7956 34822 7956 0 _008_
rlabel metal1 27370 11159 27370 11159 0 _009_
rlabel metal2 20838 9911 20838 9911 0 _010_
rlabel metal1 28205 6698 28205 6698 0 _011_
rlabel metal2 32890 4624 32890 4624 0 _012_
rlabel metal1 30130 2455 30130 2455 0 _013_
rlabel metal1 32706 4998 32706 4998 0 _014_
rlabel metal1 27370 7242 27370 7242 0 _015_
rlabel metal1 30498 8534 30498 8534 0 _016_
rlabel metal1 27830 2312 27830 2312 0 _017_
rlabel metal1 33817 3434 33817 3434 0 _018_
rlabel metal1 29309 2414 29309 2414 0 _019_
rlabel metal1 23237 3502 23237 3502 0 _020_
rlabel metal1 26450 8602 26450 8602 0 _021_
rlabel metal2 25530 7820 25530 7820 0 _022_
rlabel metal1 33879 6358 33879 6358 0 _023_
rlabel metal2 23966 4318 23966 4318 0 _024_
rlabel metal1 20792 5270 20792 5270 0 _025_
rlabel metal1 18630 5882 18630 5882 0 _026_
rlabel metal2 13754 9248 13754 9248 0 _027_
rlabel metal2 20194 7752 20194 7752 0 _028_
rlabel metal2 31832 3638 31832 3638 0 _029_
rlabel metal1 33679 5678 33679 5678 0 _030_
rlabel metal1 34178 5576 34178 5576 0 _031_
rlabel metal1 34822 8806 34822 8806 0 _032_
rlabel metal1 29447 8534 29447 8534 0 _033_
rlabel metal1 33258 9928 33258 9928 0 _034_
rlabel metal1 23644 5542 23644 5542 0 _035_
rlabel metal1 37444 3638 37444 3638 0 _036_
rlabel metal1 31609 3434 31609 3434 0 _037_
rlabel metal1 22080 4998 22080 4998 0 _038_
rlabel metal2 19642 7293 19642 7293 0 _039_
rlabel metal1 13708 5882 13708 5882 0 _040_
rlabel metal1 15318 6766 15318 6766 0 _041_
rlabel metal2 18170 3808 18170 3808 0 _042_
rlabel metal2 18814 3145 18814 3145 0 _043_
rlabel metal1 16376 4794 16376 4794 0 _044_
rlabel metal1 22126 7956 22126 7956 0 _045_
rlabel metal2 19550 7412 19550 7412 0 _046_
rlabel via2 17066 6715 17066 6715 0 _047_
rlabel metal1 15824 7378 15824 7378 0 _048_
rlabel metal1 16054 7922 16054 7922 0 _049_
rlabel metal1 15824 6426 15824 6426 0 _050_
rlabel metal1 13662 6970 13662 6970 0 _051_
rlabel metal2 20516 5134 20516 5134 0 _052_
rlabel metal2 20470 5916 20470 5916 0 _053_
rlabel metal2 27278 6936 27278 6936 0 _054_
rlabel via2 16238 5627 16238 5627 0 _055_
rlabel metal1 13846 6426 13846 6426 0 _056_
rlabel metal1 12512 6426 12512 6426 0 _057_
rlabel metal1 20194 6222 20194 6222 0 _058_
rlabel metal1 16054 6834 16054 6834 0 _059_
rlabel metal1 12259 3706 12259 3706 0 _060_
rlabel metal2 15226 5457 15226 5457 0 _061_
rlabel metal1 12834 8840 12834 8840 0 _062_
rlabel metal2 18170 7888 18170 7888 0 _063_
rlabel metal1 12788 7174 12788 7174 0 _064_
rlabel metal2 19182 6919 19182 6919 0 _065_
rlabel metal1 15180 4114 15180 4114 0 _066_
rlabel metal1 12351 2958 12351 2958 0 _067_
rlabel metal2 19734 8976 19734 8976 0 _068_
rlabel metal1 20930 5202 20930 5202 0 _069_
rlabel metal2 33166 7854 33166 7854 0 _070_
rlabel metal1 15502 4148 15502 4148 0 _071_
rlabel via2 21942 4811 21942 4811 0 _072_
rlabel metal2 21022 16558 21022 16558 0 _073_
rlabel metal2 21390 14688 21390 14688 0 _074_
rlabel metal1 19688 15538 19688 15538 0 _075_
rlabel metal1 17572 14450 17572 14450 0 _076_
rlabel metal1 16468 14790 16468 14790 0 _077_
rlabel via2 27738 12053 27738 12053 0 _078_
rlabel metal1 18998 11832 18998 11832 0 _079_
rlabel metal1 18952 8058 18952 8058 0 _080_
rlabel metal2 20102 13668 20102 13668 0 _081_
rlabel via2 17066 13923 17066 13923 0 _082_
rlabel metal2 16882 11696 16882 11696 0 _083_
rlabel metal1 20792 13226 20792 13226 0 _084_
rlabel metal1 31326 13838 31326 13838 0 _085_
rlabel metal1 19826 11016 19826 11016 0 _086_
rlabel metal1 15088 11798 15088 11798 0 _087_
rlabel metal1 29210 12886 29210 12886 0 _088_
rlabel metal1 24104 11866 24104 11866 0 _089_
rlabel metal2 18998 12240 18998 12240 0 _090_
rlabel metal1 28198 9928 28198 9928 0 _091_
rlabel metal1 17158 10710 17158 10710 0 _092_
rlabel via2 30958 11747 30958 11747 0 _093_
rlabel metal1 14904 12682 14904 12682 0 _094_
rlabel metal1 23690 9622 23690 9622 0 _095_
rlabel metal1 21666 12886 21666 12886 0 _096_
rlabel metal2 18308 4114 18308 4114 0 _097_
rlabel metal1 18354 4794 18354 4794 0 _098_
rlabel metal2 19550 14824 19550 14824 0 _099_
rlabel metal1 24334 13974 24334 13974 0 _100_
rlabel metal1 21896 15402 21896 15402 0 _101_
rlabel metal2 27462 12716 27462 12716 0 _102_
rlabel metal1 26542 13192 26542 13192 0 _103_
rlabel metal2 26450 16592 26450 16592 0 _104_
rlabel metal1 20148 6426 20148 6426 0 _105_
rlabel metal1 29118 12648 29118 12648 0 _106_
rlabel viali 25165 15402 25165 15402 0 _107_
rlabel metal2 29670 13124 29670 13124 0 _108_
rlabel metal1 14168 7514 14168 7514 0 _109_
rlabel metal1 16652 5270 16652 5270 0 _110_
rlabel metal2 17158 15912 17158 15912 0 _111_
rlabel metal2 19458 18462 19458 18462 0 _112_
rlabel metal1 19918 16150 19918 16150 0 _113_
rlabel metal1 20240 18938 20240 18938 0 _114_
rlabel metal1 25760 14586 25760 14586 0 _115_
rlabel metal1 26082 18666 26082 18666 0 _116_
rlabel metal1 20378 9078 20378 9078 0 _117_
rlabel metal1 22172 18394 22172 18394 0 _118_
rlabel metal1 20654 18394 20654 18394 0 _119_
rlabel metal1 27646 18326 27646 18326 0 _120_
rlabel metal1 16698 6834 16698 6834 0 _121_
rlabel metal2 15594 7378 15594 7378 0 _122_
rlabel metal1 15088 9622 15088 9622 0 _123_
rlabel metal1 14490 13192 14490 13192 0 _124_
rlabel metal2 15778 14042 15778 14042 0 _125_
rlabel metal2 17986 10047 17986 10047 0 _126_
rlabel metal1 16422 16558 16422 16558 0 _127_
rlabel metal1 27416 9622 27416 9622 0 _128_
rlabel metal1 16468 7446 16468 7446 0 _129_
rlabel metal2 23782 17646 23782 17646 0 _130_
rlabel metal2 27738 14382 27738 14382 0 _131_
rlabel metal1 26312 17850 26312 17850 0 _132_
rlabel metal1 27554 13226 27554 13226 0 _133_
rlabel metal1 28796 13226 28796 13226 0 _134_
rlabel metal1 28382 12954 28382 12954 0 _135_
rlabel metal2 22586 13056 22586 13056 0 _136_
rlabel metal2 23414 14110 23414 14110 0 _137_
rlabel metal2 20654 16728 20654 16728 0 _138_
rlabel metal2 28106 14331 28106 14331 0 _139_
rlabel metal2 23506 16354 23506 16354 0 _140_
rlabel metal1 28566 11832 28566 11832 0 _141_
rlabel metal1 16330 12886 16330 12886 0 _142_
rlabel metal1 18906 12920 18906 12920 0 _143_
rlabel metal1 28014 11798 28014 11798 0 _144_
rlabel metal1 17894 6834 17894 6834 0 _145_
rlabel metal1 13294 6426 13294 6426 0 _146_
rlabel metal1 15502 10642 15502 10642 0 _147_
rlabel metal1 14214 10642 14214 10642 0 _148_
rlabel metal1 15732 8602 15732 8602 0 _149_
rlabel metal1 23046 12886 23046 12886 0 _150_
rlabel metal1 18354 12104 18354 12104 0 _151_
rlabel metal2 22126 13634 22126 13634 0 _152_
rlabel metal2 20746 8296 20746 8296 0 _153_
rlabel metal1 13616 12682 13616 12682 0 _154_
rlabel metal1 16100 11322 16100 11322 0 _155_
rlabel metal1 17480 13498 17480 13498 0 _156_
rlabel metal1 15502 5338 15502 5338 0 _157_
rlabel metal1 16698 3706 16698 3706 0 _158_
rlabel metal1 23782 16184 23782 16184 0 _159_
rlabel metal1 23230 14280 23230 14280 0 _160_
rlabel metal2 24978 17374 24978 17374 0 _161_
rlabel metal1 16928 15062 16928 15062 0 _162_
rlabel metal1 23184 9146 23184 9146 0 _163_
rlabel metal1 16744 8602 16744 8602 0 _164_
rlabel metal1 17158 3910 17158 3910 0 _165_
rlabel metal1 17756 3094 17756 3094 0 _166_
rlabel metal1 20608 8602 20608 8602 0 _167_
rlabel metal1 19642 8840 19642 8840 0 _168_
rlabel metal1 30268 14042 30268 14042 0 _169_
rlabel metal2 28750 14212 28750 14212 0 _170_
rlabel metal2 21206 17374 21206 17374 0 _171_
rlabel metal2 25622 19006 25622 19006 0 _172_
rlabel metal2 21942 16763 21942 16763 0 _173_
rlabel metal1 25622 16150 25622 16150 0 _174_
rlabel metal1 26450 15096 26450 15096 0 _175_
rlabel metal1 26312 16490 26312 16490 0 _176_
rlabel via2 31142 13515 31142 13515 0 _177_
rlabel metal1 26312 14314 26312 14314 0 _178_
rlabel metal1 18446 15062 18446 15062 0 _179_
rlabel metal2 24794 13464 24794 13464 0 _180_
rlabel metal2 30958 15946 30958 15946 0 _181_
rlabel metal1 25852 15674 25852 15674 0 _182_
rlabel metal2 18538 17374 18538 17374 0 _183_
rlabel metal1 20562 18666 20562 18666 0 _184_
rlabel metal2 22494 17102 22494 17102 0 _185_
rlabel metal2 22126 19346 22126 19346 0 _186_
rlabel metal2 25162 16728 25162 16728 0 _187_
rlabel metal2 22494 19822 22494 19822 0 _188_
rlabel metal1 25392 19414 25392 19414 0 _189_
rlabel metal1 22494 17544 22494 17544 0 _190_
rlabel metal2 23414 17544 23414 17544 0 _191_
rlabel metal1 25806 17544 25806 17544 0 _192_
rlabel metal1 15686 7514 15686 7514 0 _193_
rlabel via2 16974 5355 16974 5355 0 _194_
rlabel metal1 17894 13226 17894 13226 0 _195_
rlabel metal2 18354 9758 18354 9758 0 _196_
rlabel metal1 20838 12682 20838 12682 0 _197_
rlabel metal2 21298 12036 21298 12036 0 _198_
rlabel metal1 18262 6698 18262 6698 0 _199_
rlabel metal1 29210 12750 29210 12750 0 _200_
rlabel metal2 20838 10472 20838 10472 0 _201_
rlabel via2 1610 3485 1610 3485 0 ccff_head
rlabel metal1 37536 36890 37536 36890 0 ccff_tail
rlabel via2 1610 17765 1610 17765 0 chany_bottom_in[0]
rlabel metal1 35788 2414 35788 2414 0 chany_bottom_in[10]
rlabel metal1 14904 37298 14904 37298 0 chany_bottom_in[11]
rlabel metal2 16698 37383 16698 37383 0 chany_bottom_in[12]
rlabel metal1 17894 37434 17894 37434 0 chany_bottom_in[13]
rlabel metal1 14214 2414 14214 2414 0 chany_bottom_in[14]
rlabel metal1 37352 8398 37352 8398 0 chany_bottom_in[15]
rlabel metal1 35512 37298 35512 37298 0 chany_bottom_in[16]
rlabel metal1 21988 37298 21988 37298 0 chany_bottom_in[17]
rlabel metal2 13570 1520 13570 1520 0 chany_bottom_in[18]
rlabel metal2 38226 11679 38226 11679 0 chany_bottom_in[1]
rlabel metal2 38226 17119 38226 17119 0 chany_bottom_in[2]
rlabel metal2 37490 35513 37490 35513 0 chany_bottom_in[3]
rlabel via2 38318 32011 38318 32011 0 chany_bottom_in[4]
rlabel metal1 37444 5202 37444 5202 0 chany_bottom_in[5]
rlabel via2 1610 28645 1610 28645 0 chany_bottom_in[6]
rlabel metal1 8464 2278 8464 2278 0 chany_bottom_in[7]
rlabel metal2 38226 26775 38226 26775 0 chany_bottom_in[8]
rlabel via2 1702 30651 1702 30651 0 chany_bottom_in[9]
rlabel metal3 1188 14348 1188 14348 0 chany_bottom_out[0]
rlabel via2 38226 27931 38226 27931 0 chany_bottom_out[10]
rlabel metal2 37398 1520 37398 1520 0 chany_bottom_out[11]
rlabel metal1 25300 37094 25300 37094 0 chany_bottom_out[12]
rlabel metal1 1518 37094 1518 37094 0 chany_bottom_out[13]
rlabel via2 38226 30005 38226 30005 0 chany_bottom_out[14]
rlabel metal3 1188 19788 1188 19788 0 chany_bottom_out[15]
rlabel metal3 1188 23188 1188 23188 0 chany_bottom_out[16]
rlabel metal3 1188 1428 1188 1428 0 chany_bottom_out[17]
rlabel metal2 30314 1520 30314 1520 0 chany_bottom_out[18]
rlabel metal3 1188 34068 1188 34068 0 chany_bottom_out[1]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[2]
rlabel metal1 28520 37094 28520 37094 0 chany_bottom_out[3]
rlabel metal1 34408 2822 34408 2822 0 chany_bottom_out[4]
rlabel metal1 20102 37094 20102 37094 0 chany_bottom_out[5]
rlabel via2 38226 33371 38226 33371 0 chany_bottom_out[6]
rlabel metal2 23874 2064 23874 2064 0 chany_bottom_out[7]
rlabel metal3 1188 21148 1188 21148 0 chany_bottom_out[8]
rlabel metal1 37030 2278 37030 2278 0 chany_bottom_out[9]
rlabel metal2 38226 15895 38226 15895 0 chany_top_in[0]
rlabel metal1 2346 36754 2346 36754 0 chany_top_in[10]
rlabel via2 1610 10251 1610 10251 0 chany_top_in[11]
rlabel via2 1610 32011 1610 32011 0 chany_top_in[12]
rlabel metal3 1142 6868 1142 6868 0 chany_top_in[13]
rlabel metal2 38318 37383 38318 37383 0 chany_top_in[14]
rlabel metal1 7866 37230 7866 37230 0 chany_top_in[15]
rlabel metal1 3312 2278 3312 2278 0 chany_top_in[16]
rlabel metal1 9798 2414 9798 2414 0 chany_top_in[17]
rlabel metal2 32246 1761 32246 1761 0 chany_top_in[18]
rlabel metal2 38318 13583 38318 13583 0 chany_top_in[1]
rlabel metal2 38226 6239 38226 6239 0 chany_top_in[2]
rlabel metal2 33902 3808 33902 3808 0 chany_top_in[3]
rlabel metal1 2668 36822 2668 36822 0 chany_top_in[4]
rlabel metal1 38272 3502 38272 3502 0 chany_top_in[5]
rlabel via2 1610 8925 1610 8925 0 chany_top_in[6]
rlabel metal2 38318 10455 38318 10455 0 chany_top_in[7]
rlabel via2 1610 25245 1610 25245 0 chany_top_in[8]
rlabel metal2 34086 6018 34086 6018 0 chany_top_in[9]
rlabel via2 38226 24565 38226 24565 0 chany_top_out[0]
rlabel metal1 11730 37094 11730 37094 0 chany_top_out[10]
rlabel metal1 6578 37094 6578 37094 0 chany_top_out[11]
rlabel metal2 18722 1520 18722 1520 0 chany_top_out[12]
rlabel metal2 46 1656 46 1656 0 chany_top_out[13]
rlabel metal2 21942 1435 21942 1435 0 chany_top_out[14]
rlabel metal1 13018 37094 13018 37094 0 chany_top_out[15]
rlabel metal1 23368 37094 23368 37094 0 chany_top_out[16]
rlabel metal1 33672 37094 33672 37094 0 chany_top_out[17]
rlabel metal3 1188 26588 1188 26588 0 chany_top_out[18]
rlabel metal2 4554 1520 4554 1520 0 chany_top_out[1]
rlabel metal2 1334 1520 1334 1520 0 chany_top_out[2]
rlabel metal1 38456 36346 38456 36346 0 chany_top_out[3]
rlabel metal1 30498 37094 30498 37094 0 chany_top_out[4]
rlabel metal2 16790 1520 16790 1520 0 chany_top_out[5]
rlabel metal1 37352 36346 37352 36346 0 chany_top_out[6]
rlabel metal1 38272 2822 38272 2822 0 chany_top_out[7]
rlabel metal1 4692 37094 4692 37094 0 chany_top_out[8]
rlabel metal2 38226 21233 38226 21233 0 chany_top_out[9]
rlabel metal2 6486 1520 6486 1520 0 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 11638 1520 11638 1520 0 left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal3 1188 15708 1188 15708 0 left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel via2 38226 22491 38226 22491 0 left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20148 3366 20148 3366 0 left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal3 1188 4828 1188 4828 0 left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal1 32338 37094 32338 37094 0 left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_
rlabel metal2 2806 37145 2806 37145 0 left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_
rlabel metal1 19090 4590 19090 4590 0 mem_left_ipin_0.DFFR_0_.Q
rlabel metal2 18078 15572 18078 15572 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal1 19366 17646 19366 17646 0 mem_left_ipin_0.DFFR_2_.Q
rlabel metal1 20976 6902 20976 6902 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal2 28934 5933 28934 5933 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal3 19458 7820 19458 7820 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal1 21114 12818 21114 12818 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal1 16284 12818 16284 12818 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal2 18906 11322 18906 11322 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal1 31372 7990 31372 7990 0 mem_left_ipin_1.DFFR_3_.Q
rlabel metal1 33856 3162 33856 3162 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal2 29900 12716 29900 12716 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal2 20930 9860 20930 9860 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal1 17250 12818 17250 12818 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal1 23460 11798 23460 11798 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal2 21758 7242 21758 7242 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal2 15042 7174 15042 7174 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal1 19550 4216 19550 4216 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal1 27048 2278 27048 2278 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal1 29302 14994 29302 14994 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal1 36501 2550 36501 2550 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal1 31188 2346 31188 2346 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal1 29348 2482 29348 2482 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal1 21298 4488 21298 4488 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal1 20838 18292 20838 18292 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal1 18538 15980 18538 15980 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal1 19550 18802 19550 18802 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal1 24794 2516 24794 2516 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal1 28796 2618 28796 2618 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal2 20010 4658 20010 4658 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal1 24472 20230 24472 20230 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal1 14030 14790 14030 14790 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal1 22655 1870 22655 1870 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal1 16376 7378 16376 7378 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal2 16974 6596 16974 6596 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal1 21390 3944 21390 3944 0 mem_right_ipin_2.DFFR_5_.Q
rlabel metal2 15502 13158 15502 13158 0 mem_right_ipin_3.DFFR_0_.Q
rlabel metal1 30498 14382 30498 14382 0 mem_right_ipin_3.DFFR_1_.Q
rlabel metal1 18722 13328 18722 13328 0 mem_right_ipin_3.DFFR_2_.Q
rlabel metal1 30544 5746 30544 5746 0 mem_right_ipin_3.DFFR_3_.Q
rlabel metal1 30176 16082 30176 16082 0 mem_right_ipin_3.DFFR_4_.Q
rlabel metal1 29854 9622 29854 9622 0 mem_right_ipin_3.DFFR_5_.Q
rlabel metal1 17020 13294 17020 13294 0 mem_right_ipin_4.DFFR_0_.Q
rlabel metal1 15502 8432 15502 8432 0 mem_right_ipin_4.DFFR_1_.Q
rlabel metal1 17112 1870 17112 1870 0 mem_right_ipin_4.DFFR_2_.Q
rlabel metal1 30038 3400 30038 3400 0 mem_right_ipin_4.DFFR_3_.Q
rlabel metal2 17894 5729 17894 5729 0 mem_right_ipin_4.DFFR_4_.Q
rlabel metal1 25576 6222 25576 6222 0 mem_right_ipin_4.DFFR_5_.Q
rlabel metal1 14720 10030 14720 10030 0 mem_right_ipin_5.DFFR_0_.Q
rlabel metal1 24472 17646 24472 17646 0 mem_right_ipin_5.DFFR_1_.Q
rlabel metal2 16422 15674 16422 15674 0 mem_right_ipin_5.DFFR_2_.Q
rlabel metal1 22034 2958 22034 2958 0 mem_right_ipin_5.DFFR_3_.Q
rlabel metal1 19596 2822 19596 2822 0 mem_right_ipin_5.DFFR_4_.Q
rlabel via2 21666 3587 21666 3587 0 mem_right_ipin_5.DFFR_5_.Q
rlabel metal1 18906 15436 18906 15436 0 mem_right_ipin_6.DFFR_0_.Q
rlabel metal1 21804 8058 21804 8058 0 mem_right_ipin_6.DFFR_1_.Q
rlabel metal1 27094 17646 27094 17646 0 mem_right_ipin_6.DFFR_2_.Q
rlabel metal1 30912 13294 30912 13294 0 mem_right_ipin_6.DFFR_3_.Q
rlabel metal1 29854 13974 29854 13974 0 mem_right_ipin_6.DFFR_4_.Q
rlabel metal1 27508 10778 27508 10778 0 mem_right_ipin_6.DFFR_5_.Q
rlabel metal1 23828 17646 23828 17646 0 mem_right_ipin_7.DFFR_0_.Q
rlabel metal1 21344 18258 21344 18258 0 mem_right_ipin_7.DFFR_1_.Q
rlabel metal2 21114 20128 21114 20128 0 mem_right_ipin_7.DFFR_2_.Q
rlabel metal1 26680 9554 26680 9554 0 mem_right_ipin_7.DFFR_3_.Q
rlabel metal1 31142 12818 31142 12818 0 mem_right_ipin_7.DFFR_4_.Q
rlabel metal2 20286 13532 20286 13532 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal2 18354 14076 18354 14076 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 22080 21318 22080 21318 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal2 16882 13991 16882 13991 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal1 19734 14382 19734 14382 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 20608 25126 20608 25126 0 mux_left_ipin_0.INVTX1_5_.out
rlabel metal1 17204 12750 17204 12750 0 mux_left_ipin_0.INVTX1_6_.out
rlabel metal2 30222 12886 30222 12886 0 mux_left_ipin_0.INVTX1_7_.out
rlabel metal1 21022 13226 21022 13226 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 19182 14654 19182 14654 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 18952 11662 18952 11662 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 2806 34578 2806 34578 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 20516 10574 20516 10574 0 mux_left_ipin_1.INVTX1_2_.out
rlabel metal1 23276 9486 23276 9486 0 mux_left_ipin_1.INVTX1_3_.out
rlabel metal1 18584 10574 18584 10574 0 mux_left_ipin_1.INVTX1_4_.out
rlabel metal1 24012 12750 24012 12750 0 mux_left_ipin_1.INVTX1_5_.out
rlabel metal1 14582 12138 14582 12138 0 mux_left_ipin_1.INVTX1_6_.out
rlabel metal1 15686 10540 15686 10540 0 mux_left_ipin_1.INVTX1_7_.out
rlabel metal1 24426 12342 24426 12342 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20838 10506 20838 10506 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 21114 13498 21114 13498 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 28934 16048 28934 16048 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27002 12954 27002 12954 0 mux_left_ipin_2.INVTX1_2_.out
rlabel metal1 26956 14926 26956 14926 0 mux_left_ipin_2.INVTX1_3_.out
rlabel metal1 16100 27846 16100 27846 0 mux_left_ipin_2.INVTX1_4_.out
rlabel metal1 18078 9486 18078 9486 0 mux_left_ipin_2.INVTX1_5_.out
rlabel metal2 20286 8993 20286 8993 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16882 7956 16882 7956 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15410 7786 15410 7786 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 29256 27302 29256 27302 0 mux_right_ipin_0.INVTX1_2_.out
rlabel metal1 25898 16626 25898 16626 0 mux_right_ipin_0.INVTX1_3_.out
rlabel metal2 21758 17918 21758 17918 0 mux_right_ipin_0.INVTX1_4_.out
rlabel metal1 25576 16014 25576 16014 0 mux_right_ipin_0.INVTX1_5_.out
rlabel metal1 27094 14314 27094 14314 0 mux_right_ipin_0.INVTX1_6_.out
rlabel metal2 19412 14926 19412 14926 0 mux_right_ipin_0.INVTX1_7_.out
rlabel metal2 21482 8092 21482 8092 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18952 6222 18952 6222 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20010 13639 20010 13639 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 8418 3060 8418 3060 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27232 25126 27232 25126 0 mux_right_ipin_1.INVTX1_2_.out
rlabel metal2 18722 17986 18722 17986 0 mux_right_ipin_1.INVTX1_3_.out
rlabel via1 22218 15997 22218 15997 0 mux_right_ipin_1.INVTX1_4_.out
rlabel metal1 20332 22406 20332 22406 0 mux_right_ipin_1.INVTX1_5_.out
rlabel metal1 22172 29002 22172 29002 0 mux_right_ipin_1.INVTX1_6_.out
rlabel metal2 10534 15844 10534 15844 0 mux_right_ipin_1.INVTX1_7_.out
rlabel metal1 24012 14858 24012 14858 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19688 15946 19688 15946 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19780 18190 19780 18190 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 18676 10166 18676 10166 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 27830 11492 27830 11492 0 mux_right_ipin_2.INVTX1_2_.out
rlabel metal2 27830 14110 27830 14110 0 mux_right_ipin_2.INVTX1_3_.out
rlabel metal1 23184 29002 23184 29002 0 mux_right_ipin_2.INVTX1_6_.out
rlabel metal2 15686 8160 15686 8160 0 mux_right_ipin_2.INVTX1_7_.out
rlabel metal1 17572 17102 17572 17102 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16330 13260 16330 13260 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15180 13294 15180 13294 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 10718 13396 10718 13396 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 25300 13974 25300 13974 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 21206 13515 21206 13515 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 24794 12716 24794 12716 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 29210 16320 29210 16320 0 mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 21344 13430 21344 13430 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18446 11594 18446 11594 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 15226 9180 15226 9180 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 18446 2482 18446 2482 0 mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 25070 18768 25070 18768 0 mux_right_ipin_5.INVTX1_4_.out
rlabel metal1 16744 14926 16744 14926 0 mux_right_ipin_5.INVTX1_5_.out
rlabel metal2 17158 3230 17158 3230 0 mux_right_ipin_5.INVTX1_6_.out
rlabel metal2 32062 20621 32062 20621 0 mux_right_ipin_5.INVTX1_7_.out
rlabel metal2 18722 7140 18722 7140 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 21068 14756 21068 14756 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17618 13044 17618 13044 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 17710 4488 17710 4488 0 mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 25760 14926 25760 14926 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19826 14892 19826 14892 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 24978 18190 24978 18190 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 30360 32402 30360 32402 0 mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 24012 19278 24012 19278 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 22816 16694 22816 16694 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20930 17952 20930 17952 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 12466 29546 12466 29546 0 mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 1794 3417 1794 3417 0 net1
rlabel metal2 22310 37026 22310 37026 0 net10
rlabel metal2 20286 19244 20286 19244 0 net100
rlabel metal1 18170 5746 18170 5746 0 net101
rlabel metal1 8418 20774 8418 20774 0 net11
rlabel metal1 12006 5678 12006 5678 0 net12
rlabel metal2 38042 14994 38042 14994 0 net13
rlabel metal2 37766 35326 37766 35326 0 net14
rlabel metal1 29026 25466 29026 25466 0 net15
rlabel metal2 28566 2278 28566 2278 0 net16
rlabel metal1 20700 29546 20700 29546 0 net17
rlabel metal1 11224 2550 11224 2550 0 net18
rlabel metal1 22678 28390 22678 28390 0 net19
rlabel metal1 7153 18326 7153 18326 0 net2
rlabel metal2 1886 25432 1886 25432 0 net20
rlabel metal2 38134 15708 38134 15708 0 net21
rlabel metal1 1978 36618 1978 36618 0 net22
rlabel metal2 1794 10336 1794 10336 0 net23
rlabel metal1 21160 25466 21160 25466 0 net24
rlabel metal1 2024 25874 2024 25874 0 net25
rlabel metal1 37950 37230 37950 37230 0 net26
rlabel metal1 5198 18734 5198 18734 0 net27
rlabel metal1 4462 2482 4462 2482 0 net28
rlabel metal1 5911 3026 5911 3026 0 net29
rlabel metal2 35742 2176 35742 2176 0 net3
rlabel metal1 32890 4794 32890 4794 0 net30
rlabel metal1 35604 13838 35604 13838 0 net31
rlabel metal1 25806 24684 25806 24684 0 net32
rlabel viali 27002 16559 27002 16559 0 net33
rlabel metal1 10074 36618 10074 36618 0 net34
rlabel metal1 37490 3570 37490 3570 0 net35
rlabel metal2 4094 11424 4094 11424 0 net36
rlabel metal2 33442 10948 33442 10948 0 net37
rlabel metal2 1978 19584 1978 19584 0 net38
rlabel metal1 30176 14994 30176 14994 0 net39
rlabel metal2 15226 36992 15226 36992 0 net4
rlabel metal2 9982 20604 9982 20604 0 net40
rlabel metal1 37168 36754 37168 36754 0 net41
rlabel metal1 4393 14382 4393 14382 0 net42
rlabel metal1 20148 27098 20148 27098 0 net43
rlabel metal1 37444 7718 37444 7718 0 net44
rlabel metal1 24334 37230 24334 37230 0 net45
rlabel metal1 1840 37230 1840 37230 0 net46
rlabel metal2 38042 30022 38042 30022 0 net47
rlabel metal2 4738 19380 4738 19380 0 net48
rlabel metal1 2392 23698 2392 23698 0 net49
rlabel metal1 16974 37298 16974 37298 0 net5
rlabel metal1 3312 3026 3312 3026 0 net50
rlabel metal1 34638 2414 34638 2414 0 net51
rlabel metal1 2116 33830 2116 33830 0 net52
rlabel metal1 26588 24650 26588 24650 0 net53
rlabel metal1 28244 37230 28244 37230 0 net54
rlabel metal1 20838 15980 20838 15980 0 net55
rlabel metal1 20838 37264 20838 37264 0 net56
rlabel metal1 37766 33490 37766 33490 0 net57
rlabel metal2 33534 7854 33534 7854 0 net58
rlabel metal2 1794 21318 1794 21318 0 net59
rlabel metal1 16376 37366 16376 37366 0 net6
rlabel metal1 36662 2380 36662 2380 0 net60
rlabel metal2 38042 22780 38042 22780 0 net61
rlabel metal1 16652 24106 16652 24106 0 net62
rlabel metal1 8924 36550 8924 36550 0 net63
rlabel metal1 18584 2414 18584 2414 0 net64
rlabel metal1 2622 2482 2622 2482 0 net65
rlabel metal2 19642 3910 19642 3910 0 net66
rlabel metal1 13340 36550 13340 36550 0 net67
rlabel metal2 22586 37060 22586 37060 0 net68
rlabel metal1 30774 36890 30774 36890 0 net69
rlabel metal1 14444 2278 14444 2278 0 net7
rlabel metal1 4370 26962 4370 26962 0 net70
rlabel metal1 5566 2448 5566 2448 0 net71
rlabel metal1 2162 2414 2162 2414 0 net72
rlabel metal2 38042 35700 38042 35700 0 net73
rlabel metal1 30452 37230 30452 37230 0 net74
rlabel metal1 16606 2414 16606 2414 0 net75
rlabel metal1 37030 36142 37030 36142 0 net76
rlabel metal1 37490 3026 37490 3026 0 net77
rlabel metal2 5474 36992 5474 36992 0 net78
rlabel metal2 37490 20604 37490 20604 0 net79
rlabel metal1 37306 8466 37306 8466 0 net8
rlabel metal2 7590 2618 7590 2618 0 net80
rlabel metal1 12006 2448 12006 2448 0 net81
rlabel metal2 10626 14790 10626 14790 0 net82
rlabel metal2 34086 21046 34086 21046 0 net83
rlabel metal1 18722 2618 18722 2618 0 net84
rlabel metal2 10350 4998 10350 4998 0 net85
rlabel metal2 32614 34884 32614 34884 0 net86
rlabel metal1 3542 37230 3542 37230 0 net87
rlabel metal2 10994 11526 10994 11526 0 net88
rlabel metal1 2162 34714 2162 34714 0 net89
rlabel metal2 23138 36448 23138 36448 0 net9
rlabel metal1 37812 18394 37812 18394 0 net90
rlabel metal1 15824 12274 15824 12274 0 net91
rlabel metal1 18262 10540 18262 10540 0 net92
rlabel metal1 24702 13838 24702 13838 0 net93
rlabel metal1 19458 18190 19458 18190 0 net94
rlabel metal2 14398 13804 14398 13804 0 net95
rlabel metal1 24288 10098 24288 10098 0 net96
rlabel metal1 14352 10574 14352 10574 0 net97
rlabel metal1 23368 12274 23368 12274 0 net98
rlabel metal2 25714 18462 25714 18462 0 net99
rlabel metal1 9798 37230 9798 37230 0 pReset
rlabel metal1 27140 2414 27140 2414 0 prog_clk
rlabel metal3 1188 12308 1188 12308 0 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
rlabel metal3 1188 36108 1188 36108 0 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
rlabel via2 38226 19125 38226 19125 0 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
