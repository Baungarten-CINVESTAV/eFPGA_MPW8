magic
tech sky130A
magscale 1 2
timestamp 1672416551
<< viali >>
rect 16221 37417 16255 37451
rect 26525 37417 26559 37451
rect 2421 37281 2455 37315
rect 9321 37281 9355 37315
rect 13277 37281 13311 37315
rect 17141 37281 17175 37315
rect 19441 37281 19475 37315
rect 27169 37281 27203 37315
rect 2145 37213 2179 37247
rect 3433 37213 3467 37247
rect 4169 37213 4203 37247
rect 4721 37213 4755 37247
rect 6009 37213 6043 37247
rect 6653 37213 6687 37247
rect 7849 37213 7883 37247
rect 9873 37213 9907 37247
rect 11989 37213 12023 37247
rect 12541 37213 12575 37247
rect 13093 37213 13127 37247
rect 15209 37213 15243 37247
rect 16957 37213 16991 37247
rect 18429 37213 18463 37247
rect 19717 37213 19751 37247
rect 22017 37213 22051 37247
rect 22753 37213 22787 37247
rect 24593 37213 24627 37247
rect 27445 37213 27479 37247
rect 28457 37213 28491 37247
rect 30021 37213 30055 37247
rect 31033 37213 31067 37247
rect 32965 37213 32999 37247
rect 35173 37213 35207 37247
rect 36093 37213 36127 37247
rect 3249 37077 3283 37111
rect 4813 37077 4847 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 9965 37077 9999 37111
rect 11805 37077 11839 37111
rect 15025 37077 15059 37111
rect 15669 37077 15703 37111
rect 18245 37077 18279 37111
rect 22201 37077 22235 37111
rect 22937 37077 22971 37111
rect 24777 37077 24811 37111
rect 28641 37077 28675 37111
rect 29837 37077 29871 37111
rect 31217 37077 31251 37111
rect 33149 37077 33183 37111
rect 34989 37077 35023 37111
rect 36277 37077 36311 37111
rect 2513 36873 2547 36907
rect 7665 36873 7699 36907
rect 12081 36873 12115 36907
rect 19349 36873 19383 36907
rect 27353 36873 27387 36907
rect 29837 36873 29871 36907
rect 35541 36873 35575 36907
rect 36277 36873 36311 36907
rect 1685 36805 1719 36839
rect 2329 36737 2363 36771
rect 7849 36737 7883 36771
rect 12265 36737 12299 36771
rect 12725 36737 12759 36771
rect 27169 36737 27203 36771
rect 29745 36737 29779 36771
rect 30389 36737 30423 36771
rect 34897 36737 34931 36771
rect 35357 36737 35391 36771
rect 36093 36737 36127 36771
rect 1869 36601 1903 36635
rect 3525 36533 3559 36567
rect 8309 36533 8343 36567
rect 18521 36533 18555 36567
rect 2329 36329 2363 36363
rect 35081 36125 35115 36159
rect 35541 36125 35575 36159
rect 35817 36125 35851 36159
rect 1685 36057 1719 36091
rect 1869 36057 1903 36091
rect 1685 35785 1719 35819
rect 2237 35785 2271 35819
rect 27353 35785 27387 35819
rect 36093 35785 36127 35819
rect 27169 35649 27203 35683
rect 27813 35649 27847 35683
rect 35909 35649 35943 35683
rect 21005 35241 21039 35275
rect 1869 35037 1903 35071
rect 20821 35037 20855 35071
rect 36093 35037 36127 35071
rect 36369 35037 36403 35071
rect 1685 34901 1719 34935
rect 21557 34901 21591 34935
rect 36369 34697 36403 34731
rect 36093 32861 36127 32895
rect 36369 32861 36403 32895
rect 1685 32793 1719 32827
rect 1869 32793 1903 32827
rect 1685 32521 1719 32555
rect 22201 32521 22235 32555
rect 36369 32521 36403 32555
rect 22017 32385 22051 32419
rect 22661 32385 22695 32419
rect 36093 31909 36127 31943
rect 1869 31773 1903 31807
rect 35633 31773 35667 31807
rect 36277 31773 36311 31807
rect 1685 31705 1719 31739
rect 29469 31433 29503 31467
rect 1593 31365 1627 31399
rect 29285 31297 29319 31331
rect 29929 31093 29963 31127
rect 29929 30277 29963 30311
rect 30021 30209 30055 30243
rect 30481 30209 30515 30243
rect 23949 29801 23983 29835
rect 34989 29801 35023 29835
rect 23765 29597 23799 29631
rect 34897 29597 34931 29631
rect 35541 29597 35575 29631
rect 1685 29529 1719 29563
rect 1869 29529 1903 29563
rect 36093 29529 36127 29563
rect 36277 29529 36311 29563
rect 24593 29461 24627 29495
rect 1593 29257 1627 29291
rect 36369 29257 36403 29291
rect 1869 28033 1903 28067
rect 13185 28033 13219 28067
rect 13829 28033 13863 28067
rect 20269 28033 20303 28067
rect 35633 28033 35667 28067
rect 36277 28033 36311 28067
rect 1685 27897 1719 27931
rect 13277 27897 13311 27931
rect 36093 27897 36127 27931
rect 2329 27829 2363 27863
rect 20361 27829 20395 27863
rect 7573 27557 7607 27591
rect 11989 27489 12023 27523
rect 7665 27421 7699 27455
rect 12081 27421 12115 27455
rect 29929 27421 29963 27455
rect 8125 27285 8159 27319
rect 29837 27285 29871 27319
rect 25697 26537 25731 26571
rect 36277 26469 36311 26503
rect 1869 26333 1903 26367
rect 25145 26333 25179 26367
rect 36093 26333 36127 26367
rect 2421 26265 2455 26299
rect 25053 26265 25087 26299
rect 1685 26197 1719 26231
rect 25973 24769 26007 24803
rect 25881 24565 25915 24599
rect 26617 24565 26651 24599
rect 35725 24157 35759 24191
rect 36369 24157 36403 24191
rect 1685 24089 1719 24123
rect 1869 24089 1903 24123
rect 36185 24021 36219 24055
rect 1593 23817 1627 23851
rect 24409 23817 24443 23851
rect 23765 23681 23799 23715
rect 23857 23477 23891 23511
rect 19533 23205 19567 23239
rect 21465 23137 21499 23171
rect 20177 23069 20211 23103
rect 20821 23001 20855 23035
rect 21373 23001 21407 23035
rect 20085 22933 20119 22967
rect 21005 22729 21039 22763
rect 1869 22593 1903 22627
rect 19809 22593 19843 22627
rect 20361 22593 20395 22627
rect 21097 22593 21131 22627
rect 27353 22593 27387 22627
rect 27813 22593 27847 22627
rect 36093 22593 36127 22627
rect 1685 22457 1719 22491
rect 36277 22457 36311 22491
rect 19717 22389 19751 22423
rect 22109 22389 22143 22423
rect 27261 22389 27295 22423
rect 22385 22049 22419 22083
rect 22477 21913 22511 21947
rect 23029 21913 23063 21947
rect 15393 21845 15427 21879
rect 20453 21845 20487 21879
rect 22845 21641 22879 21675
rect 15301 21573 15335 21607
rect 15393 21573 15427 21607
rect 15945 21573 15979 21607
rect 19993 21573 20027 21607
rect 20729 21573 20763 21607
rect 22937 21505 22971 21539
rect 23581 21505 23615 21539
rect 19441 21437 19475 21471
rect 20085 21437 20119 21471
rect 22293 21369 22327 21403
rect 24041 21369 24075 21403
rect 1593 21301 1627 21335
rect 20821 21301 20855 21335
rect 23489 21301 23523 21335
rect 25145 21301 25179 21335
rect 1593 20893 1627 20927
rect 1869 20893 1903 20927
rect 17601 20893 17635 20927
rect 18061 20893 18095 20927
rect 22477 20893 22511 20927
rect 23121 20893 23155 20927
rect 24961 20893 24995 20927
rect 25421 20893 25455 20927
rect 36093 20893 36127 20927
rect 20913 20825 20947 20859
rect 21005 20825 21039 20859
rect 21557 20825 21591 20859
rect 17509 20757 17543 20791
rect 22569 20757 22603 20791
rect 24869 20757 24903 20791
rect 25973 20757 26007 20791
rect 36277 20757 36311 20791
rect 1961 20553 1995 20587
rect 14933 20553 14967 20587
rect 21097 20553 21131 20587
rect 30021 20553 30055 20587
rect 18797 20485 18831 20519
rect 20085 20485 20119 20519
rect 20637 20485 20671 20519
rect 22753 20485 22787 20519
rect 22845 20485 22879 20519
rect 24685 20485 24719 20519
rect 26525 20485 26559 20519
rect 1777 20417 1811 20451
rect 14841 20417 14875 20451
rect 25237 20417 25271 20451
rect 25881 20417 25915 20451
rect 29929 20417 29963 20451
rect 18705 20349 18739 20383
rect 19993 20349 20027 20383
rect 23397 20349 23431 20383
rect 19257 20281 19291 20315
rect 22293 20281 22327 20315
rect 25329 20281 25363 20315
rect 2513 20213 2547 20247
rect 24593 20213 24627 20247
rect 25973 20213 26007 20247
rect 19625 20009 19659 20043
rect 23949 19941 23983 19975
rect 22201 19873 22235 19907
rect 25237 19873 25271 19907
rect 25881 19873 25915 19907
rect 16129 19805 16163 19839
rect 16589 19805 16623 19839
rect 19533 19805 19567 19839
rect 20177 19805 20211 19839
rect 20913 19805 20947 19839
rect 21373 19805 21407 19839
rect 22109 19805 22143 19839
rect 17233 19737 17267 19771
rect 18613 19737 18647 19771
rect 22753 19737 22787 19771
rect 23305 19737 23339 19771
rect 23397 19737 23431 19771
rect 24593 19737 24627 19771
rect 25145 19737 25179 19771
rect 25973 19737 26007 19771
rect 26525 19737 26559 19771
rect 27077 19737 27111 19771
rect 27169 19737 27203 19771
rect 27721 19737 27755 19771
rect 16037 19669 16071 19703
rect 17693 19669 17727 19703
rect 21465 19669 21499 19703
rect 15117 19465 15151 19499
rect 19349 19465 19383 19499
rect 22109 19465 22143 19499
rect 25789 19465 25823 19499
rect 27169 19465 27203 19499
rect 32505 19465 32539 19499
rect 17325 19397 17359 19431
rect 23397 19397 23431 19431
rect 24961 19397 24995 19431
rect 25053 19397 25087 19431
rect 1685 19329 1719 19363
rect 15669 19329 15703 19363
rect 16129 19329 16163 19363
rect 16221 19329 16255 19363
rect 19257 19329 19291 19363
rect 22017 19329 22051 19363
rect 25605 19329 25639 19363
rect 26433 19329 26467 19363
rect 32321 19329 32355 19363
rect 32965 19329 32999 19363
rect 36093 19329 36127 19363
rect 17233 19261 17267 19295
rect 17877 19261 17911 19295
rect 21373 19261 21407 19295
rect 22661 19261 22695 19295
rect 23305 19261 23339 19295
rect 23581 19261 23615 19295
rect 24409 19261 24443 19295
rect 27813 19261 27847 19295
rect 1869 19193 1903 19227
rect 14565 19125 14599 19159
rect 18705 19125 18739 19159
rect 19993 19125 20027 19159
rect 20913 19125 20947 19159
rect 26341 19125 26375 19159
rect 36277 19125 36311 19159
rect 1593 18921 1627 18955
rect 13737 18921 13771 18955
rect 16129 18921 16163 18955
rect 27813 18921 27847 18955
rect 23213 18853 23247 18887
rect 18797 18785 18831 18819
rect 25697 18785 25731 18819
rect 25973 18785 26007 18819
rect 14657 18717 14691 18751
rect 15301 18717 15335 18751
rect 16037 18717 16071 18751
rect 16681 18717 16715 18751
rect 20361 18717 20395 18751
rect 21097 18717 21131 18751
rect 21833 18717 21867 18751
rect 22385 18717 22419 18751
rect 24593 18717 24627 18751
rect 26709 18717 26743 18751
rect 27169 18717 27203 18751
rect 28365 18717 28399 18751
rect 17785 18649 17819 18683
rect 18705 18649 18739 18683
rect 23673 18649 23707 18683
rect 23765 18649 23799 18683
rect 25881 18649 25915 18683
rect 14749 18581 14783 18615
rect 15393 18581 15427 18615
rect 16773 18581 16807 18615
rect 19533 18581 19567 18615
rect 20269 18581 20303 18615
rect 21741 18581 21775 18615
rect 22477 18581 22511 18615
rect 24685 18581 24719 18615
rect 26617 18581 26651 18615
rect 27261 18581 27295 18615
rect 24041 18377 24075 18411
rect 27813 18377 27847 18411
rect 14105 18309 14139 18343
rect 14197 18309 14231 18343
rect 15393 18309 15427 18343
rect 15945 18309 15979 18343
rect 17785 18309 17819 18343
rect 18337 18309 18371 18343
rect 20269 18309 20303 18343
rect 20821 18309 20855 18343
rect 22569 18309 22603 18343
rect 22661 18309 22695 18343
rect 23581 18309 23615 18343
rect 25605 18309 25639 18343
rect 12725 18241 12759 18275
rect 13185 18241 13219 18275
rect 16957 18241 16991 18275
rect 18981 18241 19015 18275
rect 21281 18241 21315 18275
rect 27353 18241 27387 18275
rect 28365 18241 28399 18275
rect 14749 18173 14783 18207
rect 15301 18173 15335 18207
rect 17693 18173 17727 18207
rect 20177 18173 20211 18207
rect 24685 18173 24719 18207
rect 25513 18173 25547 18207
rect 26157 18173 26191 18207
rect 17049 18105 17083 18139
rect 13277 18037 13311 18071
rect 18889 18037 18923 18071
rect 19625 18037 19659 18071
rect 21373 18037 21407 18071
rect 27261 18037 27295 18071
rect 29009 18037 29043 18071
rect 10701 17833 10735 17867
rect 12449 17833 12483 17867
rect 13645 17833 13679 17867
rect 15025 17765 15059 17799
rect 26157 17765 26191 17799
rect 28641 17765 28675 17799
rect 16221 17697 16255 17731
rect 17417 17697 17451 17731
rect 19533 17697 19567 17731
rect 21373 17697 21407 17731
rect 22017 17697 22051 17731
rect 22937 17697 22971 17731
rect 23949 17697 23983 17731
rect 27445 17697 27479 17731
rect 28457 17697 28491 17731
rect 11253 17629 11287 17663
rect 13093 17629 13127 17663
rect 13553 17629 13587 17663
rect 14289 17629 14323 17663
rect 18705 17629 18739 17663
rect 20821 17629 20855 17663
rect 28273 17629 28307 17663
rect 11345 17561 11379 17595
rect 15485 17561 15519 17595
rect 15577 17561 15611 17595
rect 16313 17561 16347 17595
rect 16865 17561 16899 17595
rect 17509 17561 17543 17595
rect 18061 17561 18095 17595
rect 19625 17561 19659 17595
rect 20177 17561 20211 17595
rect 21465 17561 21499 17595
rect 23029 17561 23063 17595
rect 24685 17561 24719 17595
rect 24777 17561 24811 17595
rect 25697 17561 25731 17595
rect 27629 17561 27663 17595
rect 27721 17561 27755 17595
rect 13001 17493 13035 17527
rect 14381 17493 14415 17527
rect 18797 17493 18831 17527
rect 20729 17493 20763 17527
rect 29745 17493 29779 17527
rect 9965 17289 9999 17323
rect 16221 17289 16255 17323
rect 16957 17289 16991 17323
rect 26065 17289 26099 17323
rect 15117 17221 15151 17255
rect 17509 17221 17543 17255
rect 18061 17221 18095 17255
rect 19257 17221 19291 17255
rect 19349 17221 19383 17255
rect 20913 17221 20947 17255
rect 21005 17221 21039 17255
rect 22201 17221 22235 17255
rect 23305 17221 23339 17255
rect 23397 17221 23431 17255
rect 24961 17221 24995 17255
rect 1685 17153 1719 17187
rect 9505 17153 9539 17187
rect 12173 17153 12207 17187
rect 13277 17153 13311 17187
rect 13461 17153 13495 17187
rect 14289 17153 14323 17187
rect 16129 17153 16163 17187
rect 16865 17153 16899 17187
rect 20361 17153 20395 17187
rect 26157 17153 26191 17187
rect 27353 17153 27387 17187
rect 27997 17153 28031 17187
rect 29101 17153 29135 17187
rect 36093 17153 36127 17187
rect 15025 17085 15059 17119
rect 15301 17085 15335 17119
rect 18153 17085 18187 17119
rect 22109 17085 22143 17119
rect 24317 17085 24351 17119
rect 24869 17085 24903 17119
rect 28641 17085 28675 17119
rect 1869 17017 1903 17051
rect 12265 17017 12299 17051
rect 18797 17017 18831 17051
rect 22661 17017 22695 17051
rect 25421 17017 25455 17051
rect 27905 17017 27939 17051
rect 29285 17017 29319 17051
rect 36277 17017 36311 17051
rect 9321 16949 9355 16983
rect 11161 16949 11195 16983
rect 13093 16949 13127 16983
rect 14381 16949 14415 16983
rect 27261 16949 27295 16983
rect 29745 16949 29779 16983
rect 30297 16949 30331 16983
rect 1685 16745 1719 16779
rect 13461 16745 13495 16779
rect 17785 16745 17819 16779
rect 21189 16745 21223 16779
rect 29837 16745 29871 16779
rect 15025 16677 15059 16711
rect 16221 16677 16255 16711
rect 11253 16609 11287 16643
rect 13277 16609 13311 16643
rect 16773 16609 16807 16643
rect 20269 16609 20303 16643
rect 20545 16609 20579 16643
rect 22845 16609 22879 16643
rect 24961 16609 24995 16643
rect 25789 16609 25823 16643
rect 26433 16609 26467 16643
rect 27629 16609 27663 16643
rect 28273 16609 28307 16643
rect 30297 16609 30331 16643
rect 11805 16541 11839 16575
rect 12633 16541 12667 16575
rect 13093 16541 13127 16575
rect 14289 16541 14323 16575
rect 17693 16541 17727 16575
rect 18705 16541 18739 16575
rect 21281 16541 21315 16575
rect 23581 16541 23615 16575
rect 29009 16541 29043 16575
rect 11897 16473 11931 16507
rect 15485 16473 15519 16507
rect 15577 16473 15611 16507
rect 16681 16473 16715 16507
rect 20453 16473 20487 16507
rect 22201 16473 22235 16507
rect 22753 16473 22787 16507
rect 23489 16473 23523 16507
rect 25053 16473 25087 16507
rect 26985 16473 27019 16507
rect 27077 16473 27111 16507
rect 28181 16473 28215 16507
rect 12541 16405 12575 16439
rect 14473 16405 14507 16439
rect 18797 16405 18831 16439
rect 28917 16405 28951 16439
rect 31033 16405 31067 16439
rect 2329 16201 2363 16235
rect 11069 16201 11103 16235
rect 27905 16201 27939 16235
rect 29101 16201 29135 16235
rect 30297 16201 30331 16235
rect 31309 16201 31343 16235
rect 15301 16133 15335 16167
rect 17049 16133 17083 16167
rect 19441 16133 19475 16167
rect 22477 16133 22511 16167
rect 23029 16133 23063 16167
rect 24225 16133 24259 16167
rect 25513 16133 25547 16167
rect 1869 16065 1903 16099
rect 2513 16065 2547 16099
rect 12541 16065 12575 16099
rect 12633 16065 12667 16099
rect 13277 16065 13311 16099
rect 14197 16065 14231 16099
rect 14381 16065 14415 16099
rect 18705 16065 18739 16099
rect 20545 16065 20579 16099
rect 21373 16065 21407 16099
rect 27353 16065 27387 16099
rect 28365 16065 28399 16099
rect 28549 16065 28583 16099
rect 29193 16065 29227 16099
rect 29653 16065 29687 16099
rect 31125 16065 31159 16099
rect 36093 16065 36127 16099
rect 11897 15997 11931 16031
rect 13737 15997 13771 16031
rect 15209 15997 15243 16031
rect 16957 15997 16991 16031
rect 17601 15997 17635 16031
rect 19349 15997 19383 16031
rect 23121 15997 23155 16031
rect 23673 15997 23707 16031
rect 24317 15997 24351 16031
rect 25421 15997 25455 16031
rect 25789 15997 25823 16031
rect 10517 15929 10551 15963
rect 13185 15929 13219 15963
rect 15761 15929 15795 15963
rect 18521 15929 18555 15963
rect 19901 15929 19935 15963
rect 20637 15929 20671 15963
rect 29745 15929 29779 15963
rect 1685 15861 1719 15895
rect 2973 15861 3007 15895
rect 21281 15861 21315 15895
rect 27261 15861 27295 15895
rect 36277 15861 36311 15895
rect 3985 15657 4019 15691
rect 4721 15657 4755 15691
rect 23581 15657 23615 15691
rect 31125 15657 31159 15691
rect 11161 15589 11195 15623
rect 27077 15589 27111 15623
rect 10609 15521 10643 15555
rect 13645 15521 13679 15555
rect 18613 15521 18647 15555
rect 21189 15521 21223 15555
rect 22385 15521 22419 15555
rect 24593 15521 24627 15555
rect 25237 15521 25271 15555
rect 26433 15521 26467 15555
rect 28457 15521 28491 15555
rect 29101 15521 29135 15555
rect 4169 15453 4203 15487
rect 11621 15453 11655 15487
rect 12265 15453 12299 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 14289 15453 14323 15487
rect 15669 15453 15703 15487
rect 19533 15453 19567 15487
rect 20361 15453 20395 15487
rect 23673 15453 23707 15487
rect 29929 15453 29963 15487
rect 30389 15453 30423 15487
rect 31033 15453 31067 15487
rect 13001 15385 13035 15419
rect 15025 15385 15059 15419
rect 15117 15385 15151 15419
rect 16681 15385 16715 15419
rect 17233 15385 17267 15419
rect 17325 15385 17359 15419
rect 17969 15385 18003 15419
rect 18061 15385 18095 15419
rect 20269 15385 20303 15419
rect 21281 15385 21315 15419
rect 21833 15385 21867 15419
rect 22477 15385 22511 15419
rect 23029 15385 23063 15419
rect 25145 15385 25179 15419
rect 25789 15385 25823 15419
rect 26341 15385 26375 15419
rect 27537 15385 27571 15419
rect 27629 15385 27663 15419
rect 28549 15385 28583 15419
rect 11713 15317 11747 15351
rect 12357 15317 12391 15351
rect 14381 15317 14415 15351
rect 16129 15317 16163 15351
rect 19625 15317 19659 15351
rect 29837 15317 29871 15351
rect 30481 15317 30515 15351
rect 17233 15113 17267 15147
rect 20913 15113 20947 15147
rect 28641 15113 28675 15147
rect 36001 15113 36035 15147
rect 9965 15045 9999 15079
rect 11161 15045 11195 15079
rect 13553 15045 13587 15079
rect 14381 15045 14415 15079
rect 16221 15045 16255 15079
rect 17969 15045 18003 15079
rect 20177 15045 20211 15079
rect 20269 15045 20303 15079
rect 22569 15045 22603 15079
rect 23397 15045 23431 15079
rect 24501 15045 24535 15079
rect 24593 15045 24627 15079
rect 25789 15045 25823 15079
rect 27629 15045 27663 15079
rect 28181 15045 28215 15079
rect 30665 15045 30699 15079
rect 10609 14977 10643 15011
rect 11989 14977 12023 15011
rect 16129 14977 16163 15011
rect 17141 14977 17175 15011
rect 19165 14977 19199 15011
rect 21005 14977 21039 15011
rect 29101 14977 29135 15011
rect 31217 14977 31251 15011
rect 36093 14977 36127 15011
rect 13369 14909 13403 14943
rect 13645 14909 13679 14943
rect 14289 14909 14323 14943
rect 15117 14909 15151 14943
rect 17877 14909 17911 14943
rect 22661 14909 22695 14943
rect 23305 14909 23339 14943
rect 23949 14909 23983 14943
rect 24777 14909 24811 14943
rect 25697 14909 25731 14943
rect 26341 14909 26375 14943
rect 27537 14909 27571 14943
rect 29285 14909 29319 14943
rect 18429 14841 18463 14875
rect 19717 14841 19751 14875
rect 22109 14841 22143 14875
rect 12081 14773 12115 14807
rect 19073 14773 19107 14807
rect 29745 14773 29779 14807
rect 30389 14773 30423 14807
rect 21281 14569 21315 14603
rect 23949 14569 23983 14603
rect 29837 14569 29871 14603
rect 10609 14501 10643 14535
rect 13645 14501 13679 14535
rect 16037 14501 16071 14535
rect 17233 14501 17267 14535
rect 26249 14501 26283 14535
rect 10057 14433 10091 14467
rect 11805 14433 11839 14467
rect 18245 14433 18279 14467
rect 18889 14433 18923 14467
rect 23397 14433 23431 14467
rect 26801 14433 26835 14467
rect 11253 14365 11287 14399
rect 11713 14365 11747 14399
rect 12357 14365 12391 14399
rect 14749 14365 14783 14399
rect 21373 14365 21407 14399
rect 23857 14365 23891 14399
rect 28089 14365 28123 14399
rect 28549 14365 28583 14399
rect 29929 14365 29963 14399
rect 30389 14365 30423 14399
rect 31125 14365 31159 14399
rect 13093 14297 13127 14331
rect 13185 14297 13219 14331
rect 15485 14297 15519 14331
rect 15577 14297 15611 14331
rect 16681 14297 16715 14331
rect 16773 14297 16807 14331
rect 18337 14297 18371 14331
rect 19993 14297 20027 14331
rect 20545 14297 20579 14331
rect 20637 14297 20671 14331
rect 22385 14297 22419 14331
rect 22477 14297 22511 14331
rect 24593 14297 24627 14331
rect 25513 14297 25547 14331
rect 25605 14297 25639 14331
rect 26709 14297 26743 14331
rect 27445 14297 27479 14331
rect 27537 14297 27571 14331
rect 31585 14297 31619 14331
rect 9505 14229 9539 14263
rect 11161 14229 11195 14263
rect 12449 14229 12483 14263
rect 14841 14229 14875 14263
rect 19441 14229 19475 14263
rect 28641 14229 28675 14263
rect 30481 14229 30515 14263
rect 11069 14025 11103 14059
rect 13921 14025 13955 14059
rect 22109 14025 22143 14059
rect 22753 14025 22787 14059
rect 26249 14025 26283 14059
rect 36185 14025 36219 14059
rect 12633 13957 12667 13991
rect 13185 13957 13219 13991
rect 14565 13957 14599 13991
rect 15669 13957 15703 13991
rect 15761 13957 15795 13991
rect 17325 13957 17359 13991
rect 17417 13957 17451 13991
rect 18337 13957 18371 13991
rect 18981 13957 19015 13991
rect 19993 13957 20027 13991
rect 20545 13957 20579 13991
rect 21373 13957 21407 13991
rect 23581 13957 23615 13991
rect 25513 13957 25547 13991
rect 27261 13957 27295 13991
rect 27353 13957 27387 13991
rect 28549 13957 28583 13991
rect 29101 13957 29135 13991
rect 30297 13957 30331 13991
rect 1869 13889 1903 13923
rect 8585 13889 8619 13923
rect 9137 13889 9171 13923
rect 10149 13889 10183 13923
rect 11161 13889 11195 13923
rect 11805 13889 11839 13923
rect 21281 13889 21315 13923
rect 22201 13889 22235 13923
rect 22661 13889 22695 13923
rect 26341 13889 26375 13923
rect 29745 13889 29779 13923
rect 30205 13889 30239 13923
rect 30849 13889 30883 13923
rect 35725 13889 35759 13923
rect 36369 13889 36403 13923
rect 10241 13821 10275 13855
rect 11897 13821 11931 13855
rect 12541 13821 12575 13855
rect 14473 13821 14507 13855
rect 18889 13821 18923 13855
rect 19533 13821 19567 13855
rect 20637 13821 20671 13855
rect 23489 13821 23523 13855
rect 24409 13821 24443 13855
rect 25329 13821 25363 13855
rect 25605 13821 25639 13855
rect 27905 13821 27939 13855
rect 28457 13821 28491 13855
rect 31401 13821 31435 13855
rect 9689 13753 9723 13787
rect 15025 13753 15059 13787
rect 16221 13753 16255 13787
rect 1685 13685 1719 13719
rect 29653 13685 29687 13719
rect 18889 13481 18923 13515
rect 23857 13481 23891 13515
rect 25329 13481 25363 13515
rect 31585 13481 31619 13515
rect 8401 13413 8435 13447
rect 17509 13413 17543 13447
rect 29837 13413 29871 13447
rect 9873 13345 9907 13379
rect 11713 13345 11747 13379
rect 12173 13345 12207 13379
rect 13093 13345 13127 13379
rect 13369 13345 13403 13379
rect 14381 13345 14415 13379
rect 15761 13345 15795 13379
rect 16405 13345 16439 13379
rect 19533 13345 19567 13379
rect 19809 13345 19843 13379
rect 21097 13345 21131 13379
rect 21741 13345 21775 13379
rect 24685 13345 24719 13379
rect 27905 13345 27939 13379
rect 28181 13345 28215 13379
rect 29101 13345 29135 13379
rect 8309 13277 8343 13311
rect 9137 13277 9171 13311
rect 9781 13277 9815 13311
rect 23765 13277 23799 13311
rect 24777 13277 24811 13311
rect 25237 13277 25271 13311
rect 29009 13277 29043 13311
rect 31125 13277 31159 13311
rect 9229 13209 9263 13243
rect 10425 13209 10459 13243
rect 10977 13209 11011 13243
rect 11069 13209 11103 13243
rect 11805 13209 11839 13243
rect 13162 13209 13196 13243
rect 14473 13209 14507 13243
rect 15025 13209 15059 13243
rect 15853 13209 15887 13243
rect 16957 13209 16991 13243
rect 17049 13209 17083 13243
rect 18245 13209 18279 13243
rect 19625 13209 19659 13243
rect 21189 13209 21223 13243
rect 22293 13209 22327 13243
rect 22385 13209 22419 13243
rect 22937 13209 22971 13243
rect 26249 13209 26283 13243
rect 27169 13209 27203 13243
rect 27261 13209 27295 13243
rect 27997 13209 28031 13243
rect 30297 13209 30331 13243
rect 30389 13209 30423 13243
rect 31033 13209 31067 13243
rect 18153 13141 18187 13175
rect 2145 12937 2179 12971
rect 2881 12937 2915 12971
rect 8033 12937 8067 12971
rect 9781 12937 9815 12971
rect 12081 12937 12115 12971
rect 19257 12937 19291 12971
rect 21373 12937 21407 12971
rect 27261 12937 27295 12971
rect 28549 12937 28583 12971
rect 29837 12937 29871 12971
rect 31125 12937 31159 12971
rect 31769 12937 31803 12971
rect 12817 12869 12851 12903
rect 14933 12869 14967 12903
rect 15761 12869 15795 12903
rect 16313 12869 16347 12903
rect 17509 12869 17543 12903
rect 18429 12869 18463 12903
rect 20637 12869 20671 12903
rect 22385 12869 22419 12903
rect 25973 12869 26007 12903
rect 29101 12869 29135 12903
rect 2329 12801 2363 12835
rect 8677 12801 8711 12835
rect 9689 12801 9723 12835
rect 10517 12801 10551 12835
rect 10977 12801 11011 12835
rect 11989 12801 12023 12835
rect 19349 12801 19383 12835
rect 21281 12801 21315 12835
rect 22937 12801 22971 12835
rect 23581 12801 23615 12835
rect 24041 12801 24075 12835
rect 24777 12801 24811 12835
rect 24869 12801 24903 12835
rect 27353 12801 27387 12835
rect 27813 12801 27847 12835
rect 28641 12801 28675 12835
rect 29745 12801 29779 12835
rect 30573 12801 30607 12835
rect 31217 12801 31251 12835
rect 32321 12801 32355 12835
rect 9229 12733 9263 12767
rect 12725 12733 12759 12767
rect 13001 12733 13035 12767
rect 14381 12733 14415 12767
rect 15025 12733 15059 12767
rect 15669 12733 15703 12767
rect 17417 12733 17451 12767
rect 20453 12733 20487 12767
rect 20729 12733 20763 12767
rect 22293 12733 22327 12767
rect 25605 12733 25639 12767
rect 26065 12733 26099 12767
rect 27905 12733 27939 12767
rect 11069 12665 11103 12699
rect 23489 12665 23523 12699
rect 10425 12597 10459 12631
rect 13921 12597 13955 12631
rect 24133 12597 24167 12631
rect 30389 12597 30423 12631
rect 10701 12393 10735 12427
rect 20177 12393 20211 12427
rect 21833 12393 21867 12427
rect 30941 12393 30975 12427
rect 31585 12393 31619 12427
rect 16129 12325 16163 12359
rect 18797 12325 18831 12359
rect 21281 12325 21315 12359
rect 12081 12257 12115 12291
rect 13461 12257 13495 12291
rect 14657 12257 14691 12291
rect 17325 12257 17359 12291
rect 19533 12257 19567 12291
rect 23029 12257 23063 12291
rect 25237 12257 25271 12291
rect 28641 12257 28675 12291
rect 29837 12257 29871 12291
rect 1961 12189 1995 12223
rect 7297 12189 7331 12223
rect 7757 12189 7791 12223
rect 8401 12189 8435 12223
rect 9321 12189 9355 12223
rect 9965 12189 9999 12223
rect 10793 12189 10827 12223
rect 11253 12189 11287 12223
rect 11897 12189 11931 12223
rect 13645 12189 13679 12223
rect 15301 12189 15335 12223
rect 18705 12189 18739 12223
rect 19441 12189 19475 12223
rect 20085 12189 20119 12223
rect 21189 12189 21223 12223
rect 22385 12189 22419 12223
rect 23765 12189 23799 12223
rect 26525 12189 26559 12223
rect 26617 12189 26651 12223
rect 28733 12189 28767 12223
rect 8493 12121 8527 12155
rect 14749 12121 14783 12155
rect 16589 12121 16623 12155
rect 16681 12121 16715 12155
rect 17417 12121 17451 12155
rect 17969 12121 18003 12155
rect 22937 12121 22971 12155
rect 24593 12121 24627 12155
rect 25145 12121 25179 12155
rect 25789 12121 25823 12155
rect 25973 12121 26007 12155
rect 27445 12121 27479 12155
rect 27537 12121 27571 12155
rect 28089 12121 28123 12155
rect 29929 12121 29963 12155
rect 30481 12121 30515 12155
rect 1777 12053 1811 12087
rect 7849 12053 7883 12087
rect 9505 12053 9539 12087
rect 10057 12053 10091 12087
rect 11345 12053 11379 12087
rect 12541 12053 12575 12087
rect 13001 12053 13035 12087
rect 23673 12053 23707 12087
rect 32137 12053 32171 12087
rect 8677 11849 8711 11883
rect 9229 11849 9263 11883
rect 16221 11849 16255 11883
rect 17785 11849 17819 11883
rect 21189 11849 21223 11883
rect 22201 11849 22235 11883
rect 25881 11849 25915 11883
rect 26525 11849 26559 11883
rect 27261 11849 27295 11883
rect 27905 11849 27939 11883
rect 29837 11849 29871 11883
rect 11897 11781 11931 11815
rect 13277 11781 13311 11815
rect 14565 11781 14599 11815
rect 14657 11781 14691 11815
rect 18613 11781 18647 11815
rect 19901 11781 19935 11815
rect 20453 11781 20487 11815
rect 20545 11781 20579 11815
rect 23213 11781 23247 11815
rect 28549 11781 28583 11815
rect 30389 11781 30423 11815
rect 1869 11713 1903 11747
rect 9873 11713 9907 11747
rect 10517 11713 10551 11747
rect 10977 11713 11011 11747
rect 13829 11713 13863 11747
rect 16129 11713 16163 11747
rect 17233 11713 17267 11747
rect 17877 11713 17911 11747
rect 21281 11713 21315 11747
rect 25329 11713 25363 11747
rect 25789 11713 25823 11747
rect 26617 11713 26651 11747
rect 27353 11713 27387 11747
rect 27997 11713 28031 11747
rect 28641 11713 28675 11747
rect 29285 11713 29319 11747
rect 29745 11713 29779 11747
rect 35633 11713 35667 11747
rect 36277 11713 36311 11747
rect 11805 11645 11839 11679
rect 12081 11645 12115 11679
rect 13185 11645 13219 11679
rect 14841 11645 14875 11679
rect 18521 11645 18555 11679
rect 18797 11645 18831 11679
rect 22937 11645 22971 11679
rect 30941 11645 30975 11679
rect 1685 11577 1719 11611
rect 9781 11577 9815 11611
rect 36093 11577 36127 11611
rect 8125 11509 8159 11543
rect 10425 11509 10459 11543
rect 11069 11509 11103 11543
rect 17141 11509 17175 11543
rect 24685 11509 24719 11543
rect 25237 11509 25271 11543
rect 29193 11509 29227 11543
rect 31493 11509 31527 11543
rect 9505 11305 9539 11339
rect 14565 11305 14599 11339
rect 18153 11305 18187 11339
rect 25329 11305 25363 11339
rect 26617 11305 26651 11339
rect 27905 11305 27939 11339
rect 29837 11305 29871 11339
rect 11345 11237 11379 11271
rect 12265 11237 12299 11271
rect 18797 11237 18831 11271
rect 21465 11237 21499 11271
rect 25973 11237 26007 11271
rect 30389 11237 30423 11271
rect 10149 11169 10183 11203
rect 10793 11169 10827 11203
rect 12909 11169 12943 11203
rect 13277 11169 13311 11203
rect 16681 11169 16715 11203
rect 19717 11169 19751 11203
rect 30941 11169 30975 11203
rect 10057 11101 10091 11135
rect 12357 11101 12391 11135
rect 14473 11101 14507 11135
rect 16957 11101 16991 11135
rect 17509 11101 17543 11135
rect 17601 11101 17635 11135
rect 18061 11101 18095 11135
rect 18889 11101 18923 11135
rect 22109 11101 22143 11135
rect 22661 11101 22695 11135
rect 22753 11101 22787 11135
rect 23397 11101 23431 11135
rect 24041 11101 24075 11135
rect 24777 11101 24811 11135
rect 25421 11101 25455 11135
rect 26065 11101 26099 11135
rect 26709 11101 26743 11135
rect 27353 11101 27387 11135
rect 27813 11101 27847 11135
rect 28549 11101 28583 11135
rect 28641 11101 28675 11135
rect 29193 11101 29227 11135
rect 29745 11101 29779 11135
rect 32045 11101 32079 11135
rect 7941 11033 7975 11067
rect 8033 11033 8067 11067
rect 8585 11033 8619 11067
rect 10885 11033 10919 11067
rect 13001 11033 13035 11067
rect 19993 11033 20027 11067
rect 23305 11033 23339 11067
rect 23949 11033 23983 11067
rect 24685 11033 24719 11067
rect 31493 11033 31527 11067
rect 15209 10965 15243 10999
rect 22017 10965 22051 10999
rect 27261 10965 27295 10999
rect 8033 10761 8067 10795
rect 8769 10761 8803 10795
rect 13185 10761 13219 10795
rect 16957 10761 16991 10795
rect 25145 10761 25179 10795
rect 26433 10761 26467 10795
rect 27261 10761 27295 10795
rect 35541 10761 35575 10795
rect 10517 10693 10551 10727
rect 14749 10693 14783 10727
rect 17785 10693 17819 10727
rect 19993 10693 20027 10727
rect 23673 10693 23707 10727
rect 28089 10693 28123 10727
rect 28641 10693 28675 10727
rect 30297 10693 30331 10727
rect 1869 10625 1903 10659
rect 8861 10625 8895 10659
rect 11161 10625 11195 10659
rect 11805 10625 11839 10659
rect 13093 10625 13127 10659
rect 13829 10625 13863 10659
rect 16865 10625 16899 10659
rect 22201 10625 22235 10659
rect 22845 10625 22879 10659
rect 23397 10625 23431 10659
rect 25881 10625 25915 10659
rect 26341 10625 26375 10659
rect 27169 10625 27203 10659
rect 29745 10625 29779 10659
rect 30389 10625 30423 10659
rect 31033 10625 31067 10659
rect 36093 10625 36127 10659
rect 11069 10557 11103 10591
rect 11989 10557 12023 10591
rect 14013 10557 14047 10591
rect 14473 10557 14507 10591
rect 17509 10557 17543 10591
rect 19257 10557 19291 10591
rect 19717 10557 19751 10591
rect 22753 10557 22787 10591
rect 28733 10557 28767 10591
rect 29469 10557 29503 10591
rect 31493 10557 31527 10591
rect 9965 10489 9999 10523
rect 25789 10489 25823 10523
rect 1685 10421 1719 10455
rect 9413 10421 9447 10455
rect 12449 10421 12483 10455
rect 16221 10421 16255 10455
rect 21465 10421 21499 10455
rect 22109 10421 22143 10455
rect 30941 10421 30975 10455
rect 36277 10421 36311 10455
rect 10333 10217 10367 10251
rect 11713 10217 11747 10251
rect 12357 10217 12391 10251
rect 13645 10217 13679 10251
rect 18797 10217 18831 10251
rect 23121 10217 23155 10251
rect 27169 10217 27203 10251
rect 15117 10081 15151 10115
rect 17141 10081 17175 10115
rect 10885 10013 10919 10047
rect 11621 10013 11655 10047
rect 12265 10013 12299 10047
rect 12909 10013 12943 10047
rect 13737 10013 13771 10047
rect 14473 10013 14507 10047
rect 18061 10013 18095 10047
rect 18889 10013 18923 10047
rect 19901 10013 19935 10047
rect 20545 10013 20579 10047
rect 23213 10013 23247 10047
rect 23857 10013 23891 10047
rect 26617 10013 26651 10047
rect 27077 10013 27111 10047
rect 27905 10013 27939 10047
rect 29193 10013 29227 10047
rect 31125 10013 31159 10047
rect 31585 10013 31619 10047
rect 8493 9945 8527 9979
rect 9873 9945 9907 9979
rect 13001 9945 13035 9979
rect 15393 9945 15427 9979
rect 20821 9945 20855 9979
rect 22569 9945 22603 9979
rect 24593 9945 24627 9979
rect 26341 9945 26375 9979
rect 28917 9945 28951 9979
rect 29745 9945 29779 9979
rect 30297 9945 30331 9979
rect 30389 9945 30423 9979
rect 9321 9877 9355 9911
rect 10977 9877 11011 9911
rect 14565 9877 14599 9911
rect 18153 9877 18187 9911
rect 19993 9877 20027 9911
rect 23765 9877 23799 9911
rect 27813 9877 27847 9911
rect 31033 9877 31067 9911
rect 10609 9605 10643 9639
rect 12265 9605 12299 9639
rect 12357 9605 12391 9639
rect 13277 9605 13311 9639
rect 16957 9605 16991 9639
rect 19441 9605 19475 9639
rect 25421 9605 25455 9639
rect 30021 9605 30055 9639
rect 30573 9605 30607 9639
rect 30665 9605 30699 9639
rect 11161 9537 11195 9571
rect 13185 9537 13219 9571
rect 13829 9537 13863 9571
rect 20453 9537 20487 9571
rect 21097 9537 21131 9571
rect 24501 9537 24535 9571
rect 25513 9537 25547 9571
rect 26133 9535 26167 9569
rect 27353 9537 27387 9571
rect 27997 9537 28031 9571
rect 28641 9537 28675 9571
rect 29285 9537 29319 9571
rect 35909 9537 35943 9571
rect 10517 9469 10551 9503
rect 12081 9469 12115 9503
rect 13921 9469 13955 9503
rect 16037 9469 16071 9503
rect 16313 9469 16347 9503
rect 17417 9469 17451 9503
rect 20361 9469 20395 9503
rect 22477 9469 22511 9503
rect 24225 9469 24259 9503
rect 29193 9401 29227 9435
rect 9413 9333 9447 9367
rect 9965 9333 9999 9367
rect 14565 9333 14599 9367
rect 17680 9333 17714 9367
rect 21005 9333 21039 9367
rect 26065 9333 26099 9367
rect 27261 9333 27295 9367
rect 27905 9333 27939 9367
rect 28549 9333 28583 9367
rect 36093 9333 36127 9367
rect 9873 9129 9907 9163
rect 10517 9129 10551 9163
rect 11437 9129 11471 9163
rect 15485 9129 15519 9163
rect 19533 9129 19567 9163
rect 23397 9129 23431 9163
rect 30757 9129 30791 9163
rect 13277 9061 13311 9095
rect 14841 9061 14875 9095
rect 20177 9061 20211 9095
rect 9413 8993 9447 9027
rect 12725 8993 12759 9027
rect 16313 8993 16347 9027
rect 18521 8993 18555 9027
rect 20821 8993 20855 9027
rect 22845 8993 22879 9027
rect 24593 8993 24627 9027
rect 24869 8993 24903 9027
rect 27077 8993 27111 9027
rect 29929 8993 29963 9027
rect 31493 8993 31527 9027
rect 10425 8925 10459 8959
rect 11529 8925 11563 8959
rect 11989 8925 12023 8959
rect 14749 8925 14783 8959
rect 15393 8925 15427 8959
rect 16037 8925 16071 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 23489 8925 23523 8959
rect 29745 8925 29779 8959
rect 30665 8925 30699 8959
rect 12817 8857 12851 8891
rect 18061 8857 18095 8891
rect 22569 8857 22603 8891
rect 24041 8857 24075 8891
rect 26617 8857 26651 8891
rect 27353 8857 27387 8891
rect 31585 8857 31619 8891
rect 32137 8857 32171 8891
rect 12081 8789 12115 8823
rect 28825 8789 28859 8823
rect 11989 8585 12023 8619
rect 13369 8585 13403 8619
rect 13921 8585 13955 8619
rect 14565 8585 14599 8619
rect 21281 8585 21315 8619
rect 28273 8585 28307 8619
rect 10149 8517 10183 8551
rect 10701 8517 10735 8551
rect 10793 8517 10827 8551
rect 12817 8517 12851 8551
rect 16037 8517 16071 8551
rect 16865 8517 16899 8551
rect 23213 8517 23247 8551
rect 24961 8517 24995 8551
rect 1685 8449 1719 8483
rect 12081 8449 12115 8483
rect 14013 8449 14047 8483
rect 17417 8449 17451 8483
rect 20729 8449 20763 8483
rect 22937 8449 22971 8483
rect 27445 8449 27479 8483
rect 28365 8449 28399 8483
rect 29837 8449 29871 8483
rect 30297 8449 30331 8483
rect 31217 8449 31251 8483
rect 36093 8449 36127 8483
rect 16313 8381 16347 8415
rect 17509 8381 17543 8415
rect 18061 8381 18095 8415
rect 19809 8381 19843 8415
rect 20085 8381 20119 8415
rect 26249 8381 26283 8415
rect 29561 8381 29595 8415
rect 30481 8381 30515 8415
rect 1869 8313 1903 8347
rect 9689 8313 9723 8347
rect 20637 8313 20671 8347
rect 22293 8313 22327 8347
rect 25421 8313 25455 8347
rect 27353 8313 27387 8347
rect 36277 8313 36311 8347
rect 28825 8245 28859 8279
rect 31309 8245 31343 8279
rect 1593 8041 1627 8075
rect 10977 8041 11011 8075
rect 18521 8041 18555 8075
rect 19717 7973 19751 8007
rect 28365 7973 28399 8007
rect 17141 7905 17175 7939
rect 21465 7905 21499 7939
rect 21925 7905 21959 7939
rect 22201 7905 22235 7939
rect 24593 7905 24627 7939
rect 24869 7905 24903 7939
rect 27445 7905 27479 7939
rect 30021 7905 30055 7939
rect 6377 7837 6411 7871
rect 7021 7837 7055 7871
rect 11069 7837 11103 7871
rect 14473 7837 14507 7871
rect 15117 7837 15151 7871
rect 17785 7837 17819 7871
rect 18429 7837 18463 7871
rect 27537 7837 27571 7871
rect 28457 7837 28491 7871
rect 29101 7837 29135 7871
rect 29837 7837 29871 7871
rect 10425 7769 10459 7803
rect 11989 7769 12023 7803
rect 13737 7769 13771 7803
rect 15393 7769 15427 7803
rect 17877 7769 17911 7803
rect 21189 7769 21223 7803
rect 6561 7701 6595 7735
rect 14289 7701 14323 7735
rect 23673 7701 23707 7735
rect 26341 7701 26375 7735
rect 29009 7701 29043 7735
rect 13737 7497 13771 7531
rect 29193 7497 29227 7531
rect 1869 7429 1903 7463
rect 10425 7429 10459 7463
rect 10977 7429 11011 7463
rect 11069 7429 11103 7463
rect 12265 7429 12299 7463
rect 16313 7429 16347 7463
rect 17325 7429 17359 7463
rect 17969 7429 18003 7463
rect 20361 7429 20395 7463
rect 22017 7429 22051 7463
rect 22661 7429 22695 7463
rect 25697 7429 25731 7463
rect 36093 7429 36127 7463
rect 1685 7361 1719 7395
rect 14289 7361 14323 7395
rect 26617 7361 26651 7395
rect 27353 7361 27387 7395
rect 27997 7361 28031 7395
rect 28641 7361 28675 7395
rect 29285 7361 29319 7395
rect 29929 7361 29963 7395
rect 30389 7361 30423 7395
rect 35633 7361 35667 7395
rect 36277 7361 36311 7395
rect 11989 7293 12023 7327
rect 14565 7293 14599 7327
rect 20637 7293 20671 7327
rect 23213 7293 23247 7327
rect 23673 7293 23707 7327
rect 23949 7293 23983 7327
rect 26525 7293 26559 7327
rect 29837 7225 29871 7259
rect 18889 7157 18923 7191
rect 21281 7157 21315 7191
rect 27261 7157 27295 7191
rect 27905 7157 27939 7191
rect 28549 7157 28583 7191
rect 30481 7157 30515 7191
rect 1593 6953 1627 6987
rect 10517 6953 10551 6987
rect 12246 6953 12280 6987
rect 15196 6953 15230 6987
rect 9321 6817 9355 6851
rect 9965 6817 9999 6851
rect 11989 6817 12023 6851
rect 13737 6817 13771 6851
rect 14933 6817 14967 6851
rect 19533 6817 19567 6851
rect 20269 6817 20303 6851
rect 22293 6817 22327 6851
rect 24593 6817 24627 6851
rect 29837 6817 29871 6851
rect 10425 6749 10459 6783
rect 26341 6749 26375 6783
rect 27445 6749 27479 6783
rect 27537 6749 27571 6783
rect 28181 6749 28215 6783
rect 28825 6749 28859 6783
rect 29929 6749 29963 6783
rect 32505 6749 32539 6783
rect 9413 6681 9447 6715
rect 16957 6681 16991 6715
rect 18429 6681 18463 6715
rect 20545 6681 20579 6715
rect 26801 6681 26835 6715
rect 32781 6681 32815 6715
rect 11161 6613 11195 6647
rect 14473 6613 14507 6647
rect 17509 6613 17543 6647
rect 23213 6613 23247 6647
rect 23673 6613 23707 6647
rect 28089 6613 28123 6647
rect 28733 6613 28767 6647
rect 8493 6409 8527 6443
rect 9873 6409 9907 6443
rect 10609 6341 10643 6375
rect 19165 6341 19199 6375
rect 22293 6341 22327 6375
rect 24869 6341 24903 6375
rect 27813 6341 27847 6375
rect 8033 6273 8067 6307
rect 12357 6273 12391 6307
rect 17417 6273 17451 6307
rect 21373 6273 21407 6307
rect 22017 6273 22051 6307
rect 27905 6273 27939 6307
rect 29101 6273 29135 6307
rect 29745 6273 29779 6307
rect 30389 6273 30423 6307
rect 10517 6205 10551 6239
rect 12633 6205 12667 6239
rect 14565 6205 14599 6239
rect 16037 6205 16071 6239
rect 16313 6205 16347 6239
rect 19625 6205 19659 6239
rect 24041 6205 24075 6239
rect 24593 6205 24627 6239
rect 11069 6137 11103 6171
rect 14105 6137 14139 6171
rect 30297 6137 30331 6171
rect 7849 6069 7883 6103
rect 11805 6069 11839 6103
rect 16865 6069 16899 6103
rect 26341 6069 26375 6103
rect 27261 6069 27295 6103
rect 29009 6069 29043 6103
rect 29653 6069 29687 6103
rect 9229 5865 9263 5899
rect 11437 5865 11471 5899
rect 24593 5865 24627 5899
rect 26801 5865 26835 5899
rect 31769 5865 31803 5899
rect 14289 5797 14323 5831
rect 14933 5797 14967 5831
rect 18245 5797 18279 5831
rect 18705 5797 18739 5831
rect 11989 5729 12023 5763
rect 15577 5729 15611 5763
rect 17601 5729 17635 5763
rect 21005 5729 21039 5763
rect 22753 5729 22787 5763
rect 26341 5729 26375 5763
rect 9321 5661 9355 5695
rect 11529 5661 11563 5695
rect 23029 5661 23063 5695
rect 23765 5661 23799 5695
rect 30021 5661 30055 5695
rect 31677 5661 31711 5695
rect 12265 5593 12299 5627
rect 17325 5593 17359 5627
rect 26065 5593 26099 5627
rect 13737 5525 13771 5559
rect 19441 5525 19475 5559
rect 20545 5525 20579 5559
rect 23581 5525 23615 5559
rect 27353 5525 27387 5559
rect 29929 5525 29963 5559
rect 1777 5321 1811 5355
rect 11713 5321 11747 5355
rect 12265 5321 12299 5355
rect 16221 5321 16255 5355
rect 26341 5321 26375 5355
rect 9781 5253 9815 5287
rect 13737 5253 13771 5287
rect 14749 5253 14783 5287
rect 18153 5253 18187 5287
rect 1685 5185 1719 5219
rect 14013 5185 14047 5219
rect 17233 5185 17267 5219
rect 18981 5185 19015 5219
rect 21005 5185 21039 5219
rect 24593 5185 24627 5219
rect 29101 5185 29135 5219
rect 36093 5185 36127 5219
rect 9689 5117 9723 5151
rect 9965 5117 9999 5151
rect 14473 5117 14507 5151
rect 19257 5117 19291 5151
rect 23489 5117 23523 5151
rect 23765 5117 23799 5151
rect 24869 5117 24903 5151
rect 27169 5117 27203 5151
rect 27813 5117 27847 5151
rect 36369 5117 36403 5151
rect 11161 5049 11195 5083
rect 22017 4981 22051 5015
rect 29009 4981 29043 5015
rect 1593 4777 1627 4811
rect 9137 4777 9171 4811
rect 9781 4777 9815 4811
rect 10425 4777 10459 4811
rect 12449 4777 12483 4811
rect 18797 4777 18831 4811
rect 30849 4777 30883 4811
rect 36369 4777 36403 4811
rect 15209 4709 15243 4743
rect 18153 4709 18187 4743
rect 26801 4709 26835 4743
rect 14565 4641 14599 4675
rect 15669 4641 15703 4675
rect 17693 4641 17727 4675
rect 19993 4641 20027 4675
rect 24593 4641 24627 4675
rect 24869 4641 24903 4675
rect 9873 4573 9907 4607
rect 11437 4573 11471 4607
rect 13737 4573 13771 4607
rect 19717 4573 19751 4607
rect 22293 4573 22327 4607
rect 27537 4573 27571 4607
rect 28365 4573 28399 4607
rect 30757 4573 30791 4607
rect 10977 4505 11011 4539
rect 15945 4505 15979 4539
rect 22569 4505 22603 4539
rect 26985 4505 27019 4539
rect 21465 4437 21499 4471
rect 24041 4437 24075 4471
rect 26341 4437 26375 4471
rect 27721 4437 27755 4471
rect 28825 4437 28859 4471
rect 26525 4233 26559 4267
rect 12252 4165 12286 4199
rect 16037 4165 16071 4199
rect 19349 4165 19383 4199
rect 9413 4097 9447 4131
rect 10977 4097 11011 4131
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 19073 4097 19107 4131
rect 21097 4097 21131 4131
rect 23765 4097 23799 4131
rect 24225 4097 24259 4131
rect 26433 4097 26467 4131
rect 28917 4097 28951 4131
rect 30021 4097 30055 4131
rect 30757 4097 30791 4131
rect 31401 4097 31435 4131
rect 10517 4029 10551 4063
rect 11989 4029 12023 4063
rect 14565 4029 14599 4063
rect 17141 4029 17175 4063
rect 18613 4029 18647 4063
rect 23489 4029 23523 4063
rect 24501 4029 24535 4063
rect 25973 4029 26007 4063
rect 27169 4029 27203 4063
rect 28641 4029 28675 4063
rect 9965 3961 9999 3995
rect 35909 3961 35943 3995
rect 11069 3893 11103 3927
rect 13737 3893 13771 3927
rect 22017 3893 22051 3927
rect 29929 3893 29963 3927
rect 31217 3893 31251 3927
rect 9781 3689 9815 3723
rect 28549 3689 28583 3723
rect 31401 3689 31435 3723
rect 32045 3689 32079 3723
rect 19441 3621 19475 3655
rect 19993 3621 20027 3655
rect 29929 3621 29963 3655
rect 11253 3553 11287 3587
rect 12265 3553 12299 3587
rect 14381 3553 14415 3587
rect 18061 3553 18095 3587
rect 21741 3553 21775 3587
rect 22201 3553 22235 3587
rect 24593 3553 24627 3587
rect 24869 3553 24903 3587
rect 1869 3485 1903 3519
rect 9321 3485 9355 3519
rect 11529 3485 11563 3519
rect 11989 3485 12023 3519
rect 14289 3485 14323 3519
rect 14933 3485 14967 3519
rect 16037 3485 16071 3519
rect 18889 3485 18923 3519
rect 26801 3485 26835 3519
rect 29837 3485 29871 3519
rect 31493 3485 31527 3519
rect 32137 3485 32171 3519
rect 32781 3485 32815 3519
rect 35081 3485 35115 3519
rect 36093 3485 36127 3519
rect 16313 3417 16347 3451
rect 21465 3417 21499 3451
rect 22477 3417 22511 3451
rect 27077 3417 27111 3451
rect 30481 3417 30515 3451
rect 35173 3417 35207 3451
rect 1685 3349 1719 3383
rect 2421 3349 2455 3383
rect 8585 3349 8619 3383
rect 9137 3349 9171 3383
rect 13737 3349 13771 3383
rect 15117 3349 15151 3383
rect 18705 3349 18739 3383
rect 23949 3349 23983 3383
rect 26341 3349 26375 3383
rect 29009 3349 29043 3383
rect 32689 3349 32723 3383
rect 36277 3349 36311 3383
rect 8861 3145 8895 3179
rect 27445 3145 27479 3179
rect 32413 3145 32447 3179
rect 34437 3145 34471 3179
rect 9413 3077 9447 3111
rect 11161 3077 11195 3111
rect 13461 3077 13495 3111
rect 16037 3077 16071 3111
rect 22017 3077 22051 3111
rect 26525 3077 26559 3111
rect 28917 3077 28951 3111
rect 33057 3077 33091 3111
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 8769 3009 8803 3043
rect 13737 3009 13771 3043
rect 16313 3009 16347 3043
rect 16865 3009 16899 3043
rect 18061 3009 18095 3043
rect 18797 3009 18831 3043
rect 24041 3009 24075 3043
rect 24501 3009 24535 3043
rect 29745 3009 29779 3043
rect 31217 3009 31251 3043
rect 32505 3009 32539 3043
rect 32965 3009 32999 3043
rect 34989 3009 35023 3043
rect 35633 3009 35667 3043
rect 36277 3009 36311 3043
rect 7757 2941 7791 2975
rect 11989 2941 12023 2975
rect 19073 2941 19107 2975
rect 20821 2941 20855 2975
rect 21281 2941 21315 2975
rect 23765 2941 23799 2975
rect 24777 2941 24811 2975
rect 30021 2941 30055 2975
rect 31769 2941 31803 2975
rect 8309 2873 8343 2907
rect 33609 2873 33643 2907
rect 35449 2873 35483 2907
rect 1685 2805 1719 2839
rect 2329 2805 2363 2839
rect 2973 2805 3007 2839
rect 14565 2805 14599 2839
rect 17049 2805 17083 2839
rect 18245 2805 18279 2839
rect 31033 2805 31067 2839
rect 36185 2805 36219 2839
rect 2513 2601 2547 2635
rect 5365 2601 5399 2635
rect 28917 2601 28951 2635
rect 34253 2601 34287 2635
rect 4169 2533 4203 2567
rect 24593 2533 24627 2567
rect 11989 2465 12023 2499
rect 14565 2465 14599 2499
rect 17141 2465 17175 2499
rect 19441 2465 19475 2499
rect 21465 2465 21499 2499
rect 22109 2465 22143 2499
rect 26065 2465 26099 2499
rect 26341 2465 26375 2499
rect 27169 2465 27203 2499
rect 30297 2465 30331 2499
rect 30573 2465 30607 2499
rect 32321 2465 32355 2499
rect 1869 2397 1903 2431
rect 2329 2397 2363 2431
rect 3985 2397 4019 2431
rect 4905 2397 4939 2431
rect 6561 2397 6595 2431
rect 8125 2397 8159 2431
rect 9505 2397 9539 2431
rect 10425 2397 10459 2431
rect 10885 2397 10919 2431
rect 31309 2397 31343 2431
rect 32965 2397 32999 2431
rect 33241 2397 33275 2431
rect 34897 2397 34931 2431
rect 36093 2397 36127 2431
rect 9689 2329 9723 2363
rect 12265 2329 12299 2363
rect 14841 2329 14875 2363
rect 18889 2329 18923 2363
rect 19717 2329 19751 2363
rect 23765 2329 23799 2363
rect 27445 2329 27479 2363
rect 1685 2261 1719 2295
rect 3341 2261 3375 2295
rect 4721 2261 4755 2295
rect 6745 2261 6779 2295
rect 7389 2261 7423 2295
rect 7941 2261 7975 2295
rect 10241 2261 10275 2295
rect 11069 2261 11103 2295
rect 13737 2261 13771 2295
rect 16313 2261 16347 2295
rect 31125 2261 31159 2295
rect 35081 2261 35115 2295
rect 36277 2261 36311 2295
<< metal1 >>
rect 1104 37562 36892 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36892 37562
rect 1104 37488 36892 37510
rect 16114 37408 16120 37460
rect 16172 37448 16178 37460
rect 16209 37451 16267 37457
rect 16209 37448 16221 37451
rect 16172 37420 16221 37448
rect 16172 37408 16178 37420
rect 16209 37417 16221 37420
rect 16255 37448 16267 37451
rect 16255 37420 16574 37448
rect 16255 37417 16267 37420
rect 16209 37411 16267 37417
rect 2406 37312 2412 37324
rect 2367 37284 2412 37312
rect 2406 37272 2412 37284
rect 2464 37272 2470 37324
rect 9309 37315 9367 37321
rect 9309 37281 9321 37315
rect 9355 37312 9367 37315
rect 9355 37284 9720 37312
rect 9355 37281 9367 37284
rect 9309 37275 9367 37281
rect 9692 37256 9720 37284
rect 12434 37272 12440 37324
rect 12492 37312 12498 37324
rect 13265 37315 13323 37321
rect 13265 37312 13277 37315
rect 12492 37284 13277 37312
rect 12492 37272 12498 37284
rect 13265 37281 13277 37284
rect 13311 37281 13323 37315
rect 13265 37275 13323 37281
rect 2133 37247 2191 37253
rect 2133 37213 2145 37247
rect 2179 37213 2191 37247
rect 2133 37207 2191 37213
rect 3421 37247 3479 37253
rect 3421 37213 3433 37247
rect 3467 37244 3479 37247
rect 3510 37244 3516 37256
rect 3467 37216 3516 37244
rect 3467 37213 3479 37216
rect 3421 37207 3479 37213
rect 2148 37176 2176 37207
rect 3510 37204 3516 37216
rect 3568 37204 3574 37256
rect 4157 37247 4215 37253
rect 4157 37213 4169 37247
rect 4203 37244 4215 37247
rect 4614 37244 4620 37256
rect 4203 37216 4620 37244
rect 4203 37213 4215 37216
rect 4157 37207 4215 37213
rect 4614 37204 4620 37216
rect 4672 37244 4678 37256
rect 4709 37247 4767 37253
rect 4709 37244 4721 37247
rect 4672 37216 4721 37244
rect 4672 37204 4678 37216
rect 4709 37213 4721 37216
rect 4755 37213 4767 37247
rect 4709 37207 4767 37213
rect 5997 37247 6055 37253
rect 5997 37213 6009 37247
rect 6043 37244 6055 37247
rect 6454 37244 6460 37256
rect 6043 37216 6460 37244
rect 6043 37213 6055 37216
rect 5997 37207 6055 37213
rect 6454 37204 6460 37216
rect 6512 37244 6518 37256
rect 6641 37247 6699 37253
rect 6641 37244 6653 37247
rect 6512 37216 6653 37244
rect 6512 37204 6518 37216
rect 6641 37213 6653 37216
rect 6687 37213 6699 37247
rect 6641 37207 6699 37213
rect 7650 37204 7656 37256
rect 7708 37244 7714 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 7708 37216 7849 37244
rect 7708 37204 7714 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 7837 37207 7895 37213
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9732 37216 9873 37244
rect 9732 37204 9738 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 11977 37247 12035 37253
rect 11977 37213 11989 37247
rect 12023 37244 12035 37247
rect 12066 37244 12072 37256
rect 12023 37216 12072 37244
rect 12023 37213 12035 37216
rect 11977 37207 12035 37213
rect 12066 37204 12072 37216
rect 12124 37204 12130 37256
rect 12529 37247 12587 37253
rect 12529 37213 12541 37247
rect 12575 37244 12587 37247
rect 12894 37244 12900 37256
rect 12575 37216 12900 37244
rect 12575 37213 12587 37216
rect 12529 37207 12587 37213
rect 12894 37204 12900 37216
rect 12952 37244 12958 37256
rect 13081 37247 13139 37253
rect 13081 37244 13093 37247
rect 12952 37216 13093 37244
rect 12952 37204 12958 37216
rect 13081 37213 13093 37216
rect 13127 37213 13139 37247
rect 13081 37207 13139 37213
rect 15197 37247 15255 37253
rect 15197 37213 15209 37247
rect 15243 37244 15255 37247
rect 16546 37244 16574 37420
rect 26418 37408 26424 37460
rect 26476 37448 26482 37460
rect 26513 37451 26571 37457
rect 26513 37448 26525 37451
rect 26476 37420 26525 37448
rect 26476 37408 26482 37420
rect 26513 37417 26525 37420
rect 26559 37417 26571 37451
rect 26513 37411 26571 37417
rect 16666 37272 16672 37324
rect 16724 37312 16730 37324
rect 17129 37315 17187 37321
rect 17129 37312 17141 37315
rect 16724 37284 17141 37312
rect 16724 37272 16730 37284
rect 17129 37281 17141 37284
rect 17175 37281 17187 37315
rect 17129 37275 17187 37281
rect 19334 37272 19340 37324
rect 19392 37312 19398 37324
rect 19429 37315 19487 37321
rect 19429 37312 19441 37315
rect 19392 37284 19441 37312
rect 19392 37272 19398 37284
rect 19429 37281 19441 37284
rect 19475 37281 19487 37315
rect 26528 37312 26556 37411
rect 27157 37315 27215 37321
rect 27157 37312 27169 37315
rect 26528 37284 27169 37312
rect 19429 37275 19487 37281
rect 27157 37281 27169 37284
rect 27203 37281 27215 37315
rect 27157 37275 27215 37281
rect 16945 37247 17003 37253
rect 16945 37244 16957 37247
rect 15243 37216 15700 37244
rect 16546 37216 16957 37244
rect 15243 37213 15255 37216
rect 15197 37207 15255 37213
rect 2148 37148 12572 37176
rect 12544 37120 12572 37148
rect 15672 37120 15700 37216
rect 16945 37213 16957 37216
rect 16991 37213 17003 37247
rect 16945 37207 17003 37213
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37244 18475 37247
rect 18506 37244 18512 37256
rect 18463 37216 18512 37244
rect 18463 37213 18475 37216
rect 18417 37207 18475 37213
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 19705 37247 19763 37253
rect 19705 37213 19717 37247
rect 19751 37244 19763 37247
rect 19978 37244 19984 37256
rect 19751 37216 19984 37244
rect 19751 37213 19763 37216
rect 19705 37207 19763 37213
rect 19978 37204 19984 37216
rect 20036 37204 20042 37256
rect 22002 37244 22008 37256
rect 21963 37216 22008 37244
rect 22002 37204 22008 37216
rect 22060 37204 22066 37256
rect 22738 37244 22744 37256
rect 22699 37216 22744 37244
rect 22738 37204 22744 37216
rect 22796 37204 22802 37256
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 27430 37244 27436 37256
rect 27391 37216 27436 37244
rect 27430 37204 27436 37216
rect 27488 37204 27494 37256
rect 28442 37244 28448 37256
rect 28403 37216 28448 37244
rect 28442 37204 28448 37216
rect 28500 37204 28506 37256
rect 29914 37204 29920 37256
rect 29972 37244 29978 37256
rect 30009 37247 30067 37253
rect 30009 37244 30021 37247
rect 29972 37216 30021 37244
rect 29972 37204 29978 37216
rect 30009 37213 30021 37216
rect 30055 37213 30067 37247
rect 31018 37244 31024 37256
rect 30979 37216 31024 37244
rect 30009 37207 30067 37213
rect 31018 37204 31024 37216
rect 31076 37204 31082 37256
rect 32953 37247 33011 37253
rect 32953 37213 32965 37247
rect 32999 37213 33011 37247
rect 32953 37207 33011 37213
rect 27338 37136 27344 37188
rect 27396 37176 27402 37188
rect 32968 37176 32996 37207
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35161 37247 35219 37253
rect 35161 37244 35173 37247
rect 34848 37216 35173 37244
rect 34848 37204 34854 37216
rect 35161 37213 35173 37216
rect 35207 37213 35219 37247
rect 36078 37244 36084 37256
rect 36039 37216 36084 37244
rect 35161 37207 35219 37213
rect 36078 37204 36084 37216
rect 36136 37204 36142 37256
rect 27396 37148 32996 37176
rect 27396 37136 27402 37148
rect 3234 37108 3240 37120
rect 3195 37080 3240 37108
rect 3234 37068 3240 37080
rect 3292 37068 3298 37120
rect 4798 37108 4804 37120
rect 4759 37080 4804 37108
rect 4798 37068 4804 37080
rect 4856 37068 4862 37120
rect 6730 37108 6736 37120
rect 6691 37080 6736 37108
rect 6730 37068 6736 37080
rect 6788 37068 6794 37120
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 9950 37108 9956 37120
rect 9911 37080 9956 37108
rect 8021 37071 8079 37077
rect 9950 37068 9956 37080
rect 10008 37068 10014 37120
rect 11054 37068 11060 37120
rect 11112 37108 11118 37120
rect 11793 37111 11851 37117
rect 11793 37108 11805 37111
rect 11112 37080 11805 37108
rect 11112 37068 11118 37080
rect 11793 37077 11805 37080
rect 11839 37077 11851 37111
rect 11793 37071 11851 37077
rect 12526 37068 12532 37120
rect 12584 37068 12590 37120
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 15013 37111 15071 37117
rect 15013 37108 15025 37111
rect 14884 37080 15025 37108
rect 14884 37068 14890 37080
rect 15013 37077 15025 37080
rect 15059 37077 15071 37111
rect 15654 37108 15660 37120
rect 15615 37080 15660 37108
rect 15013 37071 15071 37077
rect 15654 37068 15660 37080
rect 15712 37068 15718 37120
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18233 37111 18291 37117
rect 18233 37108 18245 37111
rect 18104 37080 18245 37108
rect 18104 37068 18110 37080
rect 18233 37077 18245 37080
rect 18279 37077 18291 37111
rect 18233 37071 18291 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 22554 37068 22560 37120
rect 22612 37108 22618 37120
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22612 37080 22937 37108
rect 22612 37068 22618 37080
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 22925 37071 22983 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 28629 37111 28687 37117
rect 28629 37108 28641 37111
rect 27764 37080 28641 37108
rect 27764 37068 27770 37080
rect 28629 37077 28641 37080
rect 28675 37077 28687 37111
rect 28629 37071 28687 37077
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 29825 37111 29883 37117
rect 29825 37108 29837 37111
rect 29696 37080 29837 37108
rect 29696 37068 29702 37080
rect 29825 37077 29837 37080
rect 29871 37077 29883 37111
rect 29825 37071 29883 37077
rect 30926 37068 30932 37120
rect 30984 37108 30990 37120
rect 31205 37111 31263 37117
rect 31205 37108 31217 37111
rect 30984 37080 31217 37108
rect 30984 37068 30990 37080
rect 31205 37077 31217 37080
rect 31251 37077 31263 37111
rect 33134 37108 33140 37120
rect 33095 37080 33140 37108
rect 31205 37071 31263 37077
rect 33134 37068 33140 37080
rect 33192 37068 33198 37120
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 34977 37111 35035 37117
rect 34977 37108 34989 37111
rect 34572 37080 34989 37108
rect 34572 37068 34578 37080
rect 34977 37077 34989 37080
rect 35023 37077 35035 37111
rect 34977 37071 35035 37077
rect 36170 37068 36176 37120
rect 36228 37108 36234 37120
rect 36265 37111 36323 37117
rect 36265 37108 36277 37111
rect 36228 37080 36277 37108
rect 36228 37068 36234 37080
rect 36265 37077 36277 37080
rect 36311 37077 36323 37111
rect 36265 37071 36323 37077
rect 1104 37018 36892 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 36892 37018
rect 1104 36944 36892 36966
rect 2501 36907 2559 36913
rect 2501 36873 2513 36907
rect 2547 36904 2559 36907
rect 2774 36904 2780 36916
rect 2547 36876 2780 36904
rect 2547 36873 2559 36876
rect 2501 36867 2559 36873
rect 2774 36864 2780 36876
rect 2832 36864 2838 36916
rect 7650 36904 7656 36916
rect 7611 36876 7656 36904
rect 7650 36864 7656 36876
rect 7708 36864 7714 36916
rect 12066 36904 12072 36916
rect 12027 36876 12072 36904
rect 12066 36864 12072 36876
rect 12124 36864 12130 36916
rect 19334 36904 19340 36916
rect 19295 36876 19340 36904
rect 19334 36864 19340 36876
rect 19392 36864 19398 36916
rect 27338 36904 27344 36916
rect 27299 36876 27344 36904
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 29825 36907 29883 36913
rect 29825 36873 29837 36907
rect 29871 36904 29883 36907
rect 31018 36904 31024 36916
rect 29871 36876 31024 36904
rect 29871 36873 29883 36876
rect 29825 36867 29883 36873
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 35526 36904 35532 36916
rect 35487 36876 35532 36904
rect 35526 36864 35532 36876
rect 35584 36864 35590 36916
rect 36265 36907 36323 36913
rect 36265 36873 36277 36907
rect 36311 36904 36323 36907
rect 37366 36904 37372 36916
rect 36311 36876 37372 36904
rect 36311 36873 36323 36876
rect 36265 36867 36323 36873
rect 37366 36864 37372 36876
rect 37424 36864 37430 36916
rect 1302 36796 1308 36848
rect 1360 36836 1366 36848
rect 1673 36839 1731 36845
rect 1673 36836 1685 36839
rect 1360 36808 1685 36836
rect 1360 36796 1366 36808
rect 1673 36805 1685 36808
rect 1719 36805 1731 36839
rect 1673 36799 1731 36805
rect 1946 36728 1952 36780
rect 2004 36768 2010 36780
rect 2317 36771 2375 36777
rect 2317 36768 2329 36771
rect 2004 36740 2329 36768
rect 2004 36728 2010 36740
rect 2317 36737 2329 36740
rect 2363 36737 2375 36771
rect 2317 36731 2375 36737
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 8294 36768 8300 36780
rect 7883 36740 8300 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 12253 36771 12311 36777
rect 12253 36737 12265 36771
rect 12299 36768 12311 36771
rect 12526 36768 12532 36780
rect 12299 36740 12532 36768
rect 12299 36737 12311 36740
rect 12253 36731 12311 36737
rect 12526 36728 12532 36740
rect 12584 36768 12590 36780
rect 12713 36771 12771 36777
rect 12713 36768 12725 36771
rect 12584 36740 12725 36768
rect 12584 36728 12590 36740
rect 12713 36737 12725 36740
rect 12759 36768 12771 36771
rect 13170 36768 13176 36780
rect 12759 36740 13176 36768
rect 12759 36737 12771 36740
rect 12713 36731 12771 36737
rect 13170 36728 13176 36740
rect 13228 36728 13234 36780
rect 19978 36728 19984 36780
rect 20036 36768 20042 36780
rect 20254 36768 20260 36780
rect 20036 36740 20260 36768
rect 20036 36728 20042 36740
rect 20254 36728 20260 36740
rect 20312 36768 20318 36780
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 20312 36740 27169 36768
rect 20312 36728 20318 36740
rect 27157 36737 27169 36740
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 28350 36728 28356 36780
rect 28408 36768 28414 36780
rect 29733 36771 29791 36777
rect 29733 36768 29745 36771
rect 28408 36740 29745 36768
rect 28408 36728 28414 36740
rect 29733 36737 29745 36740
rect 29779 36768 29791 36771
rect 30377 36771 30435 36777
rect 30377 36768 30389 36771
rect 29779 36740 30389 36768
rect 29779 36737 29791 36740
rect 29733 36731 29791 36737
rect 30377 36737 30389 36740
rect 30423 36737 30435 36771
rect 30377 36731 30435 36737
rect 34885 36771 34943 36777
rect 34885 36737 34897 36771
rect 34931 36768 34943 36771
rect 35345 36771 35403 36777
rect 35345 36768 35357 36771
rect 34931 36740 35357 36768
rect 34931 36737 34943 36740
rect 34885 36731 34943 36737
rect 35345 36737 35357 36740
rect 35391 36768 35403 36771
rect 35986 36768 35992 36780
rect 35391 36740 35992 36768
rect 35391 36737 35403 36740
rect 35345 36731 35403 36737
rect 35986 36728 35992 36740
rect 36044 36728 36050 36780
rect 36081 36771 36139 36777
rect 36081 36737 36093 36771
rect 36127 36737 36139 36771
rect 36081 36731 36139 36737
rect 35894 36660 35900 36712
rect 35952 36700 35958 36712
rect 36096 36700 36124 36731
rect 35952 36672 36124 36700
rect 35952 36660 35958 36672
rect 1857 36635 1915 36641
rect 1857 36601 1869 36635
rect 1903 36632 1915 36635
rect 2590 36632 2596 36644
rect 1903 36604 2596 36632
rect 1903 36601 1915 36604
rect 1857 36595 1915 36601
rect 2590 36592 2596 36604
rect 2648 36592 2654 36644
rect 3510 36564 3516 36576
rect 3471 36536 3516 36564
rect 3510 36524 3516 36536
rect 3568 36524 3574 36576
rect 8294 36564 8300 36576
rect 8255 36536 8300 36564
rect 8294 36524 8300 36536
rect 8352 36524 8358 36576
rect 18506 36564 18512 36576
rect 18467 36536 18512 36564
rect 18506 36524 18512 36536
rect 18564 36524 18570 36576
rect 1104 36474 36892 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36892 36474
rect 1104 36400 36892 36422
rect 1302 36320 1308 36372
rect 1360 36360 1366 36372
rect 2317 36363 2375 36369
rect 2317 36360 2329 36363
rect 1360 36332 2329 36360
rect 1360 36320 1366 36332
rect 2317 36329 2329 36332
rect 2363 36329 2375 36363
rect 2317 36323 2375 36329
rect 35069 36159 35127 36165
rect 35069 36125 35081 36159
rect 35115 36156 35127 36159
rect 35526 36156 35532 36168
rect 35115 36128 35532 36156
rect 35115 36125 35127 36128
rect 35069 36119 35127 36125
rect 35526 36116 35532 36128
rect 35584 36116 35590 36168
rect 35802 36156 35808 36168
rect 35763 36128 35808 36156
rect 35802 36116 35808 36128
rect 35860 36116 35866 36168
rect 1670 36088 1676 36100
rect 1631 36060 1676 36088
rect 1670 36048 1676 36060
rect 1728 36048 1734 36100
rect 1857 36091 1915 36097
rect 1857 36057 1869 36091
rect 1903 36088 1915 36091
rect 1903 36060 6914 36088
rect 1903 36057 1915 36060
rect 1857 36051 1915 36057
rect 6886 36020 6914 36060
rect 17586 36020 17592 36032
rect 6886 35992 17592 36020
rect 17586 35980 17592 35992
rect 17644 35980 17650 36032
rect 1104 35930 36892 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 36892 35930
rect 1104 35856 36892 35878
rect 1670 35816 1676 35828
rect 1631 35788 1676 35816
rect 1670 35776 1676 35788
rect 1728 35776 1734 35828
rect 2225 35819 2283 35825
rect 2225 35785 2237 35819
rect 2271 35816 2283 35819
rect 2406 35816 2412 35828
rect 2271 35788 2412 35816
rect 2271 35785 2283 35788
rect 2225 35779 2283 35785
rect 2406 35776 2412 35788
rect 2464 35776 2470 35828
rect 27341 35819 27399 35825
rect 27341 35785 27353 35819
rect 27387 35816 27399 35819
rect 28442 35816 28448 35828
rect 27387 35788 28448 35816
rect 27387 35785 27399 35788
rect 27341 35779 27399 35785
rect 28442 35776 28448 35788
rect 28500 35776 28506 35828
rect 36078 35816 36084 35828
rect 36039 35788 36084 35816
rect 36078 35776 36084 35788
rect 36136 35776 36142 35828
rect 27154 35680 27160 35692
rect 27115 35652 27160 35680
rect 27154 35640 27160 35652
rect 27212 35680 27218 35692
rect 27801 35683 27859 35689
rect 27801 35680 27813 35683
rect 27212 35652 27813 35680
rect 27212 35640 27218 35652
rect 27801 35649 27813 35652
rect 27847 35649 27859 35683
rect 27801 35643 27859 35649
rect 34514 35640 34520 35692
rect 34572 35680 34578 35692
rect 35802 35680 35808 35692
rect 34572 35652 35808 35680
rect 34572 35640 34578 35652
rect 35802 35640 35808 35652
rect 35860 35680 35866 35692
rect 35897 35683 35955 35689
rect 35897 35680 35909 35683
rect 35860 35652 35909 35680
rect 35860 35640 35866 35652
rect 35897 35649 35909 35652
rect 35943 35649 35955 35683
rect 35897 35643 35955 35649
rect 1104 35386 36892 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36892 35386
rect 1104 35312 36892 35334
rect 20993 35275 21051 35281
rect 20993 35241 21005 35275
rect 21039 35272 21051 35275
rect 22002 35272 22008 35284
rect 21039 35244 22008 35272
rect 21039 35241 21051 35244
rect 20993 35235 21051 35241
rect 22002 35232 22008 35244
rect 22060 35232 22066 35284
rect 1857 35071 1915 35077
rect 1857 35037 1869 35071
rect 1903 35068 1915 35071
rect 7558 35068 7564 35080
rect 1903 35040 7564 35068
rect 1903 35037 1915 35040
rect 1857 35031 1915 35037
rect 7558 35028 7564 35040
rect 7616 35028 7622 35080
rect 20809 35071 20867 35077
rect 20809 35037 20821 35071
rect 20855 35068 20867 35071
rect 20855 35040 21588 35068
rect 20855 35037 20867 35040
rect 20809 35031 20867 35037
rect 1670 34932 1676 34944
rect 1631 34904 1676 34932
rect 1670 34892 1676 34904
rect 1728 34892 1734 34944
rect 21560 34941 21588 35040
rect 26602 35028 26608 35080
rect 26660 35068 26666 35080
rect 36081 35071 36139 35077
rect 36081 35068 36093 35071
rect 26660 35040 36093 35068
rect 26660 35028 26666 35040
rect 36081 35037 36093 35040
rect 36127 35037 36139 35071
rect 36354 35068 36360 35080
rect 36315 35040 36360 35068
rect 36081 35031 36139 35037
rect 36354 35028 36360 35040
rect 36412 35028 36418 35080
rect 21545 34935 21603 34941
rect 21545 34901 21557 34935
rect 21591 34932 21603 34935
rect 24394 34932 24400 34944
rect 21591 34904 24400 34932
rect 21591 34901 21603 34904
rect 21545 34895 21603 34901
rect 24394 34892 24400 34904
rect 24452 34892 24458 34944
rect 1104 34842 36892 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 36892 34842
rect 1104 34768 36892 34790
rect 36354 34728 36360 34740
rect 36315 34700 36360 34728
rect 36354 34688 36360 34700
rect 36412 34688 36418 34740
rect 24394 34484 24400 34536
rect 24452 34524 24458 34536
rect 36078 34524 36084 34536
rect 24452 34496 36084 34524
rect 24452 34484 24458 34496
rect 36078 34484 36084 34496
rect 36136 34484 36142 34536
rect 1104 34298 36892 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36892 34298
rect 1104 34224 36892 34246
rect 1104 33754 36892 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 36892 33754
rect 1104 33680 36892 33702
rect 1104 33210 36892 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36892 33210
rect 1104 33136 36892 33158
rect 27154 32852 27160 32904
rect 27212 32892 27218 32904
rect 36081 32895 36139 32901
rect 36081 32892 36093 32895
rect 27212 32864 36093 32892
rect 27212 32852 27218 32864
rect 36081 32861 36093 32864
rect 36127 32861 36139 32895
rect 36354 32892 36360 32904
rect 36315 32864 36360 32892
rect 36081 32855 36139 32861
rect 36354 32852 36360 32864
rect 36412 32852 36418 32904
rect 1670 32824 1676 32836
rect 1631 32796 1676 32824
rect 1670 32784 1676 32796
rect 1728 32784 1734 32836
rect 1857 32827 1915 32833
rect 1857 32793 1869 32827
rect 1903 32824 1915 32827
rect 2222 32824 2228 32836
rect 1903 32796 2228 32824
rect 1903 32793 1915 32796
rect 1857 32787 1915 32793
rect 2222 32784 2228 32796
rect 2280 32784 2286 32836
rect 1104 32666 36892 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 36892 32666
rect 1104 32592 36892 32614
rect 1670 32552 1676 32564
rect 1631 32524 1676 32552
rect 1670 32512 1676 32524
rect 1728 32512 1734 32564
rect 22189 32555 22247 32561
rect 22189 32521 22201 32555
rect 22235 32552 22247 32555
rect 22738 32552 22744 32564
rect 22235 32524 22744 32552
rect 22235 32521 22247 32524
rect 22189 32515 22247 32521
rect 22738 32512 22744 32524
rect 22796 32512 22802 32564
rect 36354 32552 36360 32564
rect 36315 32524 36360 32552
rect 36354 32512 36360 32524
rect 36412 32512 36418 32564
rect 22002 32416 22008 32428
rect 21963 32388 22008 32416
rect 22002 32376 22008 32388
rect 22060 32416 22066 32428
rect 22649 32419 22707 32425
rect 22649 32416 22661 32419
rect 22060 32388 22661 32416
rect 22060 32376 22066 32388
rect 22649 32385 22661 32388
rect 22695 32385 22707 32419
rect 22649 32379 22707 32385
rect 1104 32122 36892 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36892 32122
rect 1104 32048 36892 32070
rect 36078 31940 36084 31952
rect 36039 31912 36084 31940
rect 36078 31900 36084 31912
rect 36136 31900 36142 31952
rect 1857 31807 1915 31813
rect 1857 31773 1869 31807
rect 1903 31804 1915 31807
rect 22002 31804 22008 31816
rect 1903 31776 22008 31804
rect 1903 31773 1915 31776
rect 1857 31767 1915 31773
rect 22002 31764 22008 31776
rect 22060 31764 22066 31816
rect 35621 31807 35679 31813
rect 35621 31773 35633 31807
rect 35667 31804 35679 31807
rect 35802 31804 35808 31816
rect 35667 31776 35808 31804
rect 35667 31773 35679 31776
rect 35621 31767 35679 31773
rect 35802 31764 35808 31776
rect 35860 31804 35866 31816
rect 36265 31807 36323 31813
rect 36265 31804 36277 31807
rect 35860 31776 36277 31804
rect 35860 31764 35866 31776
rect 36265 31773 36277 31776
rect 36311 31773 36323 31807
rect 36265 31767 36323 31773
rect 1578 31696 1584 31748
rect 1636 31736 1642 31748
rect 1673 31739 1731 31745
rect 1673 31736 1685 31739
rect 1636 31708 1685 31736
rect 1636 31696 1642 31708
rect 1673 31705 1685 31708
rect 1719 31705 1731 31739
rect 1673 31699 1731 31705
rect 1104 31578 36892 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 36892 31578
rect 1104 31504 36892 31526
rect 29457 31467 29515 31473
rect 29457 31433 29469 31467
rect 29503 31464 29515 31467
rect 35894 31464 35900 31476
rect 29503 31436 35900 31464
rect 29503 31433 29515 31436
rect 29457 31427 29515 31433
rect 35894 31424 35900 31436
rect 35952 31424 35958 31476
rect 1578 31396 1584 31408
rect 1539 31368 1584 31396
rect 1578 31356 1584 31368
rect 1636 31356 1642 31408
rect 29273 31331 29331 31337
rect 29273 31297 29285 31331
rect 29319 31328 29331 31331
rect 29822 31328 29828 31340
rect 29319 31300 29828 31328
rect 29319 31297 29331 31300
rect 29273 31291 29331 31297
rect 29822 31288 29828 31300
rect 29880 31288 29886 31340
rect 29822 31084 29828 31136
rect 29880 31124 29886 31136
rect 29917 31127 29975 31133
rect 29917 31124 29929 31127
rect 29880 31096 29929 31124
rect 29880 31084 29886 31096
rect 29917 31093 29929 31096
rect 29963 31093 29975 31127
rect 29917 31087 29975 31093
rect 1104 31034 36892 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36892 31034
rect 1104 30960 36892 30982
rect 1104 30490 36892 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 36892 30490
rect 1104 30416 36892 30438
rect 29914 30308 29920 30320
rect 29875 30280 29920 30308
rect 29914 30268 29920 30280
rect 29972 30268 29978 30320
rect 24118 30200 24124 30252
rect 24176 30240 24182 30252
rect 30009 30243 30067 30249
rect 30009 30240 30021 30243
rect 24176 30212 30021 30240
rect 24176 30200 24182 30212
rect 30009 30209 30021 30212
rect 30055 30240 30067 30243
rect 30469 30243 30527 30249
rect 30469 30240 30481 30243
rect 30055 30212 30481 30240
rect 30055 30209 30067 30212
rect 30009 30203 30067 30209
rect 30469 30209 30481 30212
rect 30515 30209 30527 30243
rect 30469 30203 30527 30209
rect 1104 29946 36892 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36892 29946
rect 1104 29872 36892 29894
rect 23937 29835 23995 29841
rect 23937 29801 23949 29835
rect 23983 29832 23995 29835
rect 24578 29832 24584 29844
rect 23983 29804 24584 29832
rect 23983 29801 23995 29804
rect 23937 29795 23995 29801
rect 24578 29792 24584 29804
rect 24636 29792 24642 29844
rect 34790 29792 34796 29844
rect 34848 29832 34854 29844
rect 34977 29835 35035 29841
rect 34977 29832 34989 29835
rect 34848 29804 34989 29832
rect 34848 29792 34854 29804
rect 34977 29801 34989 29804
rect 35023 29801 35035 29835
rect 34977 29795 35035 29801
rect 23753 29631 23811 29637
rect 23753 29597 23765 29631
rect 23799 29628 23811 29631
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 23799 29600 24532 29628
rect 23799 29597 23811 29600
rect 23753 29591 23811 29597
rect 1578 29520 1584 29572
rect 1636 29560 1642 29572
rect 1673 29563 1731 29569
rect 1673 29560 1685 29563
rect 1636 29532 1685 29560
rect 1636 29520 1642 29532
rect 1673 29529 1685 29532
rect 1719 29529 1731 29563
rect 1673 29523 1731 29529
rect 1857 29563 1915 29569
rect 1857 29529 1869 29563
rect 1903 29560 1915 29563
rect 2038 29560 2044 29572
rect 1903 29532 2044 29560
rect 1903 29529 1915 29532
rect 1857 29523 1915 29529
rect 2038 29520 2044 29532
rect 2096 29520 2102 29572
rect 24504 29504 24532 29600
rect 26206 29600 34897 29628
rect 24486 29452 24492 29504
rect 24544 29492 24550 29504
rect 24581 29495 24639 29501
rect 24581 29492 24593 29495
rect 24544 29464 24593 29492
rect 24544 29452 24550 29464
rect 24581 29461 24593 29464
rect 24627 29461 24639 29495
rect 24581 29455 24639 29461
rect 25590 29452 25596 29504
rect 25648 29492 25654 29504
rect 26206 29492 26234 29600
rect 34885 29597 34897 29600
rect 34931 29628 34943 29631
rect 35529 29631 35587 29637
rect 35529 29628 35541 29631
rect 34931 29600 35541 29628
rect 34931 29597 34943 29600
rect 34885 29591 34943 29597
rect 35529 29597 35541 29600
rect 35575 29597 35587 29631
rect 35529 29591 35587 29597
rect 29730 29520 29736 29572
rect 29788 29560 29794 29572
rect 36081 29563 36139 29569
rect 36081 29560 36093 29563
rect 29788 29532 36093 29560
rect 29788 29520 29794 29532
rect 36081 29529 36093 29532
rect 36127 29529 36139 29563
rect 36081 29523 36139 29529
rect 36265 29563 36323 29569
rect 36265 29529 36277 29563
rect 36311 29560 36323 29563
rect 36354 29560 36360 29572
rect 36311 29532 36360 29560
rect 36311 29529 36323 29532
rect 36265 29523 36323 29529
rect 36354 29520 36360 29532
rect 36412 29520 36418 29572
rect 25648 29464 26234 29492
rect 25648 29452 25654 29464
rect 1104 29402 36892 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 36892 29402
rect 1104 29328 36892 29350
rect 1578 29288 1584 29300
rect 1539 29260 1584 29288
rect 1578 29248 1584 29260
rect 1636 29248 1642 29300
rect 36354 29288 36360 29300
rect 36315 29260 36360 29288
rect 36354 29248 36360 29260
rect 36412 29248 36418 29300
rect 1104 28858 36892 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36892 28858
rect 1104 28784 36892 28806
rect 1104 28314 36892 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 36892 28314
rect 1104 28240 36892 28262
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28064 1915 28067
rect 2314 28064 2320 28076
rect 1903 28036 2320 28064
rect 1903 28033 1915 28036
rect 1857 28027 1915 28033
rect 2314 28024 2320 28036
rect 2372 28024 2378 28076
rect 13170 28064 13176 28076
rect 13131 28036 13176 28064
rect 13170 28024 13176 28036
rect 13228 28064 13234 28076
rect 13817 28067 13875 28073
rect 13817 28064 13829 28067
rect 13228 28036 13829 28064
rect 13228 28024 13234 28036
rect 13817 28033 13829 28036
rect 13863 28033 13875 28067
rect 20254 28064 20260 28076
rect 20215 28036 20260 28064
rect 13817 28027 13875 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 35621 28067 35679 28073
rect 35621 28033 35633 28067
rect 35667 28064 35679 28067
rect 36262 28064 36268 28076
rect 35667 28036 36268 28064
rect 35667 28033 35679 28036
rect 35621 28027 35679 28033
rect 36262 28024 36268 28036
rect 36320 28024 36326 28076
rect 1670 27928 1676 27940
rect 1631 27900 1676 27928
rect 1670 27888 1676 27900
rect 1728 27888 1734 27940
rect 13265 27931 13323 27937
rect 13265 27897 13277 27931
rect 13311 27928 13323 27931
rect 14090 27928 14096 27940
rect 13311 27900 14096 27928
rect 13311 27897 13323 27900
rect 13265 27891 13323 27897
rect 14090 27888 14096 27900
rect 14148 27888 14154 27940
rect 35342 27888 35348 27940
rect 35400 27928 35406 27940
rect 36081 27931 36139 27937
rect 36081 27928 36093 27931
rect 35400 27900 36093 27928
rect 35400 27888 35406 27900
rect 36081 27897 36093 27900
rect 36127 27897 36139 27931
rect 36081 27891 36139 27897
rect 2314 27860 2320 27872
rect 2275 27832 2320 27860
rect 2314 27820 2320 27832
rect 2372 27820 2378 27872
rect 20349 27863 20407 27869
rect 20349 27829 20361 27863
rect 20395 27860 20407 27863
rect 21450 27860 21456 27872
rect 20395 27832 21456 27860
rect 20395 27829 20407 27832
rect 20349 27823 20407 27829
rect 21450 27820 21456 27832
rect 21508 27820 21514 27872
rect 1104 27770 36892 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36892 27770
rect 1104 27696 36892 27718
rect 7558 27588 7564 27600
rect 7519 27560 7564 27588
rect 7558 27548 7564 27560
rect 7616 27548 7622 27600
rect 3510 27480 3516 27532
rect 3568 27520 3574 27532
rect 11977 27523 12035 27529
rect 11977 27520 11989 27523
rect 3568 27492 11989 27520
rect 3568 27480 3574 27492
rect 11977 27489 11989 27492
rect 12023 27489 12035 27523
rect 11977 27483 12035 27489
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27452 7711 27455
rect 12069 27455 12127 27461
rect 7699 27424 8156 27452
rect 7699 27421 7711 27424
rect 7653 27415 7711 27421
rect 8128 27328 8156 27424
rect 12069 27421 12081 27455
rect 12115 27452 12127 27455
rect 14458 27452 14464 27464
rect 12115 27424 14464 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27452 29975 27455
rect 34514 27452 34520 27464
rect 29963 27424 34520 27452
rect 29963 27421 29975 27424
rect 29917 27415 29975 27421
rect 34514 27412 34520 27424
rect 34572 27412 34578 27464
rect 8110 27316 8116 27328
rect 8071 27288 8116 27316
rect 8110 27276 8116 27288
rect 8168 27276 8174 27328
rect 25498 27276 25504 27328
rect 25556 27316 25562 27328
rect 29825 27319 29883 27325
rect 29825 27316 29837 27319
rect 25556 27288 29837 27316
rect 25556 27276 25562 27288
rect 29825 27285 29837 27288
rect 29871 27285 29883 27319
rect 29825 27279 29883 27285
rect 1104 27226 36892 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 36892 27226
rect 1104 27152 36892 27174
rect 1104 26682 36892 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36892 26682
rect 1104 26608 36892 26630
rect 25685 26571 25743 26577
rect 25685 26537 25697 26571
rect 25731 26568 25743 26571
rect 27154 26568 27160 26580
rect 25731 26540 27160 26568
rect 25731 26537 25743 26540
rect 25685 26531 25743 26537
rect 1857 26367 1915 26373
rect 1857 26333 1869 26367
rect 1903 26364 1915 26367
rect 25133 26367 25191 26373
rect 1903 26336 2452 26364
rect 1903 26333 1915 26336
rect 1857 26327 1915 26333
rect 2424 26308 2452 26336
rect 25133 26333 25145 26367
rect 25179 26364 25191 26367
rect 25700 26364 25728 26531
rect 27154 26528 27160 26540
rect 27212 26528 27218 26580
rect 35802 26460 35808 26512
rect 35860 26500 35866 26512
rect 36265 26503 36323 26509
rect 36265 26500 36277 26503
rect 35860 26472 36277 26500
rect 35860 26460 35866 26472
rect 36265 26469 36277 26472
rect 36311 26469 36323 26503
rect 36265 26463 36323 26469
rect 36078 26364 36084 26376
rect 25179 26336 25728 26364
rect 36039 26336 36084 26364
rect 25179 26333 25191 26336
rect 25133 26327 25191 26333
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 2406 26296 2412 26308
rect 2367 26268 2412 26296
rect 2406 26256 2412 26268
rect 2464 26256 2470 26308
rect 21910 26256 21916 26308
rect 21968 26296 21974 26308
rect 25041 26299 25099 26305
rect 25041 26296 25053 26299
rect 21968 26268 25053 26296
rect 21968 26256 21974 26268
rect 25041 26265 25053 26268
rect 25087 26265 25099 26299
rect 25041 26259 25099 26265
rect 1670 26228 1676 26240
rect 1631 26200 1676 26228
rect 1670 26188 1676 26200
rect 1728 26188 1734 26240
rect 1104 26138 36892 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 36892 26138
rect 1104 26064 36892 26086
rect 1104 25594 36892 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36892 25594
rect 1104 25520 36892 25542
rect 1104 25050 36892 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 36892 25050
rect 1104 24976 36892 24998
rect 25961 24803 26019 24809
rect 25961 24769 25973 24803
rect 26007 24800 26019 24803
rect 26602 24800 26608 24812
rect 26007 24772 26608 24800
rect 26007 24769 26019 24772
rect 25961 24763 26019 24769
rect 26602 24760 26608 24772
rect 26660 24760 26666 24812
rect 2406 24556 2412 24608
rect 2464 24596 2470 24608
rect 25869 24599 25927 24605
rect 25869 24596 25881 24599
rect 2464 24568 25881 24596
rect 2464 24556 2470 24568
rect 25869 24565 25881 24568
rect 25915 24565 25927 24599
rect 26602 24596 26608 24608
rect 26563 24568 26608 24596
rect 25869 24559 25927 24565
rect 26602 24556 26608 24568
rect 26660 24556 26666 24608
rect 1104 24506 36892 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36892 24506
rect 1104 24432 36892 24454
rect 35713 24191 35771 24197
rect 35713 24157 35725 24191
rect 35759 24188 35771 24191
rect 36354 24188 36360 24200
rect 35759 24160 36360 24188
rect 35759 24157 35771 24160
rect 35713 24151 35771 24157
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 1578 24080 1584 24132
rect 1636 24120 1642 24132
rect 1673 24123 1731 24129
rect 1673 24120 1685 24123
rect 1636 24092 1685 24120
rect 1636 24080 1642 24092
rect 1673 24089 1685 24092
rect 1719 24089 1731 24123
rect 1673 24083 1731 24089
rect 1857 24123 1915 24129
rect 1857 24089 1869 24123
rect 1903 24120 1915 24123
rect 7558 24120 7564 24132
rect 1903 24092 7564 24120
rect 1903 24089 1915 24092
rect 1857 24083 1915 24089
rect 7558 24080 7564 24092
rect 7616 24080 7622 24132
rect 36170 24052 36176 24064
rect 36131 24024 36176 24052
rect 36170 24012 36176 24024
rect 36228 24012 36234 24064
rect 1104 23962 36892 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 36892 23962
rect 1104 23888 36892 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 24394 23848 24400 23860
rect 24355 23820 24400 23848
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 23753 23715 23811 23721
rect 23753 23681 23765 23715
rect 23799 23712 23811 23715
rect 24412 23712 24440 23808
rect 23799 23684 24440 23712
rect 23799 23681 23811 23684
rect 23753 23675 23811 23681
rect 23845 23511 23903 23517
rect 23845 23477 23857 23511
rect 23891 23508 23903 23511
rect 24854 23508 24860 23520
rect 23891 23480 24860 23508
rect 23891 23477 23903 23480
rect 23845 23471 23903 23477
rect 24854 23468 24860 23480
rect 24912 23468 24918 23520
rect 1104 23418 36892 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36892 23418
rect 1104 23344 36892 23366
rect 19521 23239 19579 23245
rect 19521 23205 19533 23239
rect 19567 23236 19579 23239
rect 22002 23236 22008 23248
rect 19567 23208 22008 23236
rect 19567 23205 19579 23208
rect 19521 23199 19579 23205
rect 20180 23109 20208 23208
rect 22002 23196 22008 23208
rect 22060 23196 22066 23248
rect 21450 23168 21456 23180
rect 21411 23140 21456 23168
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 20165 23103 20223 23109
rect 20165 23069 20177 23103
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 17862 22992 17868 23044
rect 17920 23032 17926 23044
rect 20809 23035 20867 23041
rect 20809 23032 20821 23035
rect 17920 23004 20821 23032
rect 17920 22992 17926 23004
rect 20809 23001 20821 23004
rect 20855 23001 20867 23035
rect 20809 22995 20867 23001
rect 20990 22992 20996 23044
rect 21048 23032 21054 23044
rect 21361 23035 21419 23041
rect 21361 23032 21373 23035
rect 21048 23004 21373 23032
rect 21048 22992 21054 23004
rect 21361 23001 21373 23004
rect 21407 23001 21419 23035
rect 21361 22995 21419 23001
rect 20070 22964 20076 22976
rect 20031 22936 20076 22964
rect 20070 22924 20076 22936
rect 20128 22924 20134 22976
rect 1104 22874 36892 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 36892 22874
rect 1104 22800 36892 22822
rect 20990 22760 20996 22772
rect 20951 22732 20996 22760
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22624 1915 22627
rect 2130 22624 2136 22636
rect 1903 22596 2136 22624
rect 1903 22593 1915 22596
rect 1857 22587 1915 22593
rect 2130 22584 2136 22596
rect 2188 22584 2194 22636
rect 19797 22627 19855 22633
rect 19797 22593 19809 22627
rect 19843 22624 19855 22627
rect 20349 22627 20407 22633
rect 20349 22624 20361 22627
rect 19843 22596 20361 22624
rect 19843 22593 19855 22596
rect 19797 22587 19855 22593
rect 20349 22593 20361 22596
rect 20395 22624 20407 22627
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20395 22596 21097 22624
rect 20395 22593 20407 22596
rect 20349 22587 20407 22593
rect 21085 22593 21097 22596
rect 21131 22624 21143 22627
rect 21131 22596 22140 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 1670 22488 1676 22500
rect 1631 22460 1676 22488
rect 1670 22448 1676 22460
rect 1728 22448 1734 22500
rect 19705 22423 19763 22429
rect 19705 22389 19717 22423
rect 19751 22420 19763 22423
rect 19978 22420 19984 22432
rect 19751 22392 19984 22420
rect 19751 22389 19763 22392
rect 19705 22383 19763 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 22112 22429 22140 22596
rect 26602 22584 26608 22636
rect 26660 22624 26666 22636
rect 27341 22627 27399 22633
rect 27341 22624 27353 22627
rect 26660 22596 27353 22624
rect 26660 22584 26666 22596
rect 27341 22593 27353 22596
rect 27387 22624 27399 22627
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 27387 22596 27813 22624
rect 27387 22593 27399 22596
rect 27341 22587 27399 22593
rect 27801 22593 27813 22596
rect 27847 22593 27859 22627
rect 27801 22587 27859 22593
rect 32490 22584 32496 22636
rect 32548 22624 32554 22636
rect 36081 22627 36139 22633
rect 36081 22624 36093 22627
rect 32548 22596 36093 22624
rect 32548 22584 32554 22596
rect 36081 22593 36093 22596
rect 36127 22593 36139 22627
rect 36081 22587 36139 22593
rect 36262 22488 36268 22500
rect 36223 22460 36268 22488
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 22097 22423 22155 22429
rect 22097 22389 22109 22423
rect 22143 22420 22155 22423
rect 23842 22420 23848 22432
rect 22143 22392 23848 22420
rect 22143 22389 22155 22392
rect 22097 22383 22155 22389
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 26602 22380 26608 22432
rect 26660 22420 26666 22432
rect 27249 22423 27307 22429
rect 27249 22420 27261 22423
rect 26660 22392 27261 22420
rect 26660 22380 26666 22392
rect 27249 22389 27261 22392
rect 27295 22389 27307 22423
rect 27249 22383 27307 22389
rect 1104 22330 36892 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36892 22330
rect 1104 22256 36892 22278
rect 21450 22040 21456 22092
rect 21508 22080 21514 22092
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 21508 22052 22385 22080
rect 21508 22040 21514 22052
rect 22373 22049 22385 22052
rect 22419 22049 22431 22083
rect 22373 22043 22431 22049
rect 22465 21947 22523 21953
rect 22465 21913 22477 21947
rect 22511 21944 22523 21947
rect 22830 21944 22836 21956
rect 22511 21916 22836 21944
rect 22511 21913 22523 21916
rect 22465 21907 22523 21913
rect 22830 21904 22836 21916
rect 22888 21904 22894 21956
rect 23017 21947 23075 21953
rect 23017 21913 23029 21947
rect 23063 21944 23075 21947
rect 23566 21944 23572 21956
rect 23063 21916 23572 21944
rect 23063 21913 23075 21916
rect 23017 21907 23075 21913
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 15381 21879 15439 21885
rect 15381 21876 15393 21879
rect 15344 21848 15393 21876
rect 15344 21836 15350 21848
rect 15381 21845 15393 21848
rect 15427 21845 15439 21879
rect 15381 21839 15439 21845
rect 17586 21836 17592 21888
rect 17644 21876 17650 21888
rect 20441 21879 20499 21885
rect 20441 21876 20453 21879
rect 17644 21848 20453 21876
rect 17644 21836 17650 21848
rect 20441 21845 20453 21848
rect 20487 21876 20499 21879
rect 20714 21876 20720 21888
rect 20487 21848 20720 21876
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 1104 21786 36892 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 36892 21786
rect 1104 21712 36892 21734
rect 22830 21672 22836 21684
rect 22791 21644 22836 21672
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 15286 21604 15292 21616
rect 15247 21576 15292 21604
rect 15286 21564 15292 21576
rect 15344 21564 15350 21616
rect 15378 21564 15384 21616
rect 15436 21604 15442 21616
rect 15933 21607 15991 21613
rect 15436 21576 15481 21604
rect 15436 21564 15442 21576
rect 15933 21573 15945 21607
rect 15979 21604 15991 21607
rect 16666 21604 16672 21616
rect 15979 21576 16672 21604
rect 15979 21573 15991 21576
rect 15933 21567 15991 21573
rect 16666 21564 16672 21576
rect 16724 21604 16730 21616
rect 17862 21604 17868 21616
rect 16724 21576 17868 21604
rect 16724 21564 16730 21576
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 19978 21604 19984 21616
rect 19939 21576 19984 21604
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 20714 21604 20720 21616
rect 20675 21576 20720 21604
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21505 23627 21539
rect 23569 21499 23627 21505
rect 19426 21468 19432 21480
rect 19387 21440 19432 21468
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21468 20131 21471
rect 21910 21468 21916 21480
rect 20119 21440 21916 21468
rect 20119 21437 20131 21440
rect 20073 21431 20131 21437
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 22281 21403 22339 21409
rect 22281 21369 22293 21403
rect 22327 21400 22339 21403
rect 22940 21400 22968 21499
rect 23584 21400 23612 21499
rect 23750 21400 23756 21412
rect 22327 21372 23756 21400
rect 22327 21369 22339 21372
rect 22281 21363 22339 21369
rect 23750 21360 23756 21372
rect 23808 21400 23814 21412
rect 24029 21403 24087 21409
rect 24029 21400 24041 21403
rect 23808 21372 24041 21400
rect 23808 21360 23814 21372
rect 24029 21369 24041 21372
rect 24075 21369 24087 21403
rect 24029 21363 24087 21369
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 20806 21332 20812 21344
rect 20767 21304 20812 21332
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 23474 21332 23480 21344
rect 23435 21304 23480 21332
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 25133 21335 25191 21341
rect 25133 21301 25145 21335
rect 25179 21332 25191 21335
rect 25314 21332 25320 21344
rect 25179 21304 25320 21332
rect 25179 21301 25191 21304
rect 25133 21295 25191 21301
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 1104 21242 36892 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36892 21242
rect 1104 21168 36892 21190
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 34238 21128 34244 21140
rect 20864 21100 34244 21128
rect 20864 21088 20870 21100
rect 34238 21088 34244 21100
rect 34296 21088 34302 21140
rect 1578 20924 1584 20936
rect 1539 20896 1584 20924
rect 1578 20884 1584 20896
rect 1636 20884 1642 20936
rect 1854 20924 1860 20936
rect 1815 20896 1860 20924
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 17586 20924 17592 20936
rect 17547 20896 17592 20924
rect 17586 20884 17592 20896
rect 17644 20924 17650 20936
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 17644 20896 18061 20924
rect 17644 20884 17650 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 22278 20884 22284 20936
rect 22336 20924 22342 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22336 20896 22477 20924
rect 22336 20884 22342 20896
rect 22465 20893 22477 20896
rect 22511 20924 22523 20927
rect 23109 20927 23167 20933
rect 23109 20924 23121 20927
rect 22511 20896 23121 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 23109 20893 23121 20896
rect 23155 20893 23167 20927
rect 24946 20924 24952 20936
rect 24907 20896 24952 20924
rect 23109 20887 23167 20893
rect 24946 20884 24952 20896
rect 25004 20924 25010 20936
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 25004 20896 25421 20924
rect 25004 20884 25010 20896
rect 25409 20893 25421 20896
rect 25455 20924 25467 20927
rect 29822 20924 29828 20936
rect 25455 20896 29828 20924
rect 25455 20893 25467 20896
rect 25409 20887 25467 20893
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 35894 20884 35900 20936
rect 35952 20924 35958 20936
rect 36081 20927 36139 20933
rect 36081 20924 36093 20927
rect 35952 20896 36093 20924
rect 35952 20884 35958 20896
rect 36081 20893 36093 20896
rect 36127 20893 36139 20927
rect 36081 20887 36139 20893
rect 20898 20856 20904 20868
rect 20859 20828 20904 20856
rect 20898 20816 20904 20828
rect 20956 20816 20962 20868
rect 20990 20816 20996 20868
rect 21048 20856 21054 20868
rect 21542 20856 21548 20868
rect 21048 20828 21093 20856
rect 21503 20828 21548 20856
rect 21048 20816 21054 20828
rect 21542 20816 21548 20828
rect 21600 20816 21606 20868
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 17276 20760 17509 20788
rect 17276 20748 17282 20760
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 17497 20751 17555 20757
rect 22557 20791 22615 20797
rect 22557 20757 22569 20791
rect 22603 20788 22615 20791
rect 22738 20788 22744 20800
rect 22603 20760 22744 20788
rect 22603 20757 22615 20760
rect 22557 20751 22615 20757
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 24857 20791 24915 20797
rect 24857 20757 24869 20791
rect 24903 20788 24915 20791
rect 25222 20788 25228 20800
rect 24903 20760 25228 20788
rect 24903 20757 24915 20760
rect 24857 20751 24915 20757
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 25866 20748 25872 20800
rect 25924 20788 25930 20800
rect 25961 20791 26019 20797
rect 25961 20788 25973 20791
rect 25924 20760 25973 20788
rect 25924 20748 25930 20760
rect 25961 20757 25973 20760
rect 26007 20757 26019 20791
rect 36262 20788 36268 20800
rect 36223 20760 36268 20788
rect 25961 20751 26019 20757
rect 36262 20748 36268 20760
rect 36320 20748 36326 20800
rect 1104 20698 36892 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 36892 20698
rect 1104 20624 36892 20646
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 14921 20587 14979 20593
rect 14921 20553 14933 20587
rect 14967 20584 14979 20587
rect 15378 20584 15384 20596
rect 14967 20556 15384 20584
rect 14967 20553 14979 20556
rect 14921 20547 14979 20553
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20956 20556 21097 20584
rect 20956 20544 20962 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 21910 20544 21916 20596
rect 21968 20584 21974 20596
rect 30009 20587 30067 20593
rect 21968 20556 22876 20584
rect 21968 20544 21974 20556
rect 16942 20476 16948 20528
rect 17000 20516 17006 20528
rect 18785 20519 18843 20525
rect 18785 20516 18797 20519
rect 17000 20488 18797 20516
rect 17000 20476 17006 20488
rect 18785 20485 18797 20488
rect 18831 20485 18843 20519
rect 18785 20479 18843 20485
rect 19610 20476 19616 20528
rect 19668 20516 19674 20528
rect 20073 20519 20131 20525
rect 20073 20516 20085 20519
rect 19668 20488 20085 20516
rect 19668 20476 19674 20488
rect 20073 20485 20085 20488
rect 20119 20485 20131 20519
rect 20073 20479 20131 20485
rect 20625 20519 20683 20525
rect 20625 20485 20637 20519
rect 20671 20516 20683 20519
rect 22370 20516 22376 20528
rect 20671 20488 22376 20516
rect 20671 20485 20683 20488
rect 20625 20479 20683 20485
rect 22370 20476 22376 20488
rect 22428 20476 22434 20528
rect 22738 20516 22744 20528
rect 22699 20488 22744 20516
rect 22738 20476 22744 20488
rect 22796 20476 22802 20528
rect 22848 20525 22876 20556
rect 30009 20553 30021 20587
rect 30055 20584 30067 20587
rect 36078 20584 36084 20596
rect 30055 20556 36084 20584
rect 30055 20553 30067 20556
rect 30009 20547 30067 20553
rect 36078 20544 36084 20556
rect 36136 20544 36142 20596
rect 22833 20519 22891 20525
rect 22833 20485 22845 20519
rect 22879 20516 22891 20519
rect 23382 20516 23388 20528
rect 22879 20488 23388 20516
rect 22879 20485 22891 20488
rect 22833 20479 22891 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 24673 20519 24731 20525
rect 24673 20485 24685 20519
rect 24719 20516 24731 20519
rect 26513 20519 26571 20525
rect 26513 20516 26525 20519
rect 24719 20488 26525 20516
rect 24719 20485 24731 20488
rect 24673 20479 24731 20485
rect 26513 20485 26525 20488
rect 26559 20516 26571 20519
rect 27430 20516 27436 20528
rect 26559 20488 27436 20516
rect 26559 20485 26571 20488
rect 26513 20479 26571 20485
rect 27430 20476 27436 20488
rect 27488 20476 27494 20528
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 14829 20451 14887 20457
rect 1811 20420 2544 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 2516 20253 2544 20420
rect 14829 20417 14841 20451
rect 14875 20448 14887 20451
rect 15194 20448 15200 20460
rect 14875 20420 15200 20448
rect 14875 20417 14887 20420
rect 14829 20411 14887 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 25225 20451 25283 20457
rect 25225 20417 25237 20451
rect 25271 20448 25283 20451
rect 25314 20448 25320 20460
rect 25271 20420 25320 20448
rect 25271 20417 25283 20420
rect 25225 20411 25283 20417
rect 25314 20408 25320 20420
rect 25372 20408 25378 20460
rect 25866 20448 25872 20460
rect 25827 20420 25872 20448
rect 25866 20408 25872 20420
rect 25924 20408 25930 20460
rect 29086 20408 29092 20460
rect 29144 20448 29150 20460
rect 29917 20451 29975 20457
rect 29917 20448 29929 20451
rect 29144 20420 29929 20448
rect 29144 20408 29150 20420
rect 29917 20417 29929 20420
rect 29963 20417 29975 20451
rect 29917 20411 29975 20417
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 19334 20380 19340 20392
rect 18739 20352 19340 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 19334 20340 19340 20352
rect 19392 20380 19398 20392
rect 19981 20383 20039 20389
rect 19981 20380 19993 20383
rect 19392 20352 19993 20380
rect 19392 20340 19398 20352
rect 19981 20349 19993 20352
rect 20027 20380 20039 20383
rect 20070 20380 20076 20392
rect 20027 20352 20076 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23385 20383 23443 20389
rect 23385 20380 23397 20383
rect 23348 20352 23397 20380
rect 23348 20340 23354 20352
rect 23385 20349 23397 20352
rect 23431 20349 23443 20383
rect 23385 20343 23443 20349
rect 19245 20315 19303 20321
rect 19245 20281 19257 20315
rect 19291 20312 19303 20315
rect 22186 20312 22192 20324
rect 19291 20284 22192 20312
rect 19291 20281 19303 20284
rect 19245 20275 19303 20281
rect 22186 20272 22192 20284
rect 22244 20312 22250 20324
rect 22281 20315 22339 20321
rect 22281 20312 22293 20315
rect 22244 20284 22293 20312
rect 22244 20272 22250 20284
rect 22281 20281 22293 20284
rect 22327 20281 22339 20315
rect 22281 20275 22339 20281
rect 25317 20315 25375 20321
rect 25317 20281 25329 20315
rect 25363 20312 25375 20315
rect 27154 20312 27160 20324
rect 25363 20284 27160 20312
rect 25363 20281 25375 20284
rect 25317 20275 25375 20281
rect 27154 20272 27160 20284
rect 27212 20272 27218 20324
rect 2501 20247 2559 20253
rect 2501 20213 2513 20247
rect 2547 20244 2559 20247
rect 2682 20244 2688 20256
rect 2547 20216 2688 20244
rect 2547 20213 2559 20216
rect 2501 20207 2559 20213
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 24581 20247 24639 20253
rect 24581 20244 24593 20247
rect 18564 20216 24593 20244
rect 18564 20204 18570 20216
rect 24581 20213 24593 20216
rect 24627 20213 24639 20247
rect 25958 20244 25964 20256
rect 25919 20216 25964 20244
rect 24581 20207 24639 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 1104 20154 36892 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36892 20154
rect 1104 20080 36892 20102
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 25866 20040 25872 20052
rect 20180 20012 25872 20040
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 20180 19845 20208 20012
rect 25866 20000 25872 20012
rect 25924 20000 25930 20052
rect 22278 19932 22284 19984
rect 22336 19972 22342 19984
rect 23937 19975 23995 19981
rect 23937 19972 23949 19975
rect 22336 19944 23949 19972
rect 22336 19932 22342 19944
rect 23937 19941 23949 19944
rect 23983 19941 23995 19975
rect 23937 19935 23995 19941
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19904 22247 19907
rect 25222 19904 25228 19916
rect 22235 19876 23704 19904
rect 25183 19876 25228 19904
rect 22235 19873 22247 19876
rect 22189 19867 22247 19873
rect 16117 19839 16175 19845
rect 16117 19836 16129 19839
rect 14700 19808 16129 19836
rect 14700 19796 14706 19808
rect 16117 19805 16129 19808
rect 16163 19836 16175 19839
rect 16577 19839 16635 19845
rect 16577 19836 16589 19839
rect 16163 19808 16589 19836
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 16577 19805 16589 19808
rect 16623 19836 16635 19839
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 16623 19808 19533 19836
rect 16623 19805 16635 19808
rect 16577 19799 16635 19805
rect 19521 19805 19533 19808
rect 19567 19836 19579 19839
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 19567 19808 20177 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20898 19836 20904 19848
rect 20811 19808 20904 19836
rect 20165 19799 20223 19805
rect 20898 19796 20904 19808
rect 20956 19836 20962 19848
rect 21361 19839 21419 19845
rect 21361 19836 21373 19839
rect 20956 19808 21373 19836
rect 20956 19796 20962 19808
rect 21361 19805 21373 19808
rect 21407 19805 21419 19839
rect 21361 19799 21419 19805
rect 22094 19796 22100 19848
rect 22152 19836 22158 19848
rect 22152 19808 22197 19836
rect 22152 19796 22158 19808
rect 17221 19771 17279 19777
rect 17221 19737 17233 19771
rect 17267 19768 17279 19771
rect 17954 19768 17960 19780
rect 17267 19740 17960 19768
rect 17267 19737 17279 19740
rect 17221 19731 17279 19737
rect 17954 19728 17960 19740
rect 18012 19728 18018 19780
rect 18601 19771 18659 19777
rect 18601 19737 18613 19771
rect 18647 19768 18659 19771
rect 18690 19768 18696 19780
rect 18647 19740 18696 19768
rect 18647 19737 18659 19740
rect 18601 19731 18659 19737
rect 18690 19728 18696 19740
rect 18748 19768 18754 19780
rect 22278 19768 22284 19780
rect 18748 19740 22284 19768
rect 18748 19728 18754 19740
rect 22278 19728 22284 19740
rect 22336 19728 22342 19780
rect 22741 19771 22799 19777
rect 22741 19737 22753 19771
rect 22787 19768 22799 19771
rect 22922 19768 22928 19780
rect 22787 19740 22928 19768
rect 22787 19737 22799 19740
rect 22741 19731 22799 19737
rect 22922 19728 22928 19740
rect 22980 19728 22986 19780
rect 23293 19771 23351 19777
rect 23293 19737 23305 19771
rect 23339 19737 23351 19771
rect 23293 19731 23351 19737
rect 2130 19660 2136 19712
rect 2188 19700 2194 19712
rect 2314 19700 2320 19712
rect 2188 19672 2320 19700
rect 2188 19660 2194 19672
rect 2314 19660 2320 19672
rect 2372 19660 2378 19712
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 16025 19703 16083 19709
rect 16025 19700 16037 19703
rect 15344 19672 16037 19700
rect 15344 19660 15350 19672
rect 16025 19669 16037 19672
rect 16071 19669 16083 19703
rect 17678 19700 17684 19712
rect 17639 19672 17684 19700
rect 16025 19663 16083 19669
rect 17678 19660 17684 19672
rect 17736 19660 17742 19712
rect 21450 19700 21456 19712
rect 21411 19672 21456 19700
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 23308 19700 23336 19731
rect 23382 19728 23388 19780
rect 23440 19768 23446 19780
rect 23676 19768 23704 19876
rect 25222 19864 25228 19876
rect 25280 19904 25286 19916
rect 25869 19907 25927 19913
rect 25869 19904 25881 19907
rect 25280 19876 25881 19904
rect 25280 19864 25286 19876
rect 25869 19873 25881 19876
rect 25915 19873 25927 19907
rect 25869 19867 25927 19873
rect 23440 19740 23485 19768
rect 23676 19740 24532 19768
rect 23440 19728 23446 19740
rect 23474 19700 23480 19712
rect 23308 19672 23480 19700
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 24504 19700 24532 19740
rect 24578 19728 24584 19780
rect 24636 19768 24642 19780
rect 25133 19771 25191 19777
rect 24636 19740 24681 19768
rect 24636 19728 24642 19740
rect 25133 19737 25145 19771
rect 25179 19737 25191 19771
rect 25133 19731 25191 19737
rect 25148 19700 25176 19731
rect 25958 19728 25964 19780
rect 26016 19768 26022 19780
rect 26513 19771 26571 19777
rect 26016 19740 26061 19768
rect 26016 19728 26022 19740
rect 26513 19737 26525 19771
rect 26559 19737 26571 19771
rect 27062 19768 27068 19780
rect 27023 19740 27068 19768
rect 26513 19731 26571 19737
rect 24504 19672 25176 19700
rect 26528 19700 26556 19731
rect 27062 19728 27068 19740
rect 27120 19728 27126 19780
rect 27154 19728 27160 19780
rect 27212 19768 27218 19780
rect 27709 19771 27767 19777
rect 27709 19768 27721 19771
rect 27212 19740 27257 19768
rect 27632 19740 27721 19768
rect 27212 19728 27218 19740
rect 27632 19712 27660 19740
rect 27709 19737 27721 19740
rect 27755 19737 27767 19771
rect 27709 19731 27767 19737
rect 27614 19700 27620 19712
rect 26528 19672 27620 19700
rect 27614 19660 27620 19672
rect 27672 19660 27678 19712
rect 1104 19610 36892 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 36892 19610
rect 1104 19536 36892 19558
rect 15105 19499 15163 19505
rect 15105 19465 15117 19499
rect 15151 19496 15163 19499
rect 15470 19496 15476 19508
rect 15151 19468 15476 19496
rect 15151 19465 15163 19468
rect 15105 19459 15163 19465
rect 15470 19456 15476 19468
rect 15528 19496 15534 19508
rect 19337 19499 19395 19505
rect 15528 19468 17448 19496
rect 15528 19456 15534 19468
rect 17310 19428 17316 19440
rect 17271 19400 17316 19428
rect 17310 19388 17316 19400
rect 17368 19388 17374 19440
rect 17420 19428 17448 19468
rect 19337 19465 19349 19499
rect 19383 19496 19395 19499
rect 20990 19496 20996 19508
rect 19383 19468 20996 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 25777 19499 25835 19505
rect 22143 19468 24992 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 20898 19428 20904 19440
rect 17420 19400 20904 19428
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 21450 19388 21456 19440
rect 21508 19428 21514 19440
rect 24964 19437 24992 19468
rect 25777 19465 25789 19499
rect 25823 19465 25835 19499
rect 25777 19459 25835 19465
rect 23385 19431 23443 19437
rect 23385 19428 23397 19431
rect 21508 19400 23397 19428
rect 21508 19388 21514 19400
rect 23385 19397 23397 19400
rect 23431 19397 23443 19431
rect 23385 19391 23443 19397
rect 24949 19431 25007 19437
rect 24949 19397 24961 19431
rect 24995 19397 25007 19431
rect 24949 19391 25007 19397
rect 25041 19431 25099 19437
rect 25041 19397 25053 19431
rect 25087 19428 25099 19431
rect 25498 19428 25504 19440
rect 25087 19400 25504 19428
rect 25087 19397 25099 19400
rect 25041 19391 25099 19397
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 25792 19428 25820 19459
rect 27062 19456 27068 19508
rect 27120 19496 27126 19508
rect 27157 19499 27215 19505
rect 27157 19496 27169 19499
rect 27120 19468 27169 19496
rect 27120 19456 27126 19468
rect 27157 19465 27169 19468
rect 27203 19465 27215 19499
rect 32490 19496 32496 19508
rect 32451 19468 32496 19496
rect 27157 19459 27215 19465
rect 32490 19456 32496 19468
rect 32548 19456 32554 19508
rect 35894 19428 35900 19440
rect 25792 19400 35900 19428
rect 35894 19388 35900 19400
rect 35952 19388 35958 19440
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1636 19332 1685 19360
rect 1636 19320 1642 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 16022 19360 16028 19372
rect 15703 19332 16028 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 16022 19320 16028 19332
rect 16080 19360 16086 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 16080 19332 16129 19360
rect 16080 19320 16086 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16209 19363 16267 19369
rect 16209 19329 16221 19363
rect 16255 19360 16267 19363
rect 17034 19360 17040 19372
rect 16255 19332 17040 19360
rect 16255 19329 16267 19332
rect 16209 19323 16267 19329
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 20622 19360 20628 19372
rect 19291 19332 20628 19360
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21376 19332 22017 19360
rect 17218 19292 17224 19304
rect 17179 19264 17224 19292
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 19426 19292 19432 19304
rect 17911 19264 19432 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 1857 19227 1915 19233
rect 1857 19193 1869 19227
rect 1903 19224 1915 19227
rect 6822 19224 6828 19236
rect 1903 19196 6828 19224
rect 1903 19193 1915 19196
rect 1857 19187 1915 19193
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 15378 19184 15384 19236
rect 15436 19224 15442 19236
rect 17880 19224 17908 19255
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21376 19301 21404 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 25593 19363 25651 19369
rect 25593 19329 25605 19363
rect 25639 19329 25651 19363
rect 25593 19323 25651 19329
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19329 26479 19363
rect 32306 19360 32312 19372
rect 26421 19323 26479 19329
rect 27586 19332 27844 19360
rect 32267 19332 32312 19360
rect 21361 19295 21419 19301
rect 21361 19292 21373 19295
rect 21140 19264 21373 19292
rect 21140 19252 21146 19264
rect 21361 19261 21373 19264
rect 21407 19261 21419 19295
rect 21361 19255 21419 19261
rect 21634 19252 21640 19304
rect 21692 19292 21698 19304
rect 22094 19292 22100 19304
rect 21692 19264 22100 19292
rect 21692 19252 21698 19264
rect 22094 19252 22100 19264
rect 22152 19292 22158 19304
rect 22649 19295 22707 19301
rect 22649 19292 22661 19295
rect 22152 19264 22661 19292
rect 22152 19252 22158 19264
rect 22649 19261 22661 19264
rect 22695 19261 22707 19295
rect 23290 19292 23296 19304
rect 23251 19264 23296 19292
rect 22649 19255 22707 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 23566 19292 23572 19304
rect 23527 19264 23572 19292
rect 23566 19252 23572 19264
rect 23624 19252 23630 19304
rect 24397 19295 24455 19301
rect 24397 19292 24409 19295
rect 23768 19264 24409 19292
rect 15436 19196 17908 19224
rect 15436 19184 15442 19196
rect 18782 19184 18788 19236
rect 18840 19224 18846 19236
rect 21542 19224 21548 19236
rect 18840 19196 21548 19224
rect 18840 19184 18846 19196
rect 21542 19184 21548 19196
rect 21600 19224 21606 19236
rect 23768 19224 23796 19264
rect 24397 19261 24409 19264
rect 24443 19292 24455 19295
rect 24578 19292 24584 19304
rect 24443 19264 24584 19292
rect 24443 19261 24455 19264
rect 24397 19255 24455 19261
rect 24578 19252 24584 19264
rect 24636 19252 24642 19304
rect 25608 19236 25636 19323
rect 26428 19292 26456 19323
rect 27062 19292 27068 19304
rect 26428 19264 27068 19292
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 25590 19224 25596 19236
rect 21600 19196 23796 19224
rect 25503 19196 25596 19224
rect 21600 19184 21606 19196
rect 25590 19184 25596 19196
rect 25648 19224 25654 19236
rect 27586 19224 27614 19332
rect 27816 19301 27844 19332
rect 32306 19320 32312 19332
rect 32364 19360 32370 19372
rect 32953 19363 33011 19369
rect 32953 19360 32965 19363
rect 32364 19332 32965 19360
rect 32364 19320 32370 19332
rect 32953 19329 32965 19332
rect 32999 19329 33011 19363
rect 36078 19360 36084 19372
rect 36039 19332 36084 19360
rect 32953 19323 33011 19329
rect 36078 19320 36084 19332
rect 36136 19320 36142 19372
rect 27801 19295 27859 19301
rect 27801 19261 27813 19295
rect 27847 19292 27859 19295
rect 27847 19264 27881 19292
rect 27847 19261 27859 19264
rect 27801 19255 27859 19261
rect 25648 19196 27614 19224
rect 25648 19184 25654 19196
rect 14550 19156 14556 19168
rect 14511 19128 14556 19156
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 17954 19156 17960 19168
rect 16172 19128 17960 19156
rect 16172 19116 16178 19128
rect 17954 19116 17960 19128
rect 18012 19156 18018 19168
rect 18693 19159 18751 19165
rect 18693 19156 18705 19159
rect 18012 19128 18705 19156
rect 18012 19116 18018 19128
rect 18693 19125 18705 19128
rect 18739 19156 18751 19159
rect 19150 19156 19156 19168
rect 18739 19128 19156 19156
rect 18739 19125 18751 19128
rect 18693 19119 18751 19125
rect 19150 19116 19156 19128
rect 19208 19116 19214 19168
rect 19981 19159 20039 19165
rect 19981 19125 19993 19159
rect 20027 19156 20039 19159
rect 20070 19156 20076 19168
rect 20027 19128 20076 19156
rect 20027 19125 20039 19128
rect 19981 19119 20039 19125
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 20901 19159 20959 19165
rect 20901 19125 20913 19159
rect 20947 19156 20959 19159
rect 21266 19156 21272 19168
rect 20947 19128 21272 19156
rect 20947 19125 20959 19128
rect 20901 19119 20959 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21358 19116 21364 19168
rect 21416 19156 21422 19168
rect 22554 19156 22560 19168
rect 21416 19128 22560 19156
rect 21416 19116 21422 19128
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 25866 19116 25872 19168
rect 25924 19156 25930 19168
rect 26329 19159 26387 19165
rect 26329 19156 26341 19159
rect 25924 19128 26341 19156
rect 25924 19116 25930 19128
rect 26329 19125 26341 19128
rect 26375 19125 26387 19159
rect 36262 19156 36268 19168
rect 36223 19128 36268 19156
rect 26329 19119 26387 19125
rect 36262 19116 36268 19128
rect 36320 19116 36326 19168
rect 1104 19066 36892 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36892 19066
rect 1104 18992 36892 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 13725 18955 13783 18961
rect 13725 18921 13737 18955
rect 13771 18952 13783 18955
rect 14274 18952 14280 18964
rect 13771 18924 14280 18952
rect 13771 18921 13783 18924
rect 13725 18915 13783 18921
rect 14274 18912 14280 18924
rect 14332 18952 14338 18964
rect 15470 18952 15476 18964
rect 14332 18924 15476 18952
rect 14332 18912 14338 18924
rect 15470 18912 15476 18924
rect 15528 18952 15534 18964
rect 15838 18952 15844 18964
rect 15528 18924 15844 18952
rect 15528 18912 15534 18924
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 16117 18955 16175 18961
rect 16117 18921 16129 18955
rect 16163 18952 16175 18955
rect 17310 18952 17316 18964
rect 16163 18924 17316 18952
rect 16163 18921 16175 18924
rect 16117 18915 16175 18921
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 25590 18952 25596 18964
rect 20864 18924 25596 18952
rect 20864 18912 20870 18924
rect 25590 18912 25596 18924
rect 25648 18912 25654 18964
rect 25958 18912 25964 18964
rect 26016 18912 26022 18964
rect 27062 18912 27068 18964
rect 27120 18952 27126 18964
rect 27801 18955 27859 18961
rect 27801 18952 27813 18955
rect 27120 18924 27813 18952
rect 27120 18912 27126 18924
rect 27801 18921 27813 18924
rect 27847 18921 27859 18955
rect 27801 18915 27859 18921
rect 17972 18856 20392 18884
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14608 18720 14657 18748
rect 14608 18708 14614 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 14660 18680 14688 18711
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 15252 18720 15301 18748
rect 15252 18708 15258 18720
rect 15289 18717 15301 18720
rect 15335 18748 15347 18751
rect 15930 18748 15936 18760
rect 15335 18720 15936 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16114 18748 16120 18760
rect 16071 18720 16120 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18748 16727 18751
rect 17972 18748 18000 18856
rect 18782 18816 18788 18828
rect 18743 18788 18788 18816
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 20364 18757 20392 18856
rect 20530 18844 20536 18896
rect 20588 18884 20594 18896
rect 23201 18887 23259 18893
rect 23201 18884 23213 18887
rect 20588 18856 23213 18884
rect 20588 18844 20594 18856
rect 23201 18853 23213 18856
rect 23247 18884 23259 18887
rect 25976 18884 26004 18912
rect 23247 18856 26004 18884
rect 23247 18853 23259 18856
rect 23201 18847 23259 18853
rect 21358 18816 21364 18828
rect 21008 18788 21364 18816
rect 21008 18760 21036 18788
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 22554 18776 22560 18828
rect 22612 18816 22618 18828
rect 25700 18825 25728 18856
rect 25685 18819 25743 18825
rect 22612 18788 24624 18816
rect 22612 18776 22618 18788
rect 16715 18720 18000 18748
rect 20349 18751 20407 18757
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 20349 18717 20361 18751
rect 20395 18748 20407 18751
rect 20990 18748 20996 18760
rect 20395 18720 20996 18748
rect 20395 18717 20407 18720
rect 20349 18711 20407 18717
rect 20990 18708 20996 18720
rect 21048 18708 21054 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 21818 18748 21824 18760
rect 21131 18720 21824 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 17773 18683 17831 18689
rect 14660 18652 16896 18680
rect 14734 18612 14740 18624
rect 14695 18584 14740 18612
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 15381 18615 15439 18621
rect 15381 18581 15393 18615
rect 15427 18612 15439 18615
rect 15470 18612 15476 18624
rect 15427 18584 15476 18612
rect 15427 18581 15439 18584
rect 15381 18575 15439 18581
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 16758 18612 16764 18624
rect 16719 18584 16764 18612
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 16868 18612 16896 18652
rect 17773 18649 17785 18683
rect 17819 18680 17831 18683
rect 17954 18680 17960 18692
rect 17819 18652 17960 18680
rect 17819 18649 17831 18652
rect 17773 18643 17831 18649
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18693 18683 18751 18689
rect 18693 18649 18705 18683
rect 18739 18680 18751 18683
rect 19978 18680 19984 18692
rect 18739 18652 19984 18680
rect 18739 18649 18751 18652
rect 18693 18643 18751 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 21100 18680 21128 18711
rect 21818 18708 21824 18720
rect 21876 18708 21882 18760
rect 22278 18708 22284 18760
rect 22336 18748 22342 18760
rect 24596 18757 24624 18788
rect 25685 18785 25697 18819
rect 25731 18785 25743 18819
rect 25685 18779 25743 18785
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 26602 18816 26608 18828
rect 26007 18788 26608 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 22373 18751 22431 18757
rect 22373 18748 22385 18751
rect 22336 18720 22385 18748
rect 22336 18708 22342 18720
rect 22373 18717 22385 18720
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 26694 18748 26700 18760
rect 26655 18720 26700 18748
rect 24581 18711 24639 18717
rect 26694 18708 26700 18720
rect 26752 18708 26758 18760
rect 27154 18748 27160 18760
rect 27115 18720 27160 18748
rect 27154 18708 27160 18720
rect 27212 18748 27218 18760
rect 28353 18751 28411 18757
rect 28353 18748 28365 18751
rect 27212 18720 28365 18748
rect 27212 18708 27218 18720
rect 28353 18717 28365 18720
rect 28399 18717 28411 18751
rect 28353 18711 28411 18717
rect 20088 18652 21128 18680
rect 23661 18683 23719 18689
rect 18322 18612 18328 18624
rect 16868 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19521 18615 19579 18621
rect 19521 18612 19533 18615
rect 18656 18584 19533 18612
rect 18656 18572 18662 18584
rect 19521 18581 19533 18584
rect 19567 18612 19579 18615
rect 20088 18612 20116 18652
rect 23661 18649 23673 18683
rect 23707 18649 23719 18683
rect 23661 18643 23719 18649
rect 23753 18683 23811 18689
rect 23753 18649 23765 18683
rect 23799 18680 23811 18683
rect 24026 18680 24032 18692
rect 23799 18652 24032 18680
rect 23799 18649 23811 18652
rect 23753 18643 23811 18649
rect 20254 18612 20260 18624
rect 19567 18584 20116 18612
rect 20215 18584 20260 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 21450 18572 21456 18624
rect 21508 18612 21514 18624
rect 21729 18615 21787 18621
rect 21729 18612 21741 18615
rect 21508 18584 21741 18612
rect 21508 18572 21514 18584
rect 21729 18581 21741 18584
rect 21775 18581 21787 18615
rect 21729 18575 21787 18581
rect 22465 18615 22523 18621
rect 22465 18581 22477 18615
rect 22511 18612 22523 18615
rect 22738 18612 22744 18624
rect 22511 18584 22744 18612
rect 22511 18581 22523 18584
rect 22465 18575 22523 18581
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 23676 18612 23704 18643
rect 24026 18640 24032 18652
rect 24084 18640 24090 18692
rect 24854 18680 24860 18692
rect 24596 18652 24860 18680
rect 24596 18612 24624 18652
rect 24854 18640 24860 18652
rect 24912 18640 24918 18692
rect 25866 18680 25872 18692
rect 25827 18652 25872 18680
rect 25866 18640 25872 18652
rect 25924 18640 25930 18692
rect 23676 18584 24624 18612
rect 24673 18615 24731 18621
rect 24673 18581 24685 18615
rect 24719 18612 24731 18615
rect 24946 18612 24952 18624
rect 24719 18584 24952 18612
rect 24719 18581 24731 18584
rect 24673 18575 24731 18581
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 26605 18615 26663 18621
rect 26605 18612 26617 18615
rect 25648 18584 26617 18612
rect 25648 18572 25654 18584
rect 26605 18581 26617 18584
rect 26651 18581 26663 18615
rect 26605 18575 26663 18581
rect 27249 18615 27307 18621
rect 27249 18581 27261 18615
rect 27295 18612 27307 18615
rect 27706 18612 27712 18624
rect 27295 18584 27712 18612
rect 27295 18581 27307 18584
rect 27249 18575 27307 18581
rect 27706 18572 27712 18584
rect 27764 18572 27770 18624
rect 1104 18522 36892 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 36892 18522
rect 1104 18448 36892 18470
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15010 18408 15016 18420
rect 14516 18380 15016 18408
rect 14516 18368 14522 18380
rect 15010 18368 15016 18380
rect 15068 18408 15074 18420
rect 18782 18408 18788 18420
rect 15068 18380 15976 18408
rect 15068 18368 15074 18380
rect 14090 18340 14096 18352
rect 14051 18312 14096 18340
rect 14090 18300 14096 18312
rect 14148 18300 14154 18352
rect 14185 18343 14243 18349
rect 14185 18309 14197 18343
rect 14231 18340 14243 18343
rect 15286 18340 15292 18352
rect 14231 18312 15292 18340
rect 14231 18309 14243 18312
rect 14185 18303 14243 18309
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 15381 18343 15439 18349
rect 15381 18309 15393 18343
rect 15427 18340 15439 18343
rect 15654 18340 15660 18352
rect 15427 18312 15660 18340
rect 15427 18309 15439 18312
rect 15381 18303 15439 18309
rect 15654 18300 15660 18312
rect 15712 18300 15718 18352
rect 15948 18349 15976 18380
rect 16040 18380 18788 18408
rect 15933 18343 15991 18349
rect 15933 18309 15945 18343
rect 15979 18309 15991 18343
rect 15933 18303 15991 18309
rect 12710 18272 12716 18284
rect 12623 18244 12716 18272
rect 12710 18232 12716 18244
rect 12768 18272 12774 18284
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 12768 18244 13185 18272
rect 12768 18232 12774 18244
rect 13173 18241 13185 18244
rect 13219 18272 13231 18275
rect 13219 18244 13952 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13262 18068 13268 18080
rect 13223 18040 13268 18068
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 13924 18068 13952 18244
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 15102 18204 15108 18216
rect 14783 18176 15108 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18204 15347 18207
rect 15378 18204 15384 18216
rect 15335 18176 15384 18204
rect 15335 18173 15347 18176
rect 15289 18167 15347 18173
rect 15378 18164 15384 18176
rect 15436 18164 15442 18216
rect 16040 18136 16068 18380
rect 18782 18368 18788 18380
rect 18840 18408 18846 18420
rect 21634 18408 21640 18420
rect 18840 18380 21640 18408
rect 18840 18368 18846 18380
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 24026 18408 24032 18420
rect 23987 18380 24032 18408
rect 24026 18368 24032 18380
rect 24084 18368 24090 18420
rect 26694 18368 26700 18420
rect 26752 18408 26758 18420
rect 27801 18411 27859 18417
rect 27801 18408 27813 18411
rect 26752 18380 27813 18408
rect 26752 18368 26758 18380
rect 27801 18377 27813 18380
rect 27847 18377 27859 18411
rect 27801 18371 27859 18377
rect 28810 18368 28816 18420
rect 28868 18408 28874 18420
rect 32306 18408 32312 18420
rect 28868 18380 32312 18408
rect 28868 18368 28874 18380
rect 32306 18368 32312 18380
rect 32364 18368 32370 18420
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 17773 18343 17831 18349
rect 17773 18340 17785 18343
rect 16816 18312 17785 18340
rect 16816 18300 16822 18312
rect 17773 18309 17785 18312
rect 17819 18309 17831 18343
rect 17773 18303 17831 18309
rect 18325 18343 18383 18349
rect 18325 18309 18337 18343
rect 18371 18340 18383 18343
rect 19426 18340 19432 18352
rect 18371 18312 19432 18340
rect 18371 18309 18383 18312
rect 18325 18303 18383 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 20254 18340 20260 18352
rect 20215 18312 20260 18340
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 20809 18343 20867 18349
rect 20809 18309 20821 18343
rect 20855 18340 20867 18343
rect 22186 18340 22192 18352
rect 20855 18312 22192 18340
rect 20855 18309 20867 18312
rect 20809 18303 20867 18309
rect 22186 18300 22192 18312
rect 22244 18340 22250 18352
rect 22557 18343 22615 18349
rect 22557 18340 22569 18343
rect 22244 18312 22569 18340
rect 22244 18300 22250 18312
rect 22557 18309 22569 18312
rect 22603 18309 22615 18343
rect 22557 18303 22615 18309
rect 22649 18343 22707 18349
rect 22649 18309 22661 18343
rect 22695 18340 22707 18343
rect 23569 18343 23627 18349
rect 22695 18312 23520 18340
rect 22695 18309 22707 18312
rect 22649 18303 22707 18309
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16448 18244 16957 18272
rect 16448 18232 16454 18244
rect 16945 18241 16957 18244
rect 16991 18241 17003 18275
rect 16945 18235 17003 18241
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 18969 18275 19027 18281
rect 18969 18272 18981 18275
rect 18656 18244 18981 18272
rect 18656 18232 18662 18244
rect 18969 18241 18981 18244
rect 19015 18241 19027 18275
rect 21266 18272 21272 18284
rect 21227 18244 21272 18272
rect 18969 18235 19027 18241
rect 21266 18232 21272 18244
rect 21324 18272 21330 18284
rect 23492 18272 23520 18312
rect 23569 18309 23581 18343
rect 23615 18340 23627 18343
rect 23658 18340 23664 18352
rect 23615 18312 23664 18340
rect 23615 18309 23627 18312
rect 23569 18303 23627 18309
rect 23658 18300 23664 18312
rect 23716 18340 23722 18352
rect 24118 18340 24124 18352
rect 23716 18312 24124 18340
rect 23716 18300 23722 18312
rect 24118 18300 24124 18312
rect 24176 18300 24182 18352
rect 25590 18340 25596 18352
rect 25551 18312 25596 18340
rect 25590 18300 25596 18312
rect 25648 18300 25654 18352
rect 24762 18272 24768 18284
rect 21324 18244 22094 18272
rect 23492 18244 24768 18272
rect 21324 18232 21330 18244
rect 17218 18164 17224 18216
rect 17276 18204 17282 18216
rect 17681 18207 17739 18213
rect 17681 18204 17693 18207
rect 17276 18176 17693 18204
rect 17276 18164 17282 18176
rect 17681 18173 17693 18176
rect 17727 18173 17739 18207
rect 20162 18204 20168 18216
rect 20123 18176 20168 18204
rect 17681 18167 17739 18173
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 22066 18204 22094 18244
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27338 18232 27344 18244
rect 27396 18272 27402 18284
rect 28353 18275 28411 18281
rect 28353 18272 28365 18275
rect 27396 18244 28365 18272
rect 27396 18232 27402 18244
rect 28353 18241 28365 18244
rect 28399 18241 28411 18275
rect 28353 18235 28411 18241
rect 23750 18204 23756 18216
rect 22066 18176 23756 18204
rect 23750 18164 23756 18176
rect 23808 18204 23814 18216
rect 24118 18204 24124 18216
rect 23808 18176 24124 18204
rect 23808 18164 23814 18176
rect 24118 18164 24124 18176
rect 24176 18164 24182 18216
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24673 18207 24731 18213
rect 24673 18204 24685 18207
rect 24268 18176 24685 18204
rect 24268 18164 24274 18176
rect 24673 18173 24685 18176
rect 24719 18173 24731 18207
rect 25498 18204 25504 18216
rect 25459 18176 25504 18204
rect 24673 18167 24731 18173
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 26145 18207 26203 18213
rect 26145 18173 26157 18207
rect 26191 18204 26203 18207
rect 27614 18204 27620 18216
rect 26191 18176 27620 18204
rect 26191 18173 26203 18176
rect 26145 18167 26203 18173
rect 27614 18164 27620 18176
rect 27672 18164 27678 18216
rect 15304 18108 16068 18136
rect 17037 18139 17095 18145
rect 15304 18068 15332 18108
rect 17037 18105 17049 18139
rect 17083 18136 17095 18139
rect 18138 18136 18144 18148
rect 17083 18108 18144 18136
rect 17083 18105 17095 18108
rect 17037 18099 17095 18105
rect 18138 18096 18144 18108
rect 18196 18096 18202 18148
rect 18322 18096 18328 18148
rect 18380 18136 18386 18148
rect 25314 18136 25320 18148
rect 18380 18108 25320 18136
rect 18380 18096 18386 18108
rect 25314 18096 25320 18108
rect 25372 18096 25378 18148
rect 13924 18040 15332 18068
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 16482 18068 16488 18080
rect 15896 18040 16488 18068
rect 15896 18028 15902 18040
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 18877 18071 18935 18077
rect 18877 18068 18889 18071
rect 18104 18040 18889 18068
rect 18104 18028 18110 18040
rect 18877 18037 18889 18040
rect 18923 18037 18935 18071
rect 18877 18031 18935 18037
rect 19613 18071 19671 18077
rect 19613 18037 19625 18071
rect 19659 18068 19671 18071
rect 20806 18068 20812 18080
rect 19659 18040 20812 18068
rect 19659 18037 19671 18040
rect 19613 18031 19671 18037
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 22462 18068 22468 18080
rect 21407 18040 22468 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 22646 18028 22652 18080
rect 22704 18068 22710 18080
rect 27062 18068 27068 18080
rect 22704 18040 27068 18068
rect 22704 18028 22710 18040
rect 27062 18028 27068 18040
rect 27120 18028 27126 18080
rect 27246 18068 27252 18080
rect 27207 18040 27252 18068
rect 27246 18028 27252 18040
rect 27304 18028 27310 18080
rect 28810 18028 28816 18080
rect 28868 18068 28874 18080
rect 28997 18071 29055 18077
rect 28997 18068 29009 18071
rect 28868 18040 29009 18068
rect 28868 18028 28874 18040
rect 28997 18037 29009 18040
rect 29043 18037 29055 18071
rect 28997 18031 29055 18037
rect 1104 17978 36892 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36892 17978
rect 1104 17904 36892 17926
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 6822 17864 6828 17876
rect 6420 17836 6828 17864
rect 6420 17824 6426 17836
rect 6822 17824 6828 17836
rect 6880 17864 6886 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 6880 17836 10701 17864
rect 6880 17824 6886 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 10704 17660 10732 17827
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13170 17864 13176 17876
rect 12492 17836 13176 17864
rect 12492 17824 12498 17836
rect 13170 17824 13176 17836
rect 13228 17864 13234 17876
rect 13633 17867 13691 17873
rect 13228 17836 13584 17864
rect 13228 17824 13234 17836
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 10704 17632 11253 17660
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13446 17660 13452 17672
rect 13127 17632 13452 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 13556 17669 13584 17836
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 20162 17864 20168 17876
rect 13679 17836 20168 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 28350 17864 28356 17876
rect 27540 17836 28356 17864
rect 15013 17799 15071 17805
rect 15013 17765 15025 17799
rect 15059 17796 15071 17799
rect 15378 17796 15384 17808
rect 15059 17768 15384 17796
rect 15059 17765 15071 17768
rect 15013 17759 15071 17765
rect 15378 17756 15384 17768
rect 15436 17756 15442 17808
rect 16114 17756 16120 17808
rect 16172 17796 16178 17808
rect 21082 17796 21088 17808
rect 16172 17768 21088 17796
rect 16172 17756 16178 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 22830 17756 22836 17808
rect 22888 17796 22894 17808
rect 26145 17799 26203 17805
rect 26145 17796 26157 17799
rect 22888 17768 26157 17796
rect 22888 17756 22894 17768
rect 26145 17765 26157 17768
rect 26191 17796 26203 17799
rect 27338 17796 27344 17808
rect 26191 17768 27344 17796
rect 26191 17765 26203 17768
rect 26145 17759 26203 17765
rect 27338 17756 27344 17768
rect 27396 17756 27402 17808
rect 15286 17728 15292 17740
rect 14936 17700 15292 17728
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17629 13599 17663
rect 14274 17660 14280 17672
rect 14235 17632 14280 17660
rect 13541 17623 13599 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 11333 17595 11391 17601
rect 11333 17561 11345 17595
rect 11379 17592 11391 17595
rect 14936 17592 14964 17700
rect 15286 17688 15292 17700
rect 15344 17728 15350 17740
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15344 17700 16221 17728
rect 15344 17688 15350 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 16209 17691 16267 17697
rect 17218 17688 17224 17740
rect 17276 17728 17282 17740
rect 17405 17731 17463 17737
rect 17405 17728 17417 17731
rect 17276 17700 17417 17728
rect 17276 17688 17282 17700
rect 17405 17697 17417 17700
rect 17451 17697 17463 17731
rect 17405 17691 17463 17697
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 19392 17700 19533 17728
rect 19392 17688 19398 17700
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 20162 17688 20168 17740
rect 20220 17728 20226 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 20220 17700 21373 17728
rect 20220 17688 20226 17700
rect 21361 17697 21373 17700
rect 21407 17697 21419 17731
rect 21361 17691 21419 17697
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22370 17728 22376 17740
rect 22051 17700 22376 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 22922 17728 22928 17740
rect 22883 17700 22928 17728
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 25774 17728 25780 17740
rect 23983 17700 25780 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 27433 17731 27491 17737
rect 27433 17728 27445 17731
rect 26252 17700 27445 17728
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 19150 17660 19156 17672
rect 18739 17632 19156 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 20806 17660 20812 17672
rect 20767 17632 20812 17660
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 15470 17592 15476 17604
rect 11379 17564 14964 17592
rect 15431 17564 15476 17592
rect 11379 17561 11391 17564
rect 11333 17555 11391 17561
rect 15470 17552 15476 17564
rect 15528 17552 15534 17604
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 15620 17564 15665 17592
rect 15620 17552 15626 17564
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 16853 17595 16911 17601
rect 16356 17564 16401 17592
rect 16356 17552 16362 17564
rect 16853 17561 16865 17595
rect 16899 17561 16911 17595
rect 16853 17555 16911 17561
rect 12986 17524 12992 17536
rect 12947 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 14369 17527 14427 17533
rect 14369 17493 14381 17527
rect 14415 17524 14427 17527
rect 16482 17524 16488 17536
rect 14415 17496 16488 17524
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 16482 17484 16488 17496
rect 16540 17484 16546 17536
rect 16868 17524 16896 17555
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 17497 17595 17555 17601
rect 17497 17592 17509 17595
rect 17092 17564 17509 17592
rect 17092 17552 17098 17564
rect 17497 17561 17509 17564
rect 17543 17561 17555 17595
rect 17497 17555 17555 17561
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17561 18107 17595
rect 18049 17555 18107 17561
rect 18064 17524 18092 17555
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 19613 17595 19671 17601
rect 18196 17564 19472 17592
rect 18196 17552 18202 17564
rect 18230 17524 18236 17536
rect 16868 17496 18236 17524
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18785 17527 18843 17533
rect 18785 17493 18797 17527
rect 18831 17524 18843 17527
rect 19242 17524 19248 17536
rect 18831 17496 19248 17524
rect 18831 17493 18843 17496
rect 18785 17487 18843 17493
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 19444 17524 19472 17564
rect 19613 17561 19625 17595
rect 19659 17561 19671 17595
rect 19613 17555 19671 17561
rect 20165 17595 20223 17601
rect 20165 17561 20177 17595
rect 20211 17592 20223 17595
rect 20346 17592 20352 17604
rect 20211 17564 20352 17592
rect 20211 17561 20223 17564
rect 20165 17555 20223 17561
rect 19628 17524 19656 17555
rect 20346 17552 20352 17564
rect 20404 17552 20410 17604
rect 21450 17552 21456 17604
rect 21508 17592 21514 17604
rect 21508 17564 21553 17592
rect 21508 17552 21514 17564
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 24673 17595 24731 17601
rect 24673 17592 24685 17595
rect 23072 17564 23117 17592
rect 23216 17564 24685 17592
rect 23072 17552 23078 17564
rect 20714 17524 20720 17536
rect 19444 17496 19656 17524
rect 20675 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17524 20778 17536
rect 22094 17524 22100 17536
rect 20772 17496 22100 17524
rect 20772 17484 20778 17496
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 22370 17484 22376 17536
rect 22428 17524 22434 17536
rect 23216 17524 23244 17564
rect 24673 17561 24685 17564
rect 24719 17561 24731 17595
rect 24673 17555 24731 17561
rect 24765 17595 24823 17601
rect 24765 17561 24777 17595
rect 24811 17592 24823 17595
rect 25590 17592 25596 17604
rect 24811 17564 25596 17592
rect 24811 17561 24823 17564
rect 24765 17555 24823 17561
rect 25590 17552 25596 17564
rect 25648 17552 25654 17604
rect 25685 17595 25743 17601
rect 25685 17561 25697 17595
rect 25731 17592 25743 17595
rect 26252 17592 26280 17700
rect 27433 17697 27445 17700
rect 27479 17728 27491 17731
rect 27540 17728 27568 17836
rect 28350 17824 28356 17836
rect 28408 17824 28414 17876
rect 27890 17756 27896 17808
rect 27948 17796 27954 17808
rect 28629 17799 28687 17805
rect 28629 17796 28641 17799
rect 27948 17768 28641 17796
rect 27948 17756 27954 17768
rect 28629 17765 28641 17768
rect 28675 17765 28687 17799
rect 28629 17759 28687 17765
rect 27479 17700 27568 17728
rect 27479 17697 27491 17700
rect 27433 17691 27491 17697
rect 27706 17688 27712 17740
rect 27764 17728 27770 17740
rect 28445 17731 28503 17737
rect 28445 17728 28457 17731
rect 27764 17700 28457 17728
rect 27764 17688 27770 17700
rect 28445 17697 28457 17700
rect 28491 17697 28503 17731
rect 28445 17691 28503 17697
rect 28261 17663 28319 17669
rect 28261 17629 28273 17663
rect 28307 17629 28319 17663
rect 28261 17623 28319 17629
rect 25731 17564 26280 17592
rect 25731 17561 25743 17564
rect 25685 17555 25743 17561
rect 22428 17496 23244 17524
rect 22428 17484 22434 17496
rect 24302 17484 24308 17536
rect 24360 17524 24366 17536
rect 25700 17524 25728 17555
rect 27522 17552 27528 17604
rect 27580 17592 27586 17604
rect 27617 17595 27675 17601
rect 27617 17592 27629 17595
rect 27580 17564 27629 17592
rect 27580 17552 27586 17564
rect 27617 17561 27629 17564
rect 27663 17561 27675 17595
rect 27617 17555 27675 17561
rect 27706 17552 27712 17604
rect 27764 17592 27770 17604
rect 27764 17564 27809 17592
rect 27764 17552 27770 17564
rect 24360 17496 25728 17524
rect 24360 17484 24366 17496
rect 26602 17484 26608 17536
rect 26660 17524 26666 17536
rect 28276 17524 28304 17623
rect 26660 17496 28304 17524
rect 26660 17484 26666 17496
rect 28994 17484 29000 17536
rect 29052 17524 29058 17536
rect 29733 17527 29791 17533
rect 29733 17524 29745 17527
rect 29052 17496 29745 17524
rect 29052 17484 29058 17496
rect 29733 17493 29745 17496
rect 29779 17493 29791 17527
rect 29733 17487 29791 17493
rect 1104 17434 36892 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 36892 17434
rect 1104 17360 36892 17382
rect 9950 17320 9956 17332
rect 9911 17292 9956 17320
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 16114 17320 16120 17332
rect 12406 17292 16120 17320
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9968 17184 9996 17280
rect 9539 17156 9996 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 11330 17144 11336 17196
rect 11388 17184 11394 17196
rect 12161 17187 12219 17193
rect 12161 17184 12173 17187
rect 11388 17156 12173 17184
rect 11388 17144 11394 17156
rect 12161 17153 12173 17156
rect 12207 17184 12219 17187
rect 12406 17184 12434 17292
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16298 17320 16304 17332
rect 16255 17292 16304 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16942 17320 16948 17332
rect 16903 17292 16948 17320
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20220 17292 21036 17320
rect 20220 17280 20226 17292
rect 15105 17255 15163 17261
rect 15105 17252 15117 17255
rect 14844 17224 15117 17252
rect 13262 17184 13268 17196
rect 12207 17156 12434 17184
rect 13223 17156 13268 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17184 13507 17187
rect 14090 17184 14096 17196
rect 13495 17156 14096 17184
rect 13495 17153 13507 17156
rect 13449 17147 13507 17153
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14277 17187 14335 17193
rect 14277 17184 14289 17187
rect 14240 17156 14289 17184
rect 14240 17144 14246 17156
rect 14277 17153 14289 17156
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 14844 17184 14872 17224
rect 15105 17221 15117 17224
rect 15151 17221 15163 17255
rect 17497 17255 17555 17261
rect 17497 17252 17509 17255
rect 15105 17215 15163 17221
rect 15764 17224 17509 17252
rect 14792 17156 14872 17184
rect 14792 17144 14798 17156
rect 13078 17076 13084 17128
rect 13136 17116 13142 17128
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 13136 17088 15025 17116
rect 13136 17076 13142 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 15102 17076 15108 17128
rect 15160 17116 15166 17128
rect 15289 17119 15347 17125
rect 15289 17116 15301 17119
rect 15160 17088 15301 17116
rect 15160 17076 15166 17088
rect 15289 17085 15301 17088
rect 15335 17116 15347 17119
rect 15764 17116 15792 17224
rect 17497 17221 17509 17224
rect 17543 17221 17555 17255
rect 18046 17252 18052 17264
rect 18007 17224 18052 17252
rect 17497 17215 17555 17221
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 15896 17156 16129 17184
rect 15896 17144 15902 17156
rect 16117 17153 16129 17156
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16816 17156 16865 17184
rect 16816 17144 16822 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 15335 17088 15792 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 1857 17051 1915 17057
rect 1857 17017 1869 17051
rect 1903 17048 1915 17051
rect 2590 17048 2596 17060
rect 1903 17020 2596 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 2590 17008 2596 17020
rect 2648 17008 2654 17060
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 13354 17048 13360 17060
rect 12299 17020 13360 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 14182 17008 14188 17060
rect 14240 17048 14246 17060
rect 16758 17048 16764 17060
rect 14240 17020 16764 17048
rect 14240 17008 14246 17020
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 17512 17048 17540 17215
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 19242 17252 19248 17264
rect 19203 17224 19248 17252
rect 19242 17212 19248 17224
rect 19300 17212 19306 17264
rect 19337 17255 19395 17261
rect 19337 17221 19349 17255
rect 19383 17252 19395 17255
rect 20714 17252 20720 17264
rect 19383 17224 20720 17252
rect 19383 17221 19395 17224
rect 19337 17215 19395 17221
rect 20714 17212 20720 17224
rect 20772 17212 20778 17264
rect 20898 17252 20904 17264
rect 20859 17224 20904 17252
rect 20898 17212 20904 17224
rect 20956 17212 20962 17264
rect 21008 17261 21036 17292
rect 21192 17292 23336 17320
rect 20993 17255 21051 17261
rect 20993 17221 21005 17255
rect 21039 17221 21051 17255
rect 20993 17215 21051 17221
rect 20346 17184 20352 17196
rect 20307 17156 20352 17184
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 18138 17116 18144 17128
rect 18099 17088 18144 17116
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 21192 17116 21220 17292
rect 23308 17261 23336 17292
rect 24854 17280 24860 17332
rect 24912 17320 24918 17332
rect 26053 17323 26111 17329
rect 26053 17320 26065 17323
rect 24912 17292 26065 17320
rect 24912 17280 24918 17292
rect 26053 17289 26065 17292
rect 26099 17289 26111 17323
rect 26053 17283 26111 17289
rect 27614 17280 27620 17332
rect 27672 17320 27678 17332
rect 29730 17320 29736 17332
rect 27672 17292 29736 17320
rect 27672 17280 27678 17292
rect 29730 17280 29736 17292
rect 29788 17280 29794 17332
rect 22189 17255 22247 17261
rect 22189 17221 22201 17255
rect 22235 17252 22247 17255
rect 23293 17255 23351 17261
rect 22235 17224 23152 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 18248 17088 21220 17116
rect 18248 17048 18276 17088
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22830 17116 22836 17128
rect 22152 17088 22197 17116
rect 22572 17088 22836 17116
rect 22152 17076 22158 17088
rect 17512 17020 18276 17048
rect 18785 17051 18843 17057
rect 18785 17017 18797 17051
rect 18831 17017 18843 17051
rect 18785 17011 18843 17017
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 5408 16952 9321 16980
rect 5408 16940 5414 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 11149 16983 11207 16989
rect 11149 16949 11161 16983
rect 11195 16980 11207 16983
rect 11330 16980 11336 16992
rect 11195 16952 11336 16980
rect 11195 16949 11207 16952
rect 11149 16943 11207 16949
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 13081 16983 13139 16989
rect 13081 16949 13093 16983
rect 13127 16980 13139 16983
rect 13446 16980 13452 16992
rect 13127 16952 13452 16980
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 14369 16983 14427 16989
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 16206 16980 16212 16992
rect 14415 16952 16212 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 18800 16980 18828 17011
rect 18874 17008 18880 17060
rect 18932 17048 18938 17060
rect 22572 17048 22600 17088
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 23124 17116 23152 17224
rect 23293 17221 23305 17255
rect 23339 17221 23351 17255
rect 23293 17215 23351 17221
rect 23385 17255 23443 17261
rect 23385 17221 23397 17255
rect 23431 17252 23443 17255
rect 24946 17252 24952 17264
rect 23431 17224 24716 17252
rect 24907 17224 24952 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 23474 17116 23480 17128
rect 23124 17088 23480 17116
rect 23474 17076 23480 17088
rect 23532 17076 23538 17128
rect 24302 17116 24308 17128
rect 24263 17088 24308 17116
rect 24302 17076 24308 17088
rect 24360 17076 24366 17128
rect 18932 17020 22600 17048
rect 22649 17051 22707 17057
rect 18932 17008 18938 17020
rect 22649 17017 22661 17051
rect 22695 17048 22707 17051
rect 23566 17048 23572 17060
rect 22695 17020 23572 17048
rect 22695 17017 22707 17020
rect 22649 17011 22707 17017
rect 23566 17008 23572 17020
rect 23624 17048 23630 17060
rect 24578 17048 24584 17060
rect 23624 17020 24584 17048
rect 23624 17008 23630 17020
rect 24578 17008 24584 17020
rect 24636 17008 24642 17060
rect 24688 17048 24716 17224
rect 24946 17212 24952 17224
rect 25004 17212 25010 17264
rect 25590 17212 25596 17264
rect 25648 17252 25654 17264
rect 29178 17252 29184 17264
rect 25648 17224 29184 17252
rect 25648 17212 25654 17224
rect 29178 17212 29184 17224
rect 29236 17212 29242 17264
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 24857 17119 24915 17125
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 25038 17116 25044 17128
rect 24903 17088 25044 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 25038 17076 25044 17088
rect 25096 17116 25102 17128
rect 25682 17116 25688 17128
rect 25096 17088 25688 17116
rect 25096 17076 25102 17088
rect 25682 17076 25688 17088
rect 25740 17076 25746 17128
rect 26160 17116 26188 17147
rect 26602 17144 26608 17196
rect 26660 17184 26666 17196
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 26660 17156 27353 17184
rect 26660 17144 26666 17156
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17184 28043 17187
rect 28810 17184 28816 17196
rect 28031 17156 28816 17184
rect 28031 17153 28043 17156
rect 27985 17147 28043 17153
rect 28810 17144 28816 17156
rect 28868 17144 28874 17196
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29089 17187 29147 17193
rect 29089 17184 29101 17187
rect 29052 17156 29101 17184
rect 29052 17144 29058 17156
rect 29089 17153 29101 17156
rect 29135 17153 29147 17187
rect 36081 17187 36139 17193
rect 36081 17184 36093 17187
rect 29089 17147 29147 17153
rect 31726 17156 36093 17184
rect 28626 17116 28632 17128
rect 26160 17088 28028 17116
rect 28587 17088 28632 17116
rect 25222 17048 25228 17060
rect 24688 17020 25228 17048
rect 25222 17008 25228 17020
rect 25280 17008 25286 17060
rect 25409 17051 25467 17057
rect 25409 17017 25421 17051
rect 25455 17048 25467 17051
rect 25590 17048 25596 17060
rect 25455 17020 25596 17048
rect 25455 17017 25467 17020
rect 25409 17011 25467 17017
rect 25590 17008 25596 17020
rect 25648 17008 25654 17060
rect 27893 17051 27951 17057
rect 27893 17048 27905 17051
rect 25700 17020 27905 17048
rect 16724 16952 18828 16980
rect 16724 16940 16730 16952
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 21082 16980 21088 16992
rect 20404 16952 21088 16980
rect 20404 16940 20410 16952
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 23290 16940 23296 16992
rect 23348 16980 23354 16992
rect 25700 16980 25728 17020
rect 27893 17017 27905 17020
rect 27939 17017 27951 17051
rect 28000 17048 28028 17088
rect 28626 17076 28632 17088
rect 28684 17076 28690 17128
rect 29273 17051 29331 17057
rect 28000 17020 28764 17048
rect 27893 17011 27951 17017
rect 28736 16992 28764 17020
rect 29273 17017 29285 17051
rect 29319 17048 29331 17051
rect 31726 17048 31754 17156
rect 36081 17153 36093 17156
rect 36127 17153 36139 17187
rect 36081 17147 36139 17153
rect 36262 17048 36268 17060
rect 29319 17020 31754 17048
rect 36223 17020 36268 17048
rect 29319 17017 29331 17020
rect 29273 17011 29331 17017
rect 36262 17008 36268 17020
rect 36320 17008 36326 17060
rect 23348 16952 25728 16980
rect 23348 16940 23354 16952
rect 26970 16940 26976 16992
rect 27028 16980 27034 16992
rect 27249 16983 27307 16989
rect 27249 16980 27261 16983
rect 27028 16952 27261 16980
rect 27028 16940 27034 16952
rect 27249 16949 27261 16952
rect 27295 16949 27307 16983
rect 27249 16943 27307 16949
rect 28718 16940 28724 16992
rect 28776 16980 28782 16992
rect 29733 16983 29791 16989
rect 29733 16980 29745 16983
rect 28776 16952 29745 16980
rect 28776 16940 28782 16952
rect 29733 16949 29745 16952
rect 29779 16949 29791 16983
rect 30282 16980 30288 16992
rect 30243 16952 30288 16980
rect 29733 16943 29791 16949
rect 30282 16940 30288 16952
rect 30340 16940 30346 16992
rect 1104 16890 36892 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36892 16890
rect 1104 16816 36892 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 13446 16776 13452 16788
rect 13407 16748 13452 16776
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 15194 16776 15200 16788
rect 13556 16748 15200 16776
rect 13556 16708 13584 16748
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 17770 16776 17776 16788
rect 15620 16748 17776 16776
rect 15620 16736 15626 16748
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 20622 16776 20628 16788
rect 17880 16748 20628 16776
rect 15010 16708 15016 16720
rect 12636 16680 13584 16708
rect 14971 16680 15016 16708
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 11256 16572 11284 16603
rect 12636 16581 12664 16680
rect 15010 16668 15016 16680
rect 15068 16708 15074 16720
rect 16209 16711 16267 16717
rect 16209 16708 16221 16711
rect 15068 16680 16221 16708
rect 15068 16668 15074 16680
rect 16209 16677 16221 16680
rect 16255 16677 16267 16711
rect 17678 16708 17684 16720
rect 16209 16671 16267 16677
rect 16546 16680 17684 16708
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 13044 16612 13277 16640
rect 13044 16600 13050 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 16546 16640 16574 16680
rect 17678 16668 17684 16680
rect 17736 16668 17742 16720
rect 13265 16603 13323 16609
rect 14936 16612 16574 16640
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 6788 16544 11805 16572
rect 6788 16532 6794 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16541 12679 16575
rect 13078 16572 13084 16584
rect 13039 16544 13084 16572
rect 12621 16535 12679 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 14277 16575 14335 16581
rect 14277 16572 14289 16575
rect 13188 16544 14289 16572
rect 11885 16507 11943 16513
rect 11885 16473 11897 16507
rect 11931 16504 11943 16507
rect 13096 16504 13124 16532
rect 11931 16476 13124 16504
rect 11931 16473 11943 16476
rect 11885 16467 11943 16473
rect 2130 16396 2136 16448
rect 2188 16436 2194 16448
rect 2682 16436 2688 16448
rect 2188 16408 2688 16436
rect 2188 16396 2194 16408
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 12526 16436 12532 16448
rect 12487 16408 12532 16436
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 12986 16396 12992 16448
rect 13044 16436 13050 16448
rect 13188 16436 13216 16544
rect 14277 16541 14289 16544
rect 14323 16572 14335 16575
rect 14936 16572 14964 16612
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 16761 16643 16819 16649
rect 16761 16640 16773 16643
rect 16724 16612 16773 16640
rect 16724 16600 16730 16612
rect 16761 16609 16773 16612
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17880 16640 17908 16748
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 20956 16748 21189 16776
rect 20956 16736 20962 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 29822 16776 29828 16788
rect 29783 16748 29828 16776
rect 21177 16739 21235 16745
rect 29822 16736 29828 16748
rect 29880 16736 29886 16788
rect 18230 16668 18236 16720
rect 18288 16708 18294 16720
rect 22922 16708 22928 16720
rect 18288 16680 22928 16708
rect 18288 16668 18294 16680
rect 22922 16668 22928 16680
rect 22980 16668 22986 16720
rect 24210 16708 24216 16720
rect 23492 16680 24216 16708
rect 20254 16640 20260 16652
rect 17000 16612 17908 16640
rect 20215 16612 20260 16640
rect 17000 16600 17006 16612
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 20530 16640 20536 16652
rect 20491 16612 20536 16640
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 21542 16640 21548 16652
rect 21284 16612 21548 16640
rect 17678 16572 17684 16584
rect 14323 16544 14964 16572
rect 17639 16544 17684 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 18690 16572 18696 16584
rect 18651 16544 18696 16572
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 21284 16581 21312 16612
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 22833 16643 22891 16649
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 23492 16640 23520 16680
rect 24210 16668 24216 16680
rect 24268 16668 24274 16720
rect 24578 16668 24584 16720
rect 24636 16708 24642 16720
rect 24636 16680 24992 16708
rect 24636 16668 24642 16680
rect 24964 16649 24992 16680
rect 26602 16668 26608 16720
rect 26660 16708 26666 16720
rect 26660 16680 29040 16708
rect 26660 16668 26666 16680
rect 22879 16612 23520 16640
rect 24949 16643 25007 16649
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 24949 16609 24961 16643
rect 24995 16609 25007 16643
rect 25774 16640 25780 16652
rect 25735 16612 25780 16640
rect 24949 16603 25007 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 26418 16640 26424 16652
rect 26379 16612 26424 16640
rect 26418 16600 26424 16612
rect 26476 16640 26482 16652
rect 27617 16643 27675 16649
rect 27617 16640 27629 16643
rect 26476 16612 27629 16640
rect 26476 16600 26482 16612
rect 27617 16609 27629 16612
rect 27663 16609 27675 16643
rect 28258 16640 28264 16652
rect 28219 16612 28264 16640
rect 27617 16603 27675 16609
rect 28258 16600 28264 16612
rect 28316 16600 28322 16652
rect 29012 16640 29040 16680
rect 30282 16640 30288 16652
rect 29012 16612 30288 16640
rect 29012 16581 29040 16612
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 21269 16535 21327 16541
rect 23308 16544 23581 16572
rect 13906 16464 13912 16516
rect 13964 16504 13970 16516
rect 15473 16507 15531 16513
rect 15473 16504 15485 16507
rect 13964 16476 15485 16504
rect 13964 16464 13970 16476
rect 15473 16473 15485 16476
rect 15519 16473 15531 16507
rect 15473 16467 15531 16473
rect 15565 16507 15623 16513
rect 15565 16473 15577 16507
rect 15611 16504 15623 16507
rect 15838 16504 15844 16516
rect 15611 16476 15844 16504
rect 15611 16473 15623 16476
rect 15565 16467 15623 16473
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 16669 16507 16727 16513
rect 16669 16473 16681 16507
rect 16715 16473 16727 16507
rect 16669 16467 16727 16473
rect 13044 16408 13216 16436
rect 14461 16439 14519 16445
rect 13044 16396 13050 16408
rect 14461 16405 14473 16439
rect 14507 16436 14519 16439
rect 15010 16436 15016 16448
rect 14507 16408 15016 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 16684 16436 16712 16467
rect 18874 16464 18880 16516
rect 18932 16504 18938 16516
rect 20162 16504 20168 16516
rect 18932 16476 20168 16504
rect 18932 16464 18938 16476
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 20438 16504 20444 16516
rect 20399 16476 20444 16504
rect 20438 16464 20444 16476
rect 20496 16464 20502 16516
rect 20530 16464 20536 16516
rect 20588 16504 20594 16516
rect 22189 16507 22247 16513
rect 22189 16504 22201 16507
rect 20588 16476 22201 16504
rect 20588 16464 20594 16476
rect 22189 16473 22201 16476
rect 22235 16473 22247 16507
rect 22738 16504 22744 16516
rect 22699 16476 22744 16504
rect 22189 16467 22247 16473
rect 16942 16436 16948 16448
rect 16684 16408 16948 16436
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 18785 16439 18843 16445
rect 18785 16405 18797 16439
rect 18831 16436 18843 16439
rect 20070 16436 20076 16448
rect 18831 16408 20076 16436
rect 18831 16405 18843 16408
rect 18785 16399 18843 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 22204 16436 22232 16467
rect 22738 16464 22744 16476
rect 22796 16464 22802 16516
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 23308 16504 23336 16544
rect 23569 16541 23581 16544
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 23474 16504 23480 16516
rect 22888 16476 23336 16504
rect 23435 16476 23480 16504
rect 22888 16464 22894 16476
rect 23474 16464 23480 16476
rect 23532 16464 23538 16516
rect 25038 16464 25044 16516
rect 25096 16504 25102 16516
rect 25096 16476 25141 16504
rect 25096 16464 25102 16476
rect 25406 16464 25412 16516
rect 25464 16504 25470 16516
rect 26970 16504 26976 16516
rect 25464 16476 26648 16504
rect 26931 16476 26976 16504
rect 25464 16464 25470 16476
rect 25590 16436 25596 16448
rect 22204 16408 25596 16436
rect 25590 16396 25596 16408
rect 25648 16396 25654 16448
rect 26620 16436 26648 16476
rect 26970 16464 26976 16476
rect 27028 16464 27034 16516
rect 27062 16464 27068 16516
rect 27120 16504 27126 16516
rect 28166 16504 28172 16516
rect 27120 16476 27165 16504
rect 28127 16476 28172 16504
rect 27120 16464 27126 16476
rect 28166 16464 28172 16476
rect 28224 16464 28230 16516
rect 30282 16504 30288 16516
rect 28276 16476 30288 16504
rect 28276 16436 28304 16476
rect 30282 16464 30288 16476
rect 30340 16464 30346 16516
rect 26620 16408 28304 16436
rect 28350 16396 28356 16448
rect 28408 16436 28414 16448
rect 28905 16439 28963 16445
rect 28905 16436 28917 16439
rect 28408 16408 28917 16436
rect 28408 16396 28414 16408
rect 28905 16405 28917 16408
rect 28951 16405 28963 16439
rect 28905 16399 28963 16405
rect 31021 16439 31079 16445
rect 31021 16405 31033 16439
rect 31067 16436 31079 16439
rect 31110 16436 31116 16448
rect 31067 16408 31116 16436
rect 31067 16405 31079 16408
rect 31021 16399 31079 16405
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 1104 16346 36892 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 36892 16346
rect 1104 16272 36892 16294
rect 2314 16232 2320 16244
rect 2275 16204 2320 16232
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10008 16204 11069 16232
rect 10008 16192 10014 16204
rect 11057 16201 11069 16204
rect 11103 16232 11115 16235
rect 12342 16232 12348 16244
rect 11103 16204 12348 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 12584 16204 17172 16232
rect 12584 16192 12590 16204
rect 15289 16167 15347 16173
rect 15289 16164 15301 16167
rect 12544 16136 15301 16164
rect 1854 16096 1860 16108
rect 1815 16068 1860 16096
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 2682 16096 2688 16108
rect 2547 16068 2688 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 12544 16105 12572 16136
rect 15289 16133 15301 16136
rect 15335 16133 15347 16167
rect 15289 16127 15347 16133
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 17144 16164 17172 16204
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 19242 16232 19248 16244
rect 18196 16204 19248 16232
rect 18196 16192 18202 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 22370 16192 22376 16244
rect 22428 16232 22434 16244
rect 27246 16232 27252 16244
rect 22428 16204 22508 16232
rect 22428 16192 22434 16204
rect 17083 16136 17172 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 18046 16124 18052 16176
rect 18104 16164 18110 16176
rect 22480 16173 22508 16204
rect 24228 16204 27252 16232
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 18104 16136 19441 16164
rect 18104 16124 18110 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 22465 16167 22523 16173
rect 22465 16133 22477 16167
rect 22511 16133 22523 16167
rect 22465 16127 22523 16133
rect 23017 16167 23075 16173
rect 23017 16133 23029 16167
rect 23063 16164 23075 16167
rect 23566 16164 23572 16176
rect 23063 16136 23572 16164
rect 23063 16133 23075 16136
rect 23017 16127 23075 16133
rect 23566 16124 23572 16136
rect 23624 16124 23630 16176
rect 24228 16173 24256 16204
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 27890 16232 27896 16244
rect 27851 16204 27896 16232
rect 27890 16192 27896 16204
rect 27948 16192 27954 16244
rect 28166 16192 28172 16244
rect 28224 16232 28230 16244
rect 29089 16235 29147 16241
rect 29089 16232 29101 16235
rect 28224 16204 29101 16232
rect 28224 16192 28230 16204
rect 29089 16201 29101 16204
rect 29135 16201 29147 16235
rect 30282 16232 30288 16244
rect 30243 16204 30288 16232
rect 29089 16195 29147 16201
rect 30282 16192 30288 16204
rect 30340 16192 30346 16244
rect 31297 16235 31355 16241
rect 31297 16201 31309 16235
rect 31343 16232 31355 16235
rect 31343 16204 31754 16232
rect 31343 16201 31355 16204
rect 31297 16195 31355 16201
rect 24213 16167 24271 16173
rect 24213 16133 24225 16167
rect 24259 16133 24271 16167
rect 24213 16127 24271 16133
rect 24302 16124 24308 16176
rect 24360 16164 24366 16176
rect 25406 16164 25412 16176
rect 24360 16136 25412 16164
rect 24360 16124 24366 16136
rect 25406 16124 25412 16136
rect 25464 16124 25470 16176
rect 25501 16167 25559 16173
rect 25501 16133 25513 16167
rect 25547 16164 25559 16167
rect 26602 16164 26608 16176
rect 25547 16136 26608 16164
rect 25547 16133 25559 16136
rect 25501 16127 25559 16133
rect 26602 16124 26608 16136
rect 26660 16124 26666 16176
rect 26712 16136 29684 16164
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 12676 16068 12721 16096
rect 13096 16068 13277 16096
rect 12676 16056 12682 16068
rect 2222 15988 2228 16040
rect 2280 16028 2286 16040
rect 11885 16031 11943 16037
rect 11885 16028 11897 16031
rect 2280 16000 11897 16028
rect 2280 15988 2286 16000
rect 11885 15997 11897 16000
rect 11931 16028 11943 16031
rect 12986 16028 12992 16040
rect 11931 16000 12992 16028
rect 11931 15997 11943 16000
rect 11885 15991 11943 15997
rect 12986 15988 12992 16000
rect 13044 15988 13050 16040
rect 2038 15920 2044 15972
rect 2096 15960 2102 15972
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 2096 15932 10517 15960
rect 2096 15920 2102 15932
rect 10505 15929 10517 15932
rect 10551 15960 10563 15963
rect 11606 15960 11612 15972
rect 10551 15932 11612 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 11606 15920 11612 15932
rect 11664 15920 11670 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2682 15852 2688 15904
rect 2740 15892 2746 15904
rect 2961 15895 3019 15901
rect 2961 15892 2973 15895
rect 2740 15864 2973 15892
rect 2740 15852 2746 15864
rect 2961 15861 2973 15864
rect 3007 15861 3019 15895
rect 13096 15892 13124 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13412 16068 14197 16096
rect 13412 16056 13418 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14366 16096 14372 16108
rect 14327 16068 14372 16096
rect 14185 16059 14243 16065
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 18874 16096 18880 16108
rect 18739 16068 18880 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 20346 16056 20352 16108
rect 20404 16096 20410 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20404 16068 20545 16096
rect 20404 16056 20410 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 21361 16099 21419 16105
rect 21361 16065 21373 16099
rect 21407 16096 21419 16099
rect 21818 16096 21824 16108
rect 21407 16068 21824 16096
rect 21407 16065 21419 16068
rect 21361 16059 21419 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 13446 15988 13452 16040
rect 13504 16028 13510 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13504 16000 13737 16028
rect 13504 15988 13510 16000
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 16028 15255 16031
rect 15286 16028 15292 16040
rect 15243 16000 15292 16028
rect 15243 15997 15255 16000
rect 15197 15991 15255 15997
rect 15286 15988 15292 16000
rect 15344 16028 15350 16040
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 15344 16000 16957 16028
rect 15344 15988 15350 16000
rect 16945 15997 16957 16000
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 17589 16031 17647 16037
rect 17589 15997 17601 16031
rect 17635 16028 17647 16031
rect 17635 16000 18644 16028
rect 17635 15997 17647 16000
rect 17589 15991 17647 15997
rect 13173 15963 13231 15969
rect 13173 15929 13185 15963
rect 13219 15960 13231 15963
rect 15102 15960 15108 15972
rect 13219 15932 15108 15960
rect 13219 15929 13231 15932
rect 13173 15923 13231 15929
rect 15102 15920 15108 15932
rect 15160 15920 15166 15972
rect 15746 15960 15752 15972
rect 15707 15932 15752 15960
rect 15746 15920 15752 15932
rect 15804 15920 15810 15972
rect 15838 15920 15844 15972
rect 15896 15960 15902 15972
rect 18506 15960 18512 15972
rect 15896 15932 18276 15960
rect 18467 15932 18512 15960
rect 15896 15920 15902 15932
rect 14642 15892 14648 15904
rect 13096 15864 14648 15892
rect 2961 15855 3019 15861
rect 14642 15852 14648 15864
rect 14700 15892 14706 15904
rect 15930 15892 15936 15904
rect 14700 15864 15936 15892
rect 14700 15852 14706 15864
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 18138 15892 18144 15904
rect 16264 15864 18144 15892
rect 16264 15852 16270 15864
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 18248 15892 18276 15932
rect 18506 15920 18512 15932
rect 18564 15920 18570 15972
rect 18616 15960 18644 16000
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19392 16000 19437 16028
rect 19392 15988 19398 16000
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 22646 16028 22652 16040
rect 19576 16000 22652 16028
rect 19576 15988 19582 16000
rect 22646 15988 22652 16000
rect 22704 15988 22710 16040
rect 23109 16031 23167 16037
rect 23109 15997 23121 16031
rect 23155 16028 23167 16031
rect 23290 16028 23296 16040
rect 23155 16000 23296 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 23290 15988 23296 16000
rect 23348 15988 23354 16040
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 23532 16000 23673 16028
rect 23532 15988 23538 16000
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 24302 16028 24308 16040
rect 24263 16000 24308 16028
rect 23661 15991 23719 15997
rect 19889 15963 19947 15969
rect 19889 15960 19901 15963
rect 18616 15932 19901 15960
rect 19889 15929 19901 15932
rect 19935 15960 19947 15963
rect 20346 15960 20352 15972
rect 19935 15932 20352 15960
rect 19935 15929 19947 15932
rect 19889 15923 19947 15929
rect 20346 15920 20352 15932
rect 20404 15920 20410 15972
rect 20625 15963 20683 15969
rect 20625 15929 20637 15963
rect 20671 15960 20683 15963
rect 22462 15960 22468 15972
rect 20671 15932 22468 15960
rect 20671 15929 20683 15932
rect 20625 15923 20683 15929
rect 22462 15920 22468 15932
rect 22520 15920 22526 15972
rect 20806 15892 20812 15904
rect 18248 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 22664 15892 22692 15988
rect 23676 15960 23704 15991
rect 24302 15988 24308 16000
rect 24360 15988 24366 16040
rect 25409 16031 25467 16037
rect 25409 15997 25421 16031
rect 25455 15997 25467 16031
rect 25774 16028 25780 16040
rect 25735 16000 25780 16028
rect 25409 15991 25467 15997
rect 25424 15960 25452 15991
rect 25774 15988 25780 16000
rect 25832 15988 25838 16040
rect 25866 15988 25872 16040
rect 25924 16028 25930 16040
rect 26712 16028 26740 16136
rect 27338 16096 27344 16108
rect 27299 16068 27344 16096
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 28350 16096 28356 16108
rect 28311 16068 28356 16096
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28537 16099 28595 16105
rect 28537 16065 28549 16099
rect 28583 16096 28595 16099
rect 28626 16096 28632 16108
rect 28583 16068 28632 16096
rect 28583 16065 28595 16068
rect 28537 16059 28595 16065
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 29656 16105 29684 16136
rect 29181 16099 29239 16105
rect 29181 16065 29193 16099
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 29641 16099 29699 16105
rect 29641 16065 29653 16099
rect 29687 16065 29699 16099
rect 31110 16096 31116 16108
rect 31071 16068 31116 16096
rect 29641 16059 29699 16065
rect 25924 16000 26740 16028
rect 29196 16028 29224 16059
rect 31110 16056 31116 16068
rect 31168 16056 31174 16108
rect 31726 16096 31754 16204
rect 36081 16099 36139 16105
rect 36081 16096 36093 16099
rect 31726 16068 36093 16096
rect 36081 16065 36093 16068
rect 36127 16065 36139 16099
rect 36081 16059 36139 16065
rect 29914 16028 29920 16040
rect 29196 16000 29920 16028
rect 25924 15988 25930 16000
rect 29914 15988 29920 16000
rect 29972 15988 29978 16040
rect 23676 15932 25452 15960
rect 27522 15920 27528 15972
rect 27580 15960 27586 15972
rect 29733 15963 29791 15969
rect 29733 15960 29745 15963
rect 27580 15932 29745 15960
rect 27580 15920 27586 15932
rect 29733 15929 29745 15932
rect 29779 15929 29791 15963
rect 29733 15923 29791 15929
rect 23106 15892 23112 15904
rect 22664 15864 23112 15892
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 24302 15852 24308 15904
rect 24360 15892 24366 15904
rect 27062 15892 27068 15904
rect 24360 15864 27068 15892
rect 24360 15852 24366 15864
rect 27062 15852 27068 15864
rect 27120 15892 27126 15904
rect 27249 15895 27307 15901
rect 27249 15892 27261 15895
rect 27120 15864 27261 15892
rect 27120 15852 27126 15864
rect 27249 15861 27261 15864
rect 27295 15861 27307 15895
rect 27249 15855 27307 15861
rect 27338 15852 27344 15904
rect 27396 15892 27402 15904
rect 29822 15892 29828 15904
rect 27396 15864 29828 15892
rect 27396 15852 27402 15864
rect 29822 15852 29828 15864
rect 29880 15852 29886 15904
rect 36262 15892 36268 15904
rect 36223 15864 36268 15892
rect 36262 15852 36268 15864
rect 36320 15852 36326 15904
rect 1104 15802 36892 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36892 15802
rect 1104 15728 36892 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 3973 15691 4031 15697
rect 3973 15688 3985 15691
rect 1912 15660 3985 15688
rect 1912 15648 1918 15660
rect 3973 15657 3985 15660
rect 4019 15657 4031 15691
rect 3973 15651 4031 15657
rect 4709 15691 4767 15697
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 6730 15688 6736 15700
rect 4755 15660 6736 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4724 15484 4752 15651
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 15746 15648 15752 15700
rect 15804 15688 15810 15700
rect 15804 15660 16712 15688
rect 15804 15648 15810 15660
rect 11146 15620 11152 15632
rect 11059 15592 11152 15620
rect 11146 15580 11152 15592
rect 11204 15620 11210 15632
rect 11204 15592 14320 15620
rect 11204 15580 11210 15592
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15552 10655 15555
rect 10643 15524 12296 15552
rect 10643 15521 10655 15524
rect 10597 15515 10655 15521
rect 11606 15484 11612 15496
rect 4203 15456 4752 15484
rect 11567 15456 11612 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 12268 15493 12296 15524
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 13630 15552 13636 15564
rect 12400 15524 12940 15552
rect 13591 15524 13636 15552
rect 12400 15512 12406 15524
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12710 15484 12716 15496
rect 12299 15456 12716 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 12912 15493 12940 15524
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 13722 15484 13728 15496
rect 13587 15456 13728 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14292 15493 14320 15592
rect 14826 15580 14832 15632
rect 14884 15620 14890 15632
rect 16574 15620 16580 15632
rect 14884 15592 16580 15620
rect 14884 15580 14890 15592
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 16684 15620 16712 15660
rect 17310 15648 17316 15700
rect 17368 15688 17374 15700
rect 23290 15688 23296 15700
rect 17368 15660 23296 15688
rect 17368 15648 17374 15660
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 23566 15688 23572 15700
rect 23527 15660 23572 15688
rect 23566 15648 23572 15660
rect 23624 15648 23630 15700
rect 31113 15691 31171 15697
rect 31113 15657 31125 15691
rect 31159 15688 31171 15691
rect 36078 15688 36084 15700
rect 31159 15660 36084 15688
rect 31159 15657 31171 15660
rect 31113 15651 31171 15657
rect 36078 15648 36084 15660
rect 36136 15648 36142 15700
rect 19426 15620 19432 15632
rect 16684 15592 19432 15620
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 20806 15580 20812 15632
rect 20864 15620 20870 15632
rect 20864 15592 23060 15620
rect 20864 15580 20870 15592
rect 18230 15552 18236 15564
rect 14844 15524 18236 15552
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14844 15484 14872 15524
rect 18230 15512 18236 15524
rect 18288 15512 18294 15564
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15552 18659 15555
rect 20530 15552 20536 15564
rect 18647 15524 20536 15552
rect 18647 15521 18659 15524
rect 18601 15515 18659 15521
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 20898 15512 20904 15564
rect 20956 15552 20962 15564
rect 21177 15555 21235 15561
rect 21177 15552 21189 15555
rect 20956 15524 21189 15552
rect 20956 15512 20962 15524
rect 21177 15521 21189 15524
rect 21223 15552 21235 15555
rect 22373 15555 22431 15561
rect 22373 15552 22385 15555
rect 21223 15524 22385 15552
rect 21223 15521 21235 15524
rect 21177 15515 21235 15521
rect 22373 15521 22385 15524
rect 22419 15521 22431 15555
rect 23032 15552 23060 15592
rect 23750 15580 23756 15632
rect 23808 15620 23814 15632
rect 25498 15620 25504 15632
rect 23808 15592 25504 15620
rect 23808 15580 23814 15592
rect 25498 15580 25504 15592
rect 25556 15620 25562 15632
rect 25866 15620 25872 15632
rect 25556 15592 25872 15620
rect 25556 15580 25562 15592
rect 25866 15580 25872 15592
rect 25924 15580 25930 15632
rect 25958 15580 25964 15632
rect 26016 15620 26022 15632
rect 27065 15623 27123 15629
rect 27065 15620 27077 15623
rect 26016 15592 27077 15620
rect 26016 15580 26022 15592
rect 27065 15589 27077 15592
rect 27111 15589 27123 15623
rect 27065 15583 27123 15589
rect 28074 15580 28080 15632
rect 28132 15620 28138 15632
rect 28132 15592 31064 15620
rect 28132 15580 28138 15592
rect 24578 15552 24584 15564
rect 23032 15524 24584 15552
rect 22373 15515 22431 15521
rect 24578 15512 24584 15524
rect 24636 15512 24642 15564
rect 25225 15555 25283 15561
rect 25225 15521 25237 15555
rect 25271 15552 25283 15555
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 25271 15524 26433 15552
rect 25271 15521 25283 15524
rect 25225 15515 25283 15521
rect 26421 15521 26433 15524
rect 26467 15552 26479 15555
rect 26467 15524 27844 15552
rect 26467 15521 26479 15524
rect 26421 15515 26479 15521
rect 14323 15456 14872 15484
rect 15657 15487 15715 15493
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 15838 15484 15844 15496
rect 15703 15456 15844 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19518 15484 19524 15496
rect 19392 15456 19524 15484
rect 19392 15444 19398 15456
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 20349 15487 20407 15493
rect 20349 15484 20361 15487
rect 20220 15456 20361 15484
rect 20220 15444 20226 15456
rect 20349 15453 20361 15456
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 24394 15484 24400 15496
rect 23707 15456 24400 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 27816 15484 27844 15524
rect 27890 15512 27896 15564
rect 27948 15552 27954 15564
rect 28445 15555 28503 15561
rect 28445 15552 28457 15555
rect 27948 15524 28457 15552
rect 27948 15512 27954 15524
rect 28445 15521 28457 15524
rect 28491 15552 28503 15555
rect 28626 15552 28632 15564
rect 28491 15524 28632 15552
rect 28491 15521 28503 15524
rect 28445 15515 28503 15521
rect 28626 15512 28632 15524
rect 28684 15512 28690 15564
rect 29086 15552 29092 15564
rect 29047 15524 29092 15552
rect 29086 15512 29092 15524
rect 29144 15512 29150 15564
rect 28258 15484 28264 15496
rect 27816 15456 28264 15484
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 29914 15484 29920 15496
rect 29875 15456 29920 15484
rect 29914 15444 29920 15456
rect 29972 15484 29978 15496
rect 31036 15493 31064 15592
rect 30377 15487 30435 15493
rect 30377 15484 30389 15487
rect 29972 15456 30389 15484
rect 29972 15444 29978 15456
rect 30377 15453 30389 15456
rect 30423 15453 30435 15487
rect 30377 15447 30435 15453
rect 31021 15487 31079 15493
rect 31021 15453 31033 15487
rect 31067 15453 31079 15487
rect 31021 15447 31079 15453
rect 12989 15419 13047 15425
rect 12989 15385 13001 15419
rect 13035 15416 13047 15419
rect 14826 15416 14832 15428
rect 13035 15388 14832 15416
rect 13035 15385 13047 15388
rect 12989 15379 13047 15385
rect 14826 15376 14832 15388
rect 14884 15416 14890 15428
rect 15013 15419 15071 15425
rect 15013 15416 15025 15419
rect 14884 15388 15025 15416
rect 14884 15376 14890 15388
rect 15013 15385 15025 15388
rect 15059 15385 15071 15419
rect 15013 15379 15071 15385
rect 15102 15376 15108 15428
rect 15160 15416 15166 15428
rect 15160 15388 15205 15416
rect 15160 15376 15166 15388
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 16669 15419 16727 15425
rect 16669 15416 16681 15419
rect 15528 15388 16681 15416
rect 15528 15376 15534 15388
rect 16669 15385 16681 15388
rect 16715 15385 16727 15419
rect 17218 15416 17224 15428
rect 17179 15388 17224 15416
rect 16669 15379 16727 15385
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 17310 15376 17316 15428
rect 17368 15416 17374 15428
rect 17957 15419 18015 15425
rect 17957 15416 17969 15419
rect 17368 15388 17413 15416
rect 17880 15388 17969 15416
rect 17368 15376 17374 15388
rect 17880 15360 17908 15388
rect 17957 15385 17969 15388
rect 18003 15385 18015 15419
rect 17957 15379 18015 15385
rect 18049 15419 18107 15425
rect 18049 15385 18061 15419
rect 18095 15416 18107 15419
rect 18138 15416 18144 15428
rect 18095 15388 18144 15416
rect 18095 15385 18107 15388
rect 18049 15379 18107 15385
rect 18138 15376 18144 15388
rect 18196 15376 18202 15428
rect 19242 15376 19248 15428
rect 19300 15416 19306 15428
rect 20257 15419 20315 15425
rect 20257 15416 20269 15419
rect 19300 15388 20269 15416
rect 19300 15376 19306 15388
rect 20257 15385 20269 15388
rect 20303 15385 20315 15419
rect 20257 15379 20315 15385
rect 21266 15376 21272 15428
rect 21324 15416 21330 15428
rect 21821 15419 21879 15425
rect 21324 15388 21369 15416
rect 21324 15376 21330 15388
rect 21821 15385 21833 15419
rect 21867 15385 21879 15419
rect 21821 15379 21879 15385
rect 11701 15351 11759 15357
rect 11701 15317 11713 15351
rect 11747 15348 11759 15351
rect 11974 15348 11980 15360
rect 11747 15320 11980 15348
rect 11747 15317 11759 15320
rect 11701 15311 11759 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 12618 15348 12624 15360
rect 12391 15320 12624 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 14090 15348 14096 15360
rect 13504 15320 14096 15348
rect 13504 15308 13510 15320
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 14369 15351 14427 15357
rect 14369 15317 14381 15351
rect 14415 15348 14427 15351
rect 16022 15348 16028 15360
rect 14415 15320 16028 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 16172 15320 16217 15348
rect 16172 15308 16178 15320
rect 17862 15308 17868 15360
rect 17920 15308 17926 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 20162 15348 20168 15360
rect 19659 15320 20168 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 20346 15308 20352 15360
rect 20404 15348 20410 15360
rect 21836 15348 21864 15379
rect 22370 15376 22376 15428
rect 22428 15416 22434 15428
rect 22465 15419 22523 15425
rect 22465 15416 22477 15419
rect 22428 15388 22477 15416
rect 22428 15376 22434 15388
rect 22465 15385 22477 15388
rect 22511 15385 22523 15419
rect 22465 15379 22523 15385
rect 22830 15376 22836 15428
rect 22888 15416 22894 15428
rect 23017 15419 23075 15425
rect 23017 15416 23029 15419
rect 22888 15388 23029 15416
rect 22888 15376 22894 15388
rect 23017 15385 23029 15388
rect 23063 15416 23075 15419
rect 23474 15416 23480 15428
rect 23063 15388 23480 15416
rect 23063 15385 23075 15388
rect 23017 15379 23075 15385
rect 23474 15376 23480 15388
rect 23532 15376 23538 15428
rect 25130 15416 25136 15428
rect 25091 15388 25136 15416
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 25406 15376 25412 15428
rect 25464 15416 25470 15428
rect 25777 15419 25835 15425
rect 25777 15416 25789 15419
rect 25464 15388 25789 15416
rect 25464 15376 25470 15388
rect 25777 15385 25789 15388
rect 25823 15385 25835 15419
rect 25777 15379 25835 15385
rect 26329 15419 26387 15425
rect 26329 15385 26341 15419
rect 26375 15385 26387 15419
rect 27522 15416 27528 15428
rect 27483 15388 27528 15416
rect 26329 15379 26387 15385
rect 24670 15348 24676 15360
rect 20404 15320 24676 15348
rect 20404 15308 20410 15320
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 24854 15308 24860 15360
rect 24912 15348 24918 15360
rect 26344 15348 26372 15379
rect 27522 15376 27528 15388
rect 27580 15376 27586 15428
rect 27617 15419 27675 15425
rect 27617 15385 27629 15419
rect 27663 15416 27675 15419
rect 27798 15416 27804 15428
rect 27663 15388 27804 15416
rect 27663 15385 27675 15388
rect 27617 15379 27675 15385
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 28534 15376 28540 15428
rect 28592 15416 28598 15428
rect 28592 15388 28637 15416
rect 28592 15376 28598 15388
rect 24912 15320 26372 15348
rect 27816 15348 27844 15376
rect 29270 15348 29276 15360
rect 27816 15320 29276 15348
rect 24912 15308 24918 15320
rect 29270 15308 29276 15320
rect 29328 15308 29334 15360
rect 29822 15348 29828 15360
rect 29783 15320 29828 15348
rect 29822 15308 29828 15320
rect 29880 15308 29886 15360
rect 30466 15348 30472 15360
rect 30427 15320 30472 15348
rect 30466 15308 30472 15320
rect 30524 15308 30530 15360
rect 1104 15258 36892 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 36892 15258
rect 1104 15184 36892 15206
rect 2590 15104 2596 15156
rect 2648 15144 2654 15156
rect 17126 15144 17132 15156
rect 2648 15116 17132 15144
rect 2648 15104 2654 15116
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 17221 15147 17279 15153
rect 17221 15113 17233 15147
rect 17267 15144 17279 15147
rect 18046 15144 18052 15156
rect 17267 15116 18052 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 20898 15144 20904 15156
rect 20272 15116 20904 15144
rect 7558 15036 7564 15088
rect 7616 15076 7622 15088
rect 9950 15076 9956 15088
rect 7616 15048 9956 15076
rect 7616 15036 7622 15048
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 11146 15076 11152 15088
rect 11107 15048 11152 15076
rect 11146 15036 11152 15048
rect 11204 15036 11210 15088
rect 13541 15079 13599 15085
rect 13541 15045 13553 15079
rect 13587 15076 13599 15079
rect 13814 15076 13820 15088
rect 13587 15048 13820 15076
rect 13587 15045 13599 15048
rect 13541 15039 13599 15045
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 14366 15076 14372 15088
rect 14327 15048 14372 15076
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 16209 15079 16267 15085
rect 16209 15045 16221 15079
rect 16255 15076 16267 15079
rect 17957 15079 18015 15085
rect 17957 15076 17969 15079
rect 16255 15048 17969 15076
rect 16255 15045 16267 15048
rect 16209 15039 16267 15045
rect 17957 15045 17969 15048
rect 18003 15045 18015 15079
rect 17957 15039 18015 15045
rect 18230 15036 18236 15088
rect 18288 15076 18294 15088
rect 18288 15048 18736 15076
rect 18288 15036 18294 15048
rect 18708 15020 18736 15048
rect 20070 15036 20076 15088
rect 20128 15076 20134 15088
rect 20272 15085 20300 15116
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 22462 15104 22468 15156
rect 22520 15144 22526 15156
rect 22520 15116 24624 15144
rect 22520 15104 22526 15116
rect 20165 15079 20223 15085
rect 20165 15076 20177 15079
rect 20128 15048 20177 15076
rect 20128 15036 20134 15048
rect 20165 15045 20177 15048
rect 20211 15045 20223 15079
rect 20165 15039 20223 15045
rect 20257 15079 20315 15085
rect 20257 15045 20269 15079
rect 20303 15045 20315 15079
rect 20257 15039 20315 15045
rect 20530 15036 20536 15088
rect 20588 15076 20594 15088
rect 22554 15076 22560 15088
rect 20588 15048 21128 15076
rect 22515 15048 22560 15076
rect 20588 15036 20594 15048
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 11790 15008 11796 15020
rect 10643 14980 11796 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 11790 14968 11796 14980
rect 11848 15008 11854 15020
rect 11977 15011 12035 15017
rect 11977 15008 11989 15011
rect 11848 14980 11989 15008
rect 11848 14968 11854 14980
rect 11977 14977 11989 14980
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15436 14980 16129 15008
rect 15436 14968 15442 14980
rect 16117 14977 16129 14980
rect 16163 15008 16175 15011
rect 16390 15008 16396 15020
rect 16163 14980 16396 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17218 15008 17224 15020
rect 17175 14980 17224 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 18690 14968 18696 15020
rect 18748 15008 18754 15020
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 18748 14980 19165 15008
rect 18748 14968 18754 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 13357 14943 13415 14949
rect 13357 14940 13369 14943
rect 8168 14912 13369 14940
rect 8168 14900 8174 14912
rect 13357 14909 13369 14912
rect 13403 14940 13415 14943
rect 13538 14940 13544 14952
rect 13403 14912 13544 14940
rect 13403 14909 13415 14912
rect 13357 14903 13415 14909
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13998 14940 14004 14952
rect 13679 14912 14004 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14090 14900 14096 14952
rect 14148 14940 14154 14952
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 14148 14912 14289 14940
rect 14148 14900 14154 14912
rect 14277 14909 14289 14912
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14516 14912 15117 14940
rect 14516 14900 14522 14912
rect 15105 14909 15117 14912
rect 15151 14940 15163 14943
rect 17862 14940 17868 14952
rect 15151 14912 16896 14940
rect 17823 14912 17868 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 8294 14832 8300 14884
rect 8352 14872 8358 14884
rect 16758 14872 16764 14884
rect 8352 14844 16764 14872
rect 8352 14832 8358 14844
rect 16758 14832 16764 14844
rect 16816 14832 16822 14884
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 13630 14804 13636 14816
rect 12115 14776 13636 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 16868 14804 16896 14912
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 21008 14940 21036 14971
rect 17972 14912 21036 14940
rect 21100 14940 21128 15048
rect 22554 15036 22560 15048
rect 22612 15036 22618 15088
rect 22646 15036 22652 15088
rect 22704 15076 22710 15088
rect 23385 15079 23443 15085
rect 23385 15076 23397 15079
rect 22704 15048 23397 15076
rect 22704 15036 22710 15048
rect 23385 15045 23397 15048
rect 23431 15045 23443 15079
rect 23385 15039 23443 15045
rect 24302 15036 24308 15088
rect 24360 15076 24366 15088
rect 24596 15085 24624 15116
rect 24670 15104 24676 15156
rect 24728 15144 24734 15156
rect 26878 15144 26884 15156
rect 24728 15116 26884 15144
rect 24728 15104 24734 15116
rect 26878 15104 26884 15116
rect 26936 15104 26942 15156
rect 28626 15144 28632 15156
rect 28587 15116 28632 15144
rect 28626 15104 28632 15116
rect 28684 15104 28690 15156
rect 29086 15104 29092 15156
rect 29144 15104 29150 15156
rect 35986 15144 35992 15156
rect 35947 15116 35992 15144
rect 35986 15104 35992 15116
rect 36044 15104 36050 15156
rect 36170 15104 36176 15156
rect 36228 15104 36234 15156
rect 24489 15079 24547 15085
rect 24489 15076 24501 15079
rect 24360 15048 24501 15076
rect 24360 15036 24366 15048
rect 24489 15045 24501 15048
rect 24535 15045 24547 15079
rect 24489 15039 24547 15045
rect 24581 15079 24639 15085
rect 24581 15045 24593 15079
rect 24627 15045 24639 15079
rect 25774 15076 25780 15088
rect 25735 15048 25780 15076
rect 24581 15039 24639 15045
rect 25774 15036 25780 15048
rect 25832 15036 25838 15088
rect 27614 15076 27620 15088
rect 27575 15048 27620 15076
rect 27614 15036 27620 15048
rect 27672 15036 27678 15088
rect 28169 15079 28227 15085
rect 28169 15045 28181 15079
rect 28215 15076 28227 15079
rect 29104 15076 29132 15104
rect 28215 15048 29132 15076
rect 30653 15079 30711 15085
rect 28215 15045 28227 15048
rect 28169 15039 28227 15045
rect 30653 15045 30665 15079
rect 30699 15076 30711 15079
rect 36188 15076 36216 15104
rect 30699 15048 36216 15076
rect 30699 15045 30711 15048
rect 30653 15039 30711 15045
rect 29089 15011 29147 15017
rect 29089 14977 29101 15011
rect 29135 15008 29147 15011
rect 29822 15008 29828 15020
rect 29135 14980 29828 15008
rect 29135 14977 29147 14980
rect 29089 14971 29147 14977
rect 29822 14968 29828 14980
rect 29880 14968 29886 15020
rect 31205 15011 31263 15017
rect 31205 15008 31217 15011
rect 29932 14980 31217 15008
rect 22370 14940 22376 14952
rect 21100 14912 22376 14940
rect 17126 14832 17132 14884
rect 17184 14872 17190 14884
rect 17972 14872 18000 14912
rect 17184 14844 18000 14872
rect 18417 14875 18475 14881
rect 17184 14832 17190 14844
rect 18417 14841 18429 14875
rect 18463 14872 18475 14875
rect 18463 14844 19656 14872
rect 18463 14841 18475 14844
rect 18417 14835 18475 14841
rect 17954 14804 17960 14816
rect 16868 14776 17960 14804
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 18380 14776 19073 14804
rect 18380 14764 18386 14776
rect 19061 14773 19073 14776
rect 19107 14773 19119 14807
rect 19628 14804 19656 14844
rect 19702 14832 19708 14884
rect 19760 14872 19766 14884
rect 20530 14872 20536 14884
rect 19760 14844 20536 14872
rect 19760 14832 19766 14844
rect 20530 14832 20536 14844
rect 20588 14832 20594 14884
rect 20714 14804 20720 14816
rect 19628 14776 20720 14804
rect 19061 14767 19119 14773
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 20916 14804 20944 14912
rect 22370 14900 22376 14912
rect 22428 14900 22434 14952
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14909 22707 14943
rect 23290 14940 23296 14952
rect 23251 14912 23296 14940
rect 22649 14903 22707 14909
rect 22097 14875 22155 14881
rect 22097 14841 22109 14875
rect 22143 14872 22155 14875
rect 22186 14872 22192 14884
rect 22143 14844 22192 14872
rect 22143 14841 22155 14844
rect 22097 14835 22155 14841
rect 22186 14832 22192 14844
rect 22244 14832 22250 14884
rect 22664 14872 22692 14903
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23934 14940 23940 14952
rect 23895 14912 23940 14940
rect 23934 14900 23940 14912
rect 23992 14900 23998 14952
rect 24578 14900 24584 14952
rect 24636 14940 24642 14952
rect 24765 14943 24823 14949
rect 24765 14940 24777 14943
rect 24636 14912 24777 14940
rect 24636 14900 24642 14912
rect 24765 14909 24777 14912
rect 24811 14909 24823 14943
rect 25682 14940 25688 14952
rect 25643 14912 25688 14940
rect 24765 14903 24823 14909
rect 25682 14900 25688 14912
rect 25740 14900 25746 14952
rect 26326 14940 26332 14952
rect 26239 14912 26332 14940
rect 26326 14900 26332 14912
rect 26384 14940 26390 14952
rect 27338 14940 27344 14952
rect 26384 14912 27344 14940
rect 26384 14900 26390 14912
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 27525 14943 27583 14949
rect 27525 14909 27537 14943
rect 27571 14909 27583 14943
rect 27525 14903 27583 14909
rect 22664 14844 23152 14872
rect 22922 14804 22928 14816
rect 20916 14776 22928 14804
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 23124 14804 23152 14844
rect 23198 14832 23204 14884
rect 23256 14872 23262 14884
rect 26418 14872 26424 14884
rect 23256 14844 26424 14872
rect 23256 14832 23262 14844
rect 26418 14832 26424 14844
rect 26476 14872 26482 14884
rect 27540 14872 27568 14903
rect 27706 14900 27712 14952
rect 27764 14940 27770 14952
rect 28994 14940 29000 14952
rect 27764 14912 29000 14940
rect 27764 14900 27770 14912
rect 28994 14900 29000 14912
rect 29052 14900 29058 14952
rect 29270 14940 29276 14952
rect 29231 14912 29276 14940
rect 29270 14900 29276 14912
rect 29328 14900 29334 14952
rect 29932 14940 29960 14980
rect 31205 14977 31217 14980
rect 31251 14977 31263 15011
rect 31205 14971 31263 14977
rect 36081 15011 36139 15017
rect 36081 14977 36093 15011
rect 36127 15008 36139 15011
rect 36170 15008 36176 15020
rect 36127 14980 36176 15008
rect 36127 14977 36139 14980
rect 36081 14971 36139 14977
rect 29380 14912 29960 14940
rect 29380 14872 29408 14912
rect 31110 14872 31116 14884
rect 26476 14844 27568 14872
rect 27632 14844 29408 14872
rect 29748 14844 31116 14872
rect 26476 14832 26482 14844
rect 26786 14804 26792 14816
rect 23124 14776 26792 14804
rect 26786 14764 26792 14776
rect 26844 14804 26850 14816
rect 27632 14804 27660 14844
rect 26844 14776 27660 14804
rect 26844 14764 26850 14776
rect 28166 14764 28172 14816
rect 28224 14804 28230 14816
rect 29748 14813 29776 14844
rect 31110 14832 31116 14844
rect 31168 14832 31174 14884
rect 29733 14807 29791 14813
rect 29733 14804 29745 14807
rect 28224 14776 29745 14804
rect 28224 14764 28230 14776
rect 29733 14773 29745 14776
rect 29779 14773 29791 14807
rect 29733 14767 29791 14773
rect 30006 14764 30012 14816
rect 30064 14804 30070 14816
rect 30377 14807 30435 14813
rect 30377 14804 30389 14807
rect 30064 14776 30389 14804
rect 30064 14764 30070 14776
rect 30377 14773 30389 14776
rect 30423 14773 30435 14807
rect 31220 14804 31248 14971
rect 36170 14968 36176 14980
rect 36228 14968 36234 15020
rect 31754 14804 31760 14816
rect 31220 14776 31760 14804
rect 30377 14767 30435 14773
rect 31754 14764 31760 14776
rect 31812 14764 31818 14816
rect 1104 14714 36892 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36892 14714
rect 1104 14640 36892 14662
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 14366 14600 14372 14612
rect 11296 14572 14372 14600
rect 11296 14560 11302 14572
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 20806 14600 20812 14612
rect 14792 14572 20812 14600
rect 14792 14560 14798 14572
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 21266 14600 21272 14612
rect 21227 14572 21272 14600
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 21542 14600 21548 14612
rect 21416 14572 21548 14600
rect 21416 14560 21422 14572
rect 21542 14560 21548 14572
rect 21600 14600 21606 14612
rect 23842 14600 23848 14612
rect 21600 14572 23848 14600
rect 21600 14560 21606 14572
rect 23842 14560 23848 14572
rect 23900 14560 23906 14612
rect 23937 14603 23995 14609
rect 23937 14569 23949 14603
rect 23983 14600 23995 14603
rect 25774 14600 25780 14612
rect 23983 14572 25780 14600
rect 23983 14569 23995 14572
rect 23937 14563 23995 14569
rect 25774 14560 25780 14572
rect 25832 14560 25838 14612
rect 26786 14560 26792 14612
rect 26844 14560 26850 14612
rect 28258 14560 28264 14612
rect 28316 14600 28322 14612
rect 29825 14603 29883 14609
rect 29825 14600 29837 14603
rect 28316 14572 29837 14600
rect 28316 14560 28322 14572
rect 29825 14569 29837 14572
rect 29871 14569 29883 14603
rect 29825 14563 29883 14569
rect 10597 14535 10655 14541
rect 10597 14501 10609 14535
rect 10643 14532 10655 14535
rect 13633 14535 13691 14541
rect 10643 14504 13584 14532
rect 10643 14501 10655 14504
rect 10597 14495 10655 14501
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 11330 14464 11336 14476
rect 10091 14436 11336 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14464 11851 14467
rect 12894 14464 12900 14476
rect 11839 14436 12900 14464
rect 11839 14433 11851 14436
rect 11793 14427 11851 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13556 14464 13584 14504
rect 13633 14501 13645 14535
rect 13679 14532 13691 14535
rect 13998 14532 14004 14544
rect 13679 14504 14004 14532
rect 13679 14501 13691 14504
rect 13633 14495 13691 14501
rect 13998 14492 14004 14504
rect 14056 14532 14062 14544
rect 15470 14532 15476 14544
rect 14056 14504 15476 14532
rect 14056 14492 14062 14504
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 16025 14535 16083 14541
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 17221 14535 17279 14541
rect 17221 14532 17233 14535
rect 16071 14504 17233 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 17221 14501 17233 14504
rect 17267 14532 17279 14535
rect 26234 14532 26240 14544
rect 17267 14504 26240 14532
rect 17267 14501 17279 14504
rect 17221 14495 17279 14501
rect 26234 14492 26240 14504
rect 26292 14492 26298 14544
rect 13556 14436 14780 14464
rect 14752 14408 14780 14436
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 17678 14464 17684 14476
rect 16816 14436 17684 14464
rect 16816 14424 16822 14436
rect 17678 14424 17684 14436
rect 17736 14424 17742 14476
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 17828 14436 18245 14464
rect 17828 14424 17834 14436
rect 18233 14433 18245 14436
rect 18279 14464 18291 14467
rect 18414 14464 18420 14476
rect 18279 14436 18420 14464
rect 18279 14433 18291 14436
rect 18233 14427 18291 14433
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 18877 14467 18935 14473
rect 18877 14433 18889 14467
rect 18923 14464 18935 14467
rect 23198 14464 23204 14476
rect 18923 14436 23204 14464
rect 18923 14433 18935 14436
rect 18877 14427 18935 14433
rect 23198 14424 23204 14436
rect 23256 14424 23262 14476
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 23658 14464 23664 14476
rect 23431 14436 23664 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 23658 14424 23664 14436
rect 23716 14424 23722 14476
rect 26804 14473 26832 14560
rect 26789 14467 26847 14473
rect 26789 14433 26801 14467
rect 26835 14433 26847 14467
rect 26789 14427 26847 14433
rect 27062 14424 27068 14476
rect 27120 14464 27126 14476
rect 30466 14464 30472 14476
rect 27120 14436 30472 14464
rect 27120 14424 27126 14436
rect 30466 14424 30472 14436
rect 30524 14424 30530 14476
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 10008 14368 11253 14396
rect 10008 14356 10014 14368
rect 11241 14365 11253 14368
rect 11287 14365 11299 14399
rect 11698 14396 11704 14408
rect 11659 14368 11704 14396
rect 11241 14359 11299 14365
rect 11256 14328 11284 14359
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12342 14396 12348 14408
rect 12303 14368 12348 14396
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 14734 14396 14740 14408
rect 14695 14368 14740 14396
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 21174 14356 21180 14408
rect 21232 14396 21238 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 21232 14368 21373 14396
rect 21232 14356 21238 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 12526 14328 12532 14340
rect 11256 14300 12532 14328
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 12710 14288 12716 14340
rect 12768 14328 12774 14340
rect 13081 14331 13139 14337
rect 13081 14328 13093 14331
rect 12768 14300 13093 14328
rect 12768 14288 12774 14300
rect 13081 14297 13093 14300
rect 13127 14297 13139 14331
rect 13081 14291 13139 14297
rect 13173 14331 13231 14337
rect 13173 14297 13185 14331
rect 13219 14297 13231 14331
rect 15470 14328 15476 14340
rect 15431 14300 15476 14328
rect 13173 14291 13231 14297
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 11112 14232 11161 14260
rect 11112 14220 11118 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 12342 14260 12348 14272
rect 11388 14232 12348 14260
rect 11388 14220 11394 14232
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 12437 14263 12495 14269
rect 12437 14229 12449 14263
rect 12483 14260 12495 14263
rect 13188 14260 13216 14291
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 15565 14331 15623 14337
rect 15565 14297 15577 14331
rect 15611 14297 15623 14331
rect 16666 14328 16672 14340
rect 16627 14300 16672 14328
rect 15565 14291 15623 14297
rect 12483 14232 13216 14260
rect 14829 14263 14887 14269
rect 12483 14229 12495 14232
rect 12437 14223 12495 14229
rect 14829 14229 14841 14263
rect 14875 14260 14887 14263
rect 15580 14260 15608 14291
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 16761 14331 16819 14337
rect 16761 14297 16773 14331
rect 16807 14297 16819 14331
rect 16761 14291 16819 14297
rect 14875 14232 15608 14260
rect 14875 14229 14887 14232
rect 14829 14223 14887 14229
rect 16022 14220 16028 14272
rect 16080 14260 16086 14272
rect 16776 14260 16804 14291
rect 18322 14288 18328 14340
rect 18380 14328 18386 14340
rect 19981 14331 20039 14337
rect 18380 14300 18425 14328
rect 18380 14288 18386 14300
rect 19981 14297 19993 14331
rect 20027 14328 20039 14331
rect 20027 14300 20116 14328
rect 20027 14297 20039 14300
rect 19981 14291 20039 14297
rect 20088 14272 20116 14300
rect 20162 14288 20168 14340
rect 20220 14328 20226 14340
rect 20533 14331 20591 14337
rect 20533 14328 20545 14331
rect 20220 14300 20545 14328
rect 20220 14288 20226 14300
rect 20533 14297 20545 14300
rect 20579 14297 20591 14331
rect 20533 14291 20591 14297
rect 20625 14331 20683 14337
rect 20625 14297 20637 14331
rect 20671 14328 20683 14331
rect 21082 14328 21088 14340
rect 20671 14300 21088 14328
rect 20671 14297 20683 14300
rect 20625 14291 20683 14297
rect 21082 14288 21088 14300
rect 21140 14288 21146 14340
rect 22370 14328 22376 14340
rect 22331 14300 22376 14328
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 22465 14331 22523 14337
rect 22465 14297 22477 14331
rect 22511 14297 22523 14331
rect 23676 14328 23704 14424
rect 23842 14396 23848 14408
rect 23803 14368 23848 14396
rect 23842 14356 23848 14368
rect 23900 14356 23906 14408
rect 28074 14356 28080 14408
rect 28132 14396 28138 14408
rect 28132 14368 28177 14396
rect 28132 14356 28138 14368
rect 28350 14356 28356 14408
rect 28408 14396 28414 14408
rect 28537 14399 28595 14405
rect 28537 14396 28549 14399
rect 28408 14368 28549 14396
rect 28408 14356 28414 14368
rect 28537 14365 28549 14368
rect 28583 14365 28595 14399
rect 28537 14359 28595 14365
rect 28994 14356 29000 14408
rect 29052 14396 29058 14408
rect 29917 14399 29975 14405
rect 29917 14396 29929 14399
rect 29052 14368 29929 14396
rect 29052 14356 29058 14368
rect 29917 14365 29929 14368
rect 29963 14396 29975 14399
rect 30377 14399 30435 14405
rect 29963 14368 30328 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 24581 14331 24639 14337
rect 24581 14328 24593 14331
rect 23676 14300 24593 14328
rect 22465 14291 22523 14297
rect 24581 14297 24593 14300
rect 24627 14297 24639 14331
rect 24581 14291 24639 14297
rect 25501 14331 25559 14337
rect 25501 14297 25513 14331
rect 25547 14297 25559 14331
rect 25501 14291 25559 14297
rect 16080 14232 16804 14260
rect 16080 14220 16086 14232
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 19392 14232 19441 14260
rect 19392 14220 19398 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 20070 14220 20076 14272
rect 20128 14220 20134 14272
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21910 14260 21916 14272
rect 20772 14232 21916 14260
rect 20772 14220 20778 14232
rect 21910 14220 21916 14232
rect 21968 14220 21974 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22094 14260 22100 14272
rect 22060 14232 22100 14260
rect 22060 14220 22066 14232
rect 22094 14220 22100 14232
rect 22152 14220 22158 14272
rect 22480 14260 22508 14291
rect 25314 14260 25320 14272
rect 22480 14232 25320 14260
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 25516 14260 25544 14291
rect 25590 14288 25596 14340
rect 25648 14328 25654 14340
rect 26697 14331 26755 14337
rect 25648 14300 25693 14328
rect 25648 14288 25654 14300
rect 26697 14297 26709 14331
rect 26743 14328 26755 14331
rect 26970 14328 26976 14340
rect 26743 14300 26976 14328
rect 26743 14297 26755 14300
rect 26697 14291 26755 14297
rect 26970 14288 26976 14300
rect 27028 14288 27034 14340
rect 27246 14288 27252 14340
rect 27304 14328 27310 14340
rect 27433 14331 27491 14337
rect 27433 14328 27445 14331
rect 27304 14300 27445 14328
rect 27304 14288 27310 14300
rect 27433 14297 27445 14300
rect 27479 14297 27491 14331
rect 27433 14291 27491 14297
rect 27525 14331 27583 14337
rect 27525 14297 27537 14331
rect 27571 14328 27583 14331
rect 30098 14328 30104 14340
rect 27571 14300 30104 14328
rect 27571 14297 27583 14300
rect 27525 14291 27583 14297
rect 30098 14288 30104 14300
rect 30156 14288 30162 14340
rect 30300 14328 30328 14368
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30558 14396 30564 14408
rect 30423 14368 30564 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 30558 14356 30564 14368
rect 30616 14356 30622 14408
rect 31113 14399 31171 14405
rect 31113 14365 31125 14399
rect 31159 14396 31171 14399
rect 31754 14396 31760 14408
rect 31159 14368 31760 14396
rect 31159 14365 31171 14368
rect 31113 14359 31171 14365
rect 31754 14356 31760 14368
rect 31812 14356 31818 14408
rect 31573 14331 31631 14337
rect 31573 14328 31585 14331
rect 30300 14300 31585 14328
rect 31128 14272 31156 14300
rect 31573 14297 31585 14300
rect 31619 14297 31631 14331
rect 31573 14291 31631 14297
rect 28629 14263 28687 14269
rect 28629 14260 28641 14263
rect 25516 14232 28641 14260
rect 28629 14229 28641 14232
rect 28675 14229 28687 14263
rect 30466 14260 30472 14272
rect 30427 14232 30472 14260
rect 28629 14223 28687 14229
rect 30466 14220 30472 14232
rect 30524 14220 30530 14272
rect 31110 14220 31116 14272
rect 31168 14220 31174 14272
rect 1104 14170 36892 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 36892 14170
rect 1104 14096 36892 14118
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 13446 14056 13452 14068
rect 11103 14028 13452 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 13955 14028 15700 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 12618 13988 12624 14000
rect 12579 13960 12624 13988
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 13173 13991 13231 13997
rect 13173 13957 13185 13991
rect 13219 13988 13231 13991
rect 13998 13988 14004 14000
rect 13219 13960 14004 13988
rect 13219 13957 13231 13960
rect 13173 13951 13231 13957
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 15672 13997 15700 14028
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 20070 14056 20076 14068
rect 16448 14028 20076 14056
rect 16448 14016 16454 14028
rect 14553 13991 14611 13997
rect 14553 13957 14565 13991
rect 14599 13988 14611 13991
rect 15657 13991 15715 13997
rect 14599 13960 15516 13988
rect 14599 13957 14611 13960
rect 14553 13951 14611 13957
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 9122 13920 9128 13932
rect 8619 13892 9128 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 9122 13880 9128 13892
rect 9180 13920 9186 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 9180 13892 10149 13920
rect 9180 13880 9186 13892
rect 10137 13889 10149 13892
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11606 13920 11612 13932
rect 11195 13892 11612 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11756 13892 11805 13920
rect 11756 13880 11762 13892
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 14090 13920 14096 13932
rect 11793 13883 11851 13889
rect 13188 13892 14096 13920
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13852 10287 13855
rect 11514 13852 11520 13864
rect 10275 13824 11520 13852
rect 10275 13821 10287 13824
rect 10229 13815 10287 13821
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12342 13852 12348 13864
rect 11931 13824 12348 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12529 13855 12587 13861
rect 12529 13852 12541 13855
rect 12452 13824 12541 13852
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 10962 13784 10968 13796
rect 9723 13756 10968 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 11054 13744 11060 13796
rect 11112 13784 11118 13796
rect 12452 13784 12480 13824
rect 12529 13821 12541 13824
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 13188 13852 13216 13892
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 12676 13824 13216 13852
rect 12676 13812 12682 13824
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 13688 13824 14473 13852
rect 13688 13812 13694 13824
rect 14461 13821 14473 13824
rect 14507 13821 14519 13855
rect 15488 13852 15516 13960
rect 15657 13957 15669 13991
rect 15703 13957 15715 13991
rect 15657 13951 15715 13957
rect 15746 13948 15752 14000
rect 15804 13988 15810 14000
rect 17328 13997 17356 14028
rect 20070 14016 20076 14028
rect 20128 14056 20134 14068
rect 22002 14056 22008 14068
rect 20128 14028 22008 14056
rect 20128 14016 20134 14028
rect 22002 14016 22008 14028
rect 22060 14016 22066 14068
rect 22097 14059 22155 14065
rect 22097 14025 22109 14059
rect 22143 14056 22155 14059
rect 22554 14056 22560 14068
rect 22143 14028 22560 14056
rect 22143 14025 22155 14028
rect 22097 14019 22155 14025
rect 22554 14016 22560 14028
rect 22612 14016 22618 14068
rect 22646 14016 22652 14068
rect 22704 14016 22710 14068
rect 22741 14059 22799 14065
rect 22741 14025 22753 14059
rect 22787 14056 22799 14059
rect 23382 14056 23388 14068
rect 22787 14028 23388 14056
rect 22787 14025 22799 14028
rect 22741 14019 22799 14025
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 25222 14016 25228 14068
rect 25280 14056 25286 14068
rect 26237 14059 26295 14065
rect 26237 14056 26249 14059
rect 25280 14028 26249 14056
rect 25280 14016 25286 14028
rect 26237 14025 26249 14028
rect 26283 14025 26295 14059
rect 30466 14056 30472 14068
rect 26237 14019 26295 14025
rect 27356 14028 30472 14056
rect 17313 13991 17371 13997
rect 15804 13960 15849 13988
rect 15804 13948 15810 13960
rect 17313 13957 17325 13991
rect 17359 13957 17371 13991
rect 17313 13951 17371 13957
rect 17402 13948 17408 14000
rect 17460 13988 17466 14000
rect 17460 13960 17505 13988
rect 17460 13948 17466 13960
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 18230 13988 18236 14000
rect 17736 13960 18236 13988
rect 17736 13948 17742 13960
rect 18230 13948 18236 13960
rect 18288 13988 18294 14000
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 18288 13960 18337 13988
rect 18288 13948 18294 13960
rect 18325 13957 18337 13960
rect 18371 13957 18383 13991
rect 18966 13988 18972 14000
rect 18927 13960 18972 13988
rect 18325 13951 18383 13957
rect 18966 13948 18972 13960
rect 19024 13948 19030 14000
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 19981 13991 20039 13997
rect 19981 13988 19993 13991
rect 19116 13960 19993 13988
rect 19116 13948 19122 13960
rect 19981 13957 19993 13960
rect 20027 13957 20039 13991
rect 20530 13988 20536 14000
rect 20491 13960 20536 13988
rect 19981 13951 20039 13957
rect 20530 13948 20536 13960
rect 20588 13948 20594 14000
rect 21361 13991 21419 13997
rect 21361 13957 21373 13991
rect 21407 13988 21419 13991
rect 22664 13988 22692 14016
rect 21407 13960 22692 13988
rect 21407 13957 21419 13960
rect 21361 13951 21419 13957
rect 23566 13948 23572 14000
rect 23624 13988 23630 14000
rect 25501 13991 25559 13997
rect 23624 13960 23669 13988
rect 23624 13948 23630 13960
rect 25501 13957 25513 13991
rect 25547 13988 25559 13991
rect 26418 13988 26424 14000
rect 25547 13960 26424 13988
rect 25547 13957 25559 13960
rect 25501 13951 25559 13957
rect 26418 13948 26424 13960
rect 26476 13948 26482 14000
rect 26878 13948 26884 14000
rect 26936 13988 26942 14000
rect 27356 13997 27384 14028
rect 30466 14016 30472 14028
rect 30524 14016 30530 14068
rect 35986 14016 35992 14068
rect 36044 14056 36050 14068
rect 36173 14059 36231 14065
rect 36173 14056 36185 14059
rect 36044 14028 36185 14056
rect 36044 14016 36050 14028
rect 36173 14025 36185 14028
rect 36219 14025 36231 14059
rect 36173 14019 36231 14025
rect 27249 13991 27307 13997
rect 27249 13988 27261 13991
rect 26936 13960 27261 13988
rect 26936 13948 26942 13960
rect 27249 13957 27261 13960
rect 27295 13957 27307 13991
rect 27249 13951 27307 13957
rect 27341 13991 27399 13997
rect 27341 13957 27353 13991
rect 27387 13957 27399 13991
rect 27341 13951 27399 13957
rect 27890 13948 27896 14000
rect 27948 13988 27954 14000
rect 28537 13991 28595 13997
rect 28537 13988 28549 13991
rect 27948 13960 28549 13988
rect 27948 13948 27954 13960
rect 28537 13957 28549 13960
rect 28583 13957 28595 13991
rect 29086 13988 29092 14000
rect 29047 13960 29092 13988
rect 28537 13951 28595 13957
rect 29086 13948 29092 13960
rect 29144 13948 29150 14000
rect 29196 13960 29868 13988
rect 21174 13880 21180 13932
rect 21232 13920 21238 13932
rect 21269 13923 21327 13929
rect 21269 13920 21281 13923
rect 21232 13892 21281 13920
rect 21232 13880 21238 13892
rect 21269 13889 21281 13892
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 22094 13880 22100 13932
rect 22152 13920 22158 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 22152 13892 22201 13920
rect 22152 13880 22158 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22646 13920 22652 13932
rect 22607 13892 22652 13920
rect 22189 13883 22247 13889
rect 22646 13880 22652 13892
rect 22704 13880 22710 13932
rect 26329 13923 26387 13929
rect 24320 13892 24532 13920
rect 16758 13852 16764 13864
rect 15488 13824 16764 13852
rect 14461 13815 14519 13821
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 18414 13812 18420 13864
rect 18472 13852 18478 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18472 13824 18889 13852
rect 18472 13812 18478 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 19518 13852 19524 13864
rect 19431 13824 19524 13852
rect 18877 13815 18935 13821
rect 19518 13812 19524 13824
rect 19576 13852 19582 13864
rect 19576 13824 20208 13852
rect 19576 13812 19582 13824
rect 11112 13756 12480 13784
rect 11112 13744 11118 13756
rect 14366 13744 14372 13796
rect 14424 13784 14430 13796
rect 15010 13784 15016 13796
rect 14424 13756 15016 13784
rect 14424 13744 14430 13756
rect 15010 13744 15016 13756
rect 15068 13744 15074 13796
rect 16209 13787 16267 13793
rect 16209 13753 16221 13787
rect 16255 13784 16267 13787
rect 17954 13784 17960 13796
rect 16255 13756 17960 13784
rect 16255 13753 16267 13756
rect 16209 13747 16267 13753
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 19794 13784 19800 13796
rect 18288 13756 19800 13784
rect 18288 13744 18294 13756
rect 19794 13744 19800 13756
rect 19852 13784 19858 13796
rect 20070 13784 20076 13796
rect 19852 13756 20076 13784
rect 19852 13744 19858 13756
rect 20070 13744 20076 13756
rect 20128 13744 20134 13796
rect 20180 13784 20208 13824
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20312 13824 20637 13852
rect 20312 13812 20318 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 21726 13812 21732 13864
rect 21784 13852 21790 13864
rect 23477 13855 23535 13861
rect 23477 13852 23489 13855
rect 21784 13824 23489 13852
rect 21784 13812 21790 13824
rect 23477 13821 23489 13824
rect 23523 13852 23535 13855
rect 23658 13852 23664 13864
rect 23523 13824 23664 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 24320 13784 24348 13892
rect 24397 13855 24455 13861
rect 24397 13821 24409 13855
rect 24443 13821 24455 13855
rect 24504 13852 24532 13892
rect 26329 13889 26341 13923
rect 26375 13920 26387 13923
rect 26970 13920 26976 13932
rect 26375 13892 26976 13920
rect 26375 13889 26387 13892
rect 26329 13883 26387 13889
rect 26970 13880 26976 13892
rect 27028 13880 27034 13932
rect 25317 13855 25375 13861
rect 25317 13852 25329 13855
rect 24504 13824 25329 13852
rect 24397 13815 24455 13821
rect 25317 13821 25329 13824
rect 25363 13852 25375 13855
rect 25406 13852 25412 13864
rect 25363 13824 25412 13852
rect 25363 13821 25375 13824
rect 25317 13815 25375 13821
rect 20180 13756 24348 13784
rect 1670 13716 1676 13728
rect 1631 13688 1676 13716
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 12342 13716 12348 13728
rect 10744 13688 12348 13716
rect 10744 13676 10750 13688
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 17034 13716 17040 13728
rect 13044 13688 17040 13716
rect 13044 13676 13050 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 24412 13716 24440 13815
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25593 13855 25651 13861
rect 25593 13821 25605 13855
rect 25639 13852 25651 13855
rect 25958 13852 25964 13864
rect 25639 13824 25964 13852
rect 25639 13821 25651 13824
rect 25593 13815 25651 13821
rect 25958 13812 25964 13824
rect 26016 13812 26022 13864
rect 27893 13855 27951 13861
rect 27356 13824 27844 13852
rect 24946 13744 24952 13796
rect 25004 13784 25010 13796
rect 27356 13784 27384 13824
rect 25004 13756 27384 13784
rect 27816 13784 27844 13824
rect 27893 13821 27905 13855
rect 27939 13852 27951 13855
rect 28074 13852 28080 13864
rect 27939 13824 28080 13852
rect 27939 13821 27951 13824
rect 27893 13815 27951 13821
rect 28074 13812 28080 13824
rect 28132 13812 28138 13864
rect 28442 13852 28448 13864
rect 28403 13824 28448 13852
rect 28442 13812 28448 13824
rect 28500 13812 28506 13864
rect 29196 13852 29224 13960
rect 29733 13923 29791 13929
rect 29733 13889 29745 13923
rect 29779 13889 29791 13923
rect 29840 13920 29868 13960
rect 30098 13948 30104 14000
rect 30156 13988 30162 14000
rect 30285 13991 30343 13997
rect 30285 13988 30297 13991
rect 30156 13960 30297 13988
rect 30156 13948 30162 13960
rect 30285 13957 30297 13960
rect 30331 13957 30343 13991
rect 30285 13951 30343 13957
rect 30193 13923 30251 13929
rect 30193 13920 30205 13923
rect 29840 13892 30205 13920
rect 29733 13883 29791 13889
rect 30193 13889 30205 13892
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 28552 13824 29224 13852
rect 28552 13784 28580 13824
rect 29454 13812 29460 13864
rect 29512 13852 29518 13864
rect 29748 13852 29776 13883
rect 30374 13880 30380 13932
rect 30432 13920 30438 13932
rect 30837 13923 30895 13929
rect 30837 13920 30849 13923
rect 30432 13892 30849 13920
rect 30432 13880 30438 13892
rect 30837 13889 30849 13892
rect 30883 13889 30895 13923
rect 30837 13883 30895 13889
rect 35713 13923 35771 13929
rect 35713 13889 35725 13923
rect 35759 13920 35771 13923
rect 36354 13920 36360 13932
rect 35759 13892 36360 13920
rect 35759 13889 35771 13892
rect 35713 13883 35771 13889
rect 36354 13880 36360 13892
rect 36412 13880 36418 13932
rect 31389 13855 31447 13861
rect 31389 13852 31401 13855
rect 29512 13824 31401 13852
rect 29512 13812 29518 13824
rect 31389 13821 31401 13824
rect 31435 13821 31447 13855
rect 31389 13815 31447 13821
rect 31570 13784 31576 13796
rect 27816 13756 28580 13784
rect 29472 13756 31576 13784
rect 25004 13744 25010 13756
rect 26234 13716 26240 13728
rect 18472 13688 26240 13716
rect 18472 13676 18478 13688
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 26510 13676 26516 13728
rect 26568 13716 26574 13728
rect 29472 13716 29500 13756
rect 31570 13744 31576 13756
rect 31628 13744 31634 13796
rect 29638 13716 29644 13728
rect 26568 13688 29500 13716
rect 29599 13688 29644 13716
rect 26568 13676 26574 13688
rect 29638 13676 29644 13688
rect 29696 13676 29702 13728
rect 1104 13626 36892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36892 13626
rect 1104 13552 36892 13574
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11698 13512 11704 13524
rect 11020 13484 11704 13512
rect 11020 13472 11026 13484
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 17402 13512 17408 13524
rect 12124 13484 17408 13512
rect 12124 13472 12130 13484
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 18874 13512 18880 13524
rect 18835 13484 18880 13512
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 19306 13484 21956 13512
rect 8389 13447 8447 13453
rect 8389 13413 8401 13447
rect 8435 13444 8447 13447
rect 12710 13444 12716 13456
rect 8435 13416 12716 13444
rect 8435 13413 8447 13416
rect 8389 13407 8447 13413
rect 11716 13385 11744 13416
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 13722 13404 13728 13456
rect 13780 13444 13786 13456
rect 15838 13444 15844 13456
rect 13780 13416 15844 13444
rect 13780 13404 13786 13416
rect 15838 13404 15844 13416
rect 15896 13404 15902 13456
rect 17497 13447 17555 13453
rect 17497 13413 17509 13447
rect 17543 13444 17555 13447
rect 19306 13444 19334 13484
rect 17543 13416 19334 13444
rect 17543 13413 17555 13416
rect 17497 13407 17555 13413
rect 20714 13404 20720 13456
rect 20772 13444 20778 13456
rect 21928 13444 21956 13484
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22922 13512 22928 13524
rect 22060 13484 22928 13512
rect 22060 13472 22066 13484
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 23845 13515 23903 13521
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 24854 13512 24860 13524
rect 23891 13484 24860 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 25314 13512 25320 13524
rect 25275 13484 25320 13512
rect 25314 13472 25320 13484
rect 25372 13472 25378 13524
rect 31570 13512 31576 13524
rect 25884 13484 29868 13512
rect 31531 13484 31576 13512
rect 22830 13444 22836 13456
rect 20772 13416 21864 13444
rect 21928 13416 22836 13444
rect 20772 13404 20778 13416
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 11701 13379 11759 13385
rect 9907 13348 11284 13376
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 1946 13268 1952 13320
rect 2004 13308 2010 13320
rect 8297 13311 8355 13317
rect 8297 13308 8309 13311
rect 2004 13280 8309 13308
rect 2004 13268 2010 13280
rect 8297 13277 8309 13280
rect 8343 13277 8355 13311
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 8297 13271 8355 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9548 13280 9781 13308
rect 9548 13268 9554 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 9217 13243 9275 13249
rect 9217 13209 9229 13243
rect 9263 13240 9275 13243
rect 10413 13243 10471 13249
rect 9263 13212 10364 13240
rect 9263 13209 9275 13212
rect 9217 13203 9275 13209
rect 10336 13172 10364 13212
rect 10413 13209 10425 13243
rect 10459 13240 10471 13243
rect 10778 13240 10784 13252
rect 10459 13212 10784 13240
rect 10459 13209 10471 13212
rect 10413 13203 10471 13209
rect 10778 13200 10784 13212
rect 10836 13200 10842 13252
rect 10965 13243 11023 13249
rect 10965 13209 10977 13243
rect 11011 13209 11023 13243
rect 10965 13203 11023 13209
rect 10980 13172 11008 13203
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11112 13212 11157 13240
rect 11112 13200 11118 13212
rect 10336 13144 11008 13172
rect 11256 13172 11284 13348
rect 11701 13345 11713 13379
rect 11747 13345 11759 13379
rect 12158 13376 12164 13388
rect 12119 13348 12164 13376
rect 11701 13339 11759 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12406 13348 13093 13376
rect 11793 13243 11851 13249
rect 11793 13209 11805 13243
rect 11839 13209 11851 13243
rect 11793 13203 11851 13209
rect 11808 13172 11836 13203
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 12406 13240 12434 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13354 13376 13360 13388
rect 13315 13348 13360 13376
rect 13081 13339 13139 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 13538 13336 13544 13388
rect 13596 13376 13602 13388
rect 13998 13376 14004 13388
rect 13596 13348 14004 13376
rect 13596 13336 13602 13348
rect 13998 13336 14004 13348
rect 14056 13376 14062 13388
rect 14369 13379 14427 13385
rect 14369 13376 14381 13379
rect 14056 13348 14381 13376
rect 14056 13336 14062 13348
rect 14369 13345 14381 13348
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15620 13348 15761 13376
rect 15620 13336 15626 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 16390 13376 16396 13388
rect 16351 13348 16396 13376
rect 15749 13339 15807 13345
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 19518 13376 19524 13388
rect 19479 13348 19524 13376
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19794 13376 19800 13388
rect 19755 13348 19800 13376
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 21082 13376 21088 13388
rect 20995 13348 21088 13376
rect 21082 13336 21088 13348
rect 21140 13376 21146 13388
rect 21450 13376 21456 13388
rect 21140 13348 21456 13376
rect 21140 13336 21146 13348
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 21726 13376 21732 13388
rect 21687 13348 21732 13376
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 21836 13376 21864 13416
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 23566 13404 23572 13456
rect 23624 13444 23630 13456
rect 25884 13444 25912 13484
rect 23624 13416 25912 13444
rect 23624 13404 23630 13416
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 29840 13453 29868 13484
rect 31570 13472 31576 13484
rect 31628 13472 31634 13524
rect 29825 13447 29883 13453
rect 26016 13416 29316 13444
rect 26016 13404 26022 13416
rect 24673 13379 24731 13385
rect 24673 13376 24685 13379
rect 21836 13348 24685 13376
rect 24673 13345 24685 13348
rect 24719 13345 24731 13379
rect 24673 13339 24731 13345
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 27430 13376 27436 13388
rect 24912 13348 27436 13376
rect 24912 13336 24918 13348
rect 27430 13336 27436 13348
rect 27488 13336 27494 13388
rect 27522 13336 27528 13388
rect 27580 13376 27586 13388
rect 27893 13379 27951 13385
rect 27893 13376 27905 13379
rect 27580 13348 27905 13376
rect 27580 13336 27586 13348
rect 27893 13345 27905 13348
rect 27939 13345 27951 13379
rect 27893 13339 27951 13345
rect 28074 13336 28080 13388
rect 28132 13376 28138 13388
rect 28169 13379 28227 13385
rect 28169 13376 28181 13379
rect 28132 13348 28181 13376
rect 28132 13336 28138 13348
rect 28169 13345 28181 13348
rect 28215 13345 28227 13379
rect 28169 13339 28227 13345
rect 29089 13379 29147 13385
rect 29089 13345 29101 13379
rect 29135 13376 29147 13379
rect 29178 13376 29184 13388
rect 29135 13348 29184 13376
rect 29135 13345 29147 13348
rect 29089 13339 29147 13345
rect 29178 13336 29184 13348
rect 29236 13336 29242 13388
rect 12894 13268 12900 13320
rect 12952 13268 12958 13320
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 19334 13308 19340 13320
rect 17644 13280 19340 13308
rect 17644 13268 17650 13280
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 23750 13308 23756 13320
rect 23711 13280 23756 13308
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 24486 13268 24492 13320
rect 24544 13308 24550 13320
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 24544 13280 24777 13308
rect 24544 13268 24550 13280
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 25225 13311 25283 13317
rect 25225 13277 25237 13311
rect 25271 13308 25283 13311
rect 25682 13308 25688 13320
rect 25271 13280 25688 13308
rect 25271 13277 25283 13280
rect 25225 13271 25283 13277
rect 25682 13268 25688 13280
rect 25740 13268 25746 13320
rect 26326 13308 26332 13320
rect 25792 13280 26332 13308
rect 12032 13212 12434 13240
rect 12912 13240 12940 13268
rect 13150 13243 13208 13249
rect 13150 13240 13162 13243
rect 12912 13212 13162 13240
rect 12032 13200 12038 13212
rect 13150 13209 13162 13212
rect 13196 13209 13208 13243
rect 13150 13203 13208 13209
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13209 14519 13243
rect 15010 13240 15016 13252
rect 14923 13212 15016 13240
rect 14461 13203 14519 13209
rect 11256 13144 11836 13172
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 14476 13172 14504 13203
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 15838 13200 15844 13252
rect 15896 13240 15902 13252
rect 15896 13212 15941 13240
rect 15896 13200 15902 13212
rect 16666 13200 16672 13252
rect 16724 13240 16730 13252
rect 16945 13243 17003 13249
rect 16945 13240 16957 13243
rect 16724 13212 16957 13240
rect 16724 13200 16730 13212
rect 16945 13209 16957 13212
rect 16991 13209 17003 13243
rect 16945 13203 17003 13209
rect 17037 13243 17095 13249
rect 17037 13209 17049 13243
rect 17083 13209 17095 13243
rect 17037 13203 17095 13209
rect 12676 13144 14504 13172
rect 15028 13172 15056 13200
rect 16298 13172 16304 13184
rect 15028 13144 16304 13172
rect 12676 13132 12682 13144
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 16482 13132 16488 13184
rect 16540 13172 16546 13184
rect 17052 13172 17080 13203
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 18233 13243 18291 13249
rect 18233 13240 18245 13243
rect 17184 13212 18245 13240
rect 17184 13200 17190 13212
rect 18233 13209 18245 13212
rect 18279 13209 18291 13243
rect 18233 13203 18291 13209
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13209 19671 13243
rect 21177 13243 21235 13249
rect 21177 13240 21189 13243
rect 19613 13203 19671 13209
rect 21008 13212 21189 13240
rect 18138 13172 18144 13184
rect 16540 13144 17080 13172
rect 18099 13144 18144 13172
rect 16540 13132 16546 13144
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19621 13172 19649 13203
rect 21008 13184 21036 13212
rect 21177 13209 21189 13212
rect 21223 13209 21235 13243
rect 22278 13240 22284 13252
rect 22239 13212 22284 13240
rect 21177 13203 21235 13209
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 22373 13243 22431 13249
rect 22373 13209 22385 13243
rect 22419 13209 22431 13243
rect 22922 13240 22928 13252
rect 22835 13212 22928 13240
rect 22373 13203 22431 13209
rect 19392 13144 19649 13172
rect 19392 13132 19398 13144
rect 20990 13132 20996 13184
rect 21048 13132 21054 13184
rect 21358 13132 21364 13184
rect 21416 13172 21422 13184
rect 22388 13172 22416 13203
rect 22922 13200 22928 13212
rect 22980 13240 22986 13252
rect 25792 13240 25820 13280
rect 26326 13268 26332 13280
rect 26384 13268 26390 13320
rect 28994 13308 29000 13320
rect 28955 13280 29000 13308
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 29288 13308 29316 13416
rect 29825 13413 29837 13447
rect 29871 13444 29883 13447
rect 30374 13444 30380 13456
rect 29871 13416 30380 13444
rect 29871 13413 29883 13416
rect 29825 13407 29883 13413
rect 30374 13404 30380 13416
rect 30432 13404 30438 13456
rect 36170 13376 36176 13388
rect 31726 13348 36176 13376
rect 31113 13311 31171 13317
rect 29288 13280 29776 13308
rect 26234 13240 26240 13252
rect 22980 13212 25820 13240
rect 26195 13212 26240 13240
rect 22980 13200 22986 13212
rect 26234 13200 26240 13212
rect 26292 13200 26298 13252
rect 27157 13243 27215 13249
rect 27157 13209 27169 13243
rect 27203 13209 27215 13243
rect 27157 13203 27215 13209
rect 27249 13243 27307 13249
rect 27249 13209 27261 13243
rect 27295 13240 27307 13243
rect 27706 13240 27712 13252
rect 27295 13212 27712 13240
rect 27295 13209 27307 13212
rect 27249 13203 27307 13209
rect 21416 13144 22416 13172
rect 21416 13132 21422 13144
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 27062 13172 27068 13184
rect 22520 13144 27068 13172
rect 22520 13132 22526 13144
rect 27062 13132 27068 13144
rect 27120 13132 27126 13184
rect 27172 13172 27200 13203
rect 27706 13200 27712 13212
rect 27764 13200 27770 13252
rect 27982 13200 27988 13252
rect 28040 13240 28046 13252
rect 29638 13240 29644 13252
rect 28040 13212 28085 13240
rect 28644 13212 29644 13240
rect 28040 13200 28046 13212
rect 28644 13172 28672 13212
rect 29638 13200 29644 13212
rect 29696 13200 29702 13252
rect 27172 13144 28672 13172
rect 29748 13172 29776 13280
rect 31113 13277 31125 13311
rect 31159 13308 31171 13311
rect 31726 13308 31754 13348
rect 36170 13336 36176 13348
rect 36228 13336 36234 13388
rect 31159 13280 31754 13308
rect 31159 13277 31171 13280
rect 31113 13271 31171 13277
rect 30282 13240 30288 13252
rect 30243 13212 30288 13240
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 30377 13243 30435 13249
rect 30377 13209 30389 13243
rect 30423 13240 30435 13243
rect 31021 13243 31079 13249
rect 31021 13240 31033 13243
rect 30423 13212 31033 13240
rect 30423 13209 30435 13212
rect 30377 13203 30435 13209
rect 31021 13209 31033 13212
rect 31067 13209 31079 13243
rect 31021 13203 31079 13209
rect 30392 13172 30420 13203
rect 29748 13144 30420 13172
rect 31570 13132 31576 13184
rect 31628 13172 31634 13184
rect 35894 13172 35900 13184
rect 31628 13144 35900 13172
rect 31628 13132 31634 13144
rect 35894 13132 35900 13144
rect 35952 13132 35958 13184
rect 1104 13082 36892 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 36892 13082
rect 1104 13008 36892 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 2133 12971 2191 12977
rect 2133 12968 2145 12971
rect 1912 12940 2145 12968
rect 1912 12928 1918 12940
rect 2133 12937 2145 12940
rect 2179 12937 2191 12971
rect 2869 12971 2927 12977
rect 2869 12968 2881 12971
rect 2133 12931 2191 12937
rect 2746 12940 2881 12968
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2746 12832 2774 12940
rect 2869 12937 2881 12940
rect 2915 12968 2927 12971
rect 4798 12968 4804 12980
rect 2915 12940 4804 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 4798 12928 4804 12940
rect 4856 12968 4862 12980
rect 8021 12971 8079 12977
rect 8021 12968 8033 12971
rect 4856 12940 8033 12968
rect 4856 12928 4862 12940
rect 8021 12937 8033 12940
rect 8067 12968 8079 12971
rect 8386 12968 8392 12980
rect 8067 12940 8392 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 9769 12971 9827 12977
rect 9769 12937 9781 12971
rect 9815 12968 9827 12971
rect 11882 12968 11888 12980
rect 9815 12940 11888 12968
rect 9815 12937 9827 12940
rect 9769 12931 9827 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12066 12968 12072 12980
rect 12027 12940 12072 12968
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 12400 12940 15792 12968
rect 12400 12928 12406 12940
rect 11422 12900 11428 12912
rect 10520 12872 11428 12900
rect 2363 12804 2774 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8352 12804 8677 12832
rect 8352 12792 8358 12804
rect 8665 12801 8677 12804
rect 8711 12832 8723 12835
rect 9490 12832 9496 12844
rect 8711 12804 9496 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 9490 12792 9496 12804
rect 9548 12832 9554 12844
rect 9677 12835 9735 12841
rect 9677 12832 9689 12835
rect 9548 12804 9689 12832
rect 9548 12792 9554 12804
rect 9677 12801 9689 12804
rect 9723 12832 9735 12835
rect 9858 12832 9864 12844
rect 9723 12804 9864 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10520 12841 10548 12872
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 12805 12903 12863 12909
rect 12805 12900 12817 12903
rect 12406 12872 12817 12900
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 10980 12764 11008 12795
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 11664 12804 11989 12832
rect 11664 12792 11670 12804
rect 11977 12801 11989 12804
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 12406 12832 12434 12872
rect 12805 12869 12817 12872
rect 12851 12869 12863 12903
rect 12805 12863 12863 12869
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 14826 12900 14832 12912
rect 12952 12872 14832 12900
rect 12952 12860 12958 12872
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 14921 12903 14979 12909
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 15470 12900 15476 12912
rect 14967 12872 15476 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 15764 12909 15792 12940
rect 16316 12940 18920 12968
rect 16316 12909 16344 12940
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12869 15807 12903
rect 15749 12863 15807 12869
rect 16301 12903 16359 12909
rect 16301 12869 16313 12903
rect 16347 12869 16359 12903
rect 16301 12863 16359 12869
rect 16850 12860 16856 12912
rect 16908 12900 16914 12912
rect 17218 12900 17224 12912
rect 16908 12872 17224 12900
rect 16908 12860 16914 12872
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 17494 12900 17500 12912
rect 17455 12872 17500 12900
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 18414 12900 18420 12912
rect 18375 12872 18420 12900
rect 18414 12860 18420 12872
rect 18472 12860 18478 12912
rect 18892 12900 18920 12940
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19245 12971 19303 12977
rect 19245 12968 19257 12971
rect 19024 12940 19257 12968
rect 19024 12928 19030 12940
rect 19245 12937 19257 12940
rect 19291 12937 19303 12971
rect 21358 12968 21364 12980
rect 19245 12931 19303 12937
rect 19444 12940 20760 12968
rect 21319 12940 21364 12968
rect 19444 12900 19472 12940
rect 18892 12872 19472 12900
rect 19518 12860 19524 12912
rect 19576 12900 19582 12912
rect 20625 12903 20683 12909
rect 20625 12900 20637 12903
rect 19576 12872 20637 12900
rect 19576 12860 19582 12872
rect 20625 12869 20637 12872
rect 20671 12869 20683 12903
rect 20732 12900 20760 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 27249 12971 27307 12977
rect 27249 12968 27261 12971
rect 24872 12940 27261 12968
rect 21726 12900 21732 12912
rect 20732 12872 21732 12900
rect 20625 12863 20683 12869
rect 21726 12860 21732 12872
rect 21784 12860 21790 12912
rect 22373 12903 22431 12909
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 24872 12900 24900 12940
rect 27249 12937 27261 12940
rect 27295 12937 27307 12971
rect 27249 12931 27307 12937
rect 27430 12928 27436 12980
rect 27488 12968 27494 12980
rect 28537 12971 28595 12977
rect 28537 12968 28549 12971
rect 27488 12940 28549 12968
rect 27488 12928 27494 12940
rect 28537 12937 28549 12940
rect 28583 12937 28595 12971
rect 28537 12931 28595 12937
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 29825 12971 29883 12977
rect 29825 12968 29837 12971
rect 29788 12940 29837 12968
rect 29788 12928 29794 12940
rect 29825 12937 29837 12940
rect 29871 12937 29883 12971
rect 29825 12931 29883 12937
rect 30282 12928 30288 12980
rect 30340 12968 30346 12980
rect 31113 12971 31171 12977
rect 31113 12968 31125 12971
rect 30340 12940 31125 12968
rect 30340 12928 30346 12940
rect 31113 12937 31125 12940
rect 31159 12937 31171 12971
rect 31113 12931 31171 12937
rect 31570 12928 31576 12980
rect 31628 12968 31634 12980
rect 31757 12971 31815 12977
rect 31757 12968 31769 12971
rect 31628 12940 31769 12968
rect 31628 12928 31634 12940
rect 31757 12937 31769 12940
rect 31803 12968 31815 12971
rect 35342 12968 35348 12980
rect 31803 12940 35348 12968
rect 31803 12937 31815 12940
rect 31757 12931 31815 12937
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 22419 12872 24900 12900
rect 25961 12903 26019 12909
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 25961 12869 25973 12903
rect 26007 12900 26019 12903
rect 26050 12900 26056 12912
rect 26007 12872 26056 12900
rect 26007 12869 26019 12872
rect 25961 12863 26019 12869
rect 26050 12860 26056 12872
rect 26108 12860 26114 12912
rect 29089 12903 29147 12909
rect 29089 12900 29101 12903
rect 26252 12872 29101 12900
rect 12124 12804 12434 12832
rect 12124 12792 12130 12804
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19337 12835 19395 12841
rect 19337 12832 19349 12835
rect 18932 12804 19349 12832
rect 18932 12792 18938 12804
rect 19337 12801 19349 12804
rect 19383 12832 19395 12835
rect 19426 12832 19432 12844
rect 19383 12804 19432 12832
rect 19383 12801 19395 12804
rect 19337 12795 19395 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 21232 12804 21281 12832
rect 21232 12792 21238 12804
rect 21269 12801 21281 12804
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12832 22983 12835
rect 23474 12832 23480 12844
rect 22971 12804 23480 12832
rect 22971 12801 22983 12804
rect 22925 12795 22983 12801
rect 9263 12736 12296 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 11057 12699 11115 12705
rect 11057 12665 11069 12699
rect 11103 12696 11115 12699
rect 12268 12696 12296 12736
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 12400 12736 12725 12764
rect 12400 12724 12406 12736
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 12434 12696 12440 12708
rect 11103 12668 12204 12696
rect 12268 12668 12440 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 12066 12628 12072 12640
rect 10459 12600 12072 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 12176 12628 12204 12668
rect 12434 12656 12440 12668
rect 12492 12656 12498 12708
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 13004 12696 13032 12727
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 13412 12736 14228 12764
rect 13412 12724 13418 12736
rect 13722 12696 13728 12708
rect 12584 12668 13728 12696
rect 12584 12656 12590 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14200 12696 14228 12736
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14332 12736 14381 12764
rect 14332 12724 14338 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 15028 12696 15056 12727
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 15252 12736 15669 12764
rect 15252 12724 15258 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 15896 12736 17417 12764
rect 15896 12724 15902 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 18012 12736 20453 12764
rect 18012 12724 18018 12736
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 20714 12764 20720 12776
rect 20675 12736 20720 12764
rect 20441 12727 20499 12733
rect 19058 12696 19064 12708
rect 14200 12668 19064 12696
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 19794 12656 19800 12708
rect 19852 12696 19858 12708
rect 20456 12696 20484 12727
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 21284 12696 21312 12795
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12832 23627 12835
rect 23750 12832 23756 12844
rect 23615 12804 23756 12832
rect 23615 12801 23627 12804
rect 23569 12795 23627 12801
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 24026 12832 24032 12844
rect 23987 12804 24032 12832
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 24210 12792 24216 12844
rect 24268 12832 24274 12844
rect 24765 12835 24823 12841
rect 24765 12832 24777 12835
rect 24268 12804 24777 12832
rect 24268 12792 24274 12804
rect 24765 12801 24777 12804
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 25406 12832 25412 12844
rect 24903 12804 25412 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 21450 12724 21456 12776
rect 21508 12764 21514 12776
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 21508 12736 22293 12764
rect 21508 12724 21514 12736
rect 22281 12733 22293 12736
rect 22327 12764 22339 12767
rect 22370 12764 22376 12776
rect 22327 12736 22376 12764
rect 22327 12733 22339 12736
rect 22281 12727 22339 12733
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 25593 12767 25651 12773
rect 25593 12764 25605 12767
rect 23716 12736 25605 12764
rect 23716 12724 23722 12736
rect 25593 12733 25605 12736
rect 25639 12733 25651 12767
rect 25593 12727 25651 12733
rect 25958 12724 25964 12776
rect 26016 12764 26022 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 26016 12736 26065 12764
rect 26016 12724 26022 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 23382 12696 23388 12708
rect 19852 12668 20024 12696
rect 20456 12668 21220 12696
rect 21284 12668 23388 12696
rect 19852 12656 19858 12668
rect 13630 12628 13636 12640
rect 12176 12600 13636 12628
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12628 13967 12631
rect 16114 12628 16120 12640
rect 13955 12600 16120 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 16114 12588 16120 12600
rect 16172 12628 16178 12640
rect 18874 12628 18880 12640
rect 16172 12600 18880 12628
rect 16172 12588 16178 12600
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 19886 12628 19892 12640
rect 19024 12600 19892 12628
rect 19024 12588 19030 12600
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 19996 12628 20024 12668
rect 20438 12628 20444 12640
rect 19996 12600 20444 12628
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 21192 12628 21220 12668
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 23477 12699 23535 12705
rect 23477 12665 23489 12699
rect 23523 12696 23535 12699
rect 24578 12696 24584 12708
rect 23523 12668 24584 12696
rect 23523 12665 23535 12668
rect 23477 12659 23535 12665
rect 24578 12656 24584 12668
rect 24636 12656 24642 12708
rect 26142 12656 26148 12708
rect 26200 12696 26206 12708
rect 26252 12696 26280 12872
rect 29089 12869 29101 12872
rect 29135 12869 29147 12903
rect 29089 12863 29147 12869
rect 27062 12792 27068 12844
rect 27120 12832 27126 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 27120 12804 27353 12832
rect 27120 12792 27126 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27430 12792 27436 12844
rect 27488 12832 27494 12844
rect 27801 12835 27859 12841
rect 27801 12832 27813 12835
rect 27488 12804 27813 12832
rect 27488 12792 27494 12804
rect 27801 12801 27813 12804
rect 27847 12801 27859 12835
rect 27801 12795 27859 12801
rect 28629 12835 28687 12841
rect 28629 12801 28641 12835
rect 28675 12832 28687 12835
rect 28718 12832 28724 12844
rect 28675 12804 28724 12832
rect 28675 12801 28687 12804
rect 28629 12795 28687 12801
rect 28718 12792 28724 12804
rect 28776 12792 28782 12844
rect 29270 12792 29276 12844
rect 29328 12832 29334 12844
rect 29733 12835 29791 12841
rect 29733 12832 29745 12835
rect 29328 12804 29745 12832
rect 29328 12792 29334 12804
rect 29733 12801 29745 12804
rect 29779 12801 29791 12835
rect 29733 12795 29791 12801
rect 30466 12792 30472 12844
rect 30524 12832 30530 12844
rect 30561 12835 30619 12841
rect 30561 12832 30573 12835
rect 30524 12804 30573 12832
rect 30524 12792 30530 12804
rect 30561 12801 30573 12804
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 26326 12724 26332 12776
rect 26384 12764 26390 12776
rect 27893 12767 27951 12773
rect 27893 12764 27905 12767
rect 26384 12736 27905 12764
rect 26384 12724 26390 12736
rect 27893 12733 27905 12736
rect 27939 12733 27951 12767
rect 30576 12764 30604 12795
rect 30742 12792 30748 12844
rect 30800 12832 30806 12844
rect 31205 12835 31263 12841
rect 31205 12832 31217 12835
rect 30800 12804 31217 12832
rect 30800 12792 30806 12804
rect 31205 12801 31217 12804
rect 31251 12832 31263 12835
rect 32309 12835 32367 12841
rect 32309 12832 32321 12835
rect 31251 12804 32321 12832
rect 31251 12801 31263 12804
rect 31205 12795 31263 12801
rect 32309 12801 32321 12804
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 31570 12764 31576 12776
rect 30576 12736 31576 12764
rect 27893 12727 27951 12733
rect 31570 12724 31576 12736
rect 31628 12724 31634 12776
rect 26200 12668 26280 12696
rect 26200 12656 26206 12668
rect 27062 12656 27068 12708
rect 27120 12696 27126 12708
rect 30926 12696 30932 12708
rect 27120 12668 30932 12696
rect 27120 12656 27126 12668
rect 30926 12656 30932 12668
rect 30984 12656 30990 12708
rect 22830 12628 22836 12640
rect 21192 12600 22836 12628
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 24121 12631 24179 12637
rect 24121 12597 24133 12631
rect 24167 12628 24179 12631
rect 25130 12628 25136 12640
rect 24167 12600 25136 12628
rect 24167 12597 24179 12600
rect 24121 12591 24179 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 25314 12588 25320 12640
rect 25372 12628 25378 12640
rect 27430 12628 27436 12640
rect 25372 12600 27436 12628
rect 25372 12588 25378 12600
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 30377 12631 30435 12637
rect 30377 12597 30389 12631
rect 30423 12628 30435 12631
rect 30650 12628 30656 12640
rect 30423 12600 30656 12628
rect 30423 12597 30435 12600
rect 30377 12591 30435 12597
rect 30650 12588 30656 12600
rect 30708 12588 30714 12640
rect 1104 12538 36892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36892 12538
rect 1104 12464 36892 12486
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 13078 12424 13084 12436
rect 10796 12396 13084 12424
rect 8294 12288 8300 12300
rect 7760 12260 8300 12288
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 7760 12229 7788 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 10796 12288 10824 12396
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 13780 12396 16160 12424
rect 13780 12384 13786 12396
rect 9324 12260 10824 12288
rect 11256 12328 12204 12356
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7331 12192 7757 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 7745 12183 7803 12189
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 9324 12229 9352 12260
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8720 12192 9321 12220
rect 8720 12180 8726 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9916 12192 9965 12220
rect 9916 12180 9922 12192
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10744 12192 10793 12220
rect 10744 12180 10750 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 11256 12229 11284 12328
rect 12066 12288 12072 12300
rect 12027 12260 12072 12288
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12176 12288 12204 12328
rect 12250 12316 12256 12368
rect 12308 12356 12314 12368
rect 15194 12356 15200 12368
rect 12308 12328 15200 12356
rect 12308 12316 12314 12328
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 16132 12365 16160 12396
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 20165 12427 20223 12433
rect 16356 12396 20116 12424
rect 16356 12384 16362 12396
rect 16117 12359 16175 12365
rect 16117 12325 16129 12359
rect 16163 12325 16175 12359
rect 16117 12319 16175 12325
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 18785 12359 18843 12365
rect 16724 12328 18736 12356
rect 16724 12316 16730 12328
rect 13170 12288 13176 12300
rect 12176 12260 13176 12288
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13446 12288 13452 12300
rect 13407 12260 13452 12288
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 13556 12260 14657 12288
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 11204 12192 11253 12220
rect 11204 12180 11210 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11606 12220 11612 12232
rect 11388 12192 11612 12220
rect 11388 12180 11394 12192
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 13556 12220 13584 12260
rect 14645 12257 14657 12260
rect 14691 12288 14703 12291
rect 17313 12291 17371 12297
rect 17313 12288 17325 12291
rect 14691 12260 17325 12288
rect 14691 12257 14703 12260
rect 14645 12251 14703 12257
rect 17313 12257 17325 12260
rect 17359 12257 17371 12291
rect 18708 12288 18736 12328
rect 18785 12325 18797 12359
rect 18831 12356 18843 12359
rect 19794 12356 19800 12368
rect 18831 12328 19800 12356
rect 18831 12325 18843 12328
rect 18785 12319 18843 12325
rect 19794 12316 19800 12328
rect 19852 12316 19858 12368
rect 19242 12288 19248 12300
rect 18708 12260 19248 12288
rect 17313 12251 17371 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19518 12288 19524 12300
rect 19479 12260 19524 12288
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 20088 12288 20116 12396
rect 20165 12393 20177 12427
rect 20211 12424 20223 12427
rect 20530 12424 20536 12436
rect 20211 12396 20536 12424
rect 20211 12393 20223 12396
rect 20165 12387 20223 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 21818 12424 21824 12436
rect 21779 12396 21824 12424
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 23014 12424 23020 12436
rect 21928 12396 23020 12424
rect 21269 12359 21327 12365
rect 21269 12325 21281 12359
rect 21315 12356 21327 12359
rect 21928 12356 21956 12396
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 24762 12384 24768 12436
rect 24820 12424 24826 12436
rect 29086 12424 29092 12436
rect 24820 12396 29092 12424
rect 24820 12384 24826 12396
rect 29086 12384 29092 12396
rect 29144 12384 29150 12436
rect 30926 12424 30932 12436
rect 30887 12396 30932 12424
rect 30926 12384 30932 12396
rect 30984 12384 30990 12436
rect 31570 12424 31576 12436
rect 31531 12396 31576 12424
rect 31570 12384 31576 12396
rect 31628 12384 31634 12436
rect 30466 12356 30472 12368
rect 21315 12328 21956 12356
rect 22020 12328 26832 12356
rect 21315 12325 21327 12328
rect 21269 12319 21327 12325
rect 22020 12288 22048 12328
rect 20088 12260 22048 12288
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 23017 12291 23075 12297
rect 23017 12288 23029 12291
rect 22888 12260 23029 12288
rect 22888 12248 22894 12260
rect 23017 12257 23029 12260
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 26142 12288 26148 12300
rect 25271 12260 26148 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 26142 12248 26148 12260
rect 26200 12248 26206 12300
rect 12400 12192 13584 12220
rect 12400 12180 12406 12192
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 15289 12223 15347 12229
rect 13688 12192 13733 12220
rect 13688 12180 13694 12192
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 16022 12220 16028 12232
rect 15335 12192 16028 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12220 18751 12223
rect 19150 12220 19156 12232
rect 18739 12192 19156 12220
rect 18739 12189 18751 12192
rect 18693 12183 18751 12189
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12220 19490 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19484 12192 20085 12220
rect 19484 12180 19490 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 20312 12192 21189 12220
rect 20312 12180 20318 12192
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 21324 12192 22385 12220
rect 21324 12180 21330 12192
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 23382 12180 23388 12232
rect 23440 12220 23446 12232
rect 23753 12223 23811 12229
rect 23753 12220 23765 12223
rect 23440 12192 23765 12220
rect 23440 12180 23446 12192
rect 23753 12189 23765 12192
rect 23799 12189 23811 12223
rect 23753 12183 23811 12189
rect 25406 12180 25412 12232
rect 25464 12220 25470 12232
rect 25682 12220 25688 12232
rect 25464 12192 25688 12220
rect 25464 12180 25470 12192
rect 25682 12180 25688 12192
rect 25740 12180 25746 12232
rect 26513 12223 26571 12229
rect 26513 12189 26525 12223
rect 26559 12189 26571 12223
rect 26513 12183 26571 12189
rect 8481 12155 8539 12161
rect 8481 12121 8493 12155
rect 8527 12152 8539 12155
rect 13538 12152 13544 12164
rect 8527 12124 13544 12152
rect 8527 12121 8539 12124
rect 8481 12115 8539 12121
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 14734 12152 14740 12164
rect 14695 12124 14740 12152
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 16574 12152 16580 12164
rect 16535 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 16666 12112 16672 12164
rect 16724 12152 16730 12164
rect 16724 12124 16769 12152
rect 16724 12112 16730 12124
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 17405 12155 17463 12161
rect 17405 12152 17417 12155
rect 16908 12124 17417 12152
rect 16908 12112 16914 12124
rect 17405 12121 17417 12124
rect 17451 12121 17463 12155
rect 17405 12115 17463 12121
rect 17957 12155 18015 12161
rect 17957 12121 17969 12155
rect 18003 12152 18015 12155
rect 22922 12152 22928 12164
rect 18003 12124 22784 12152
rect 22883 12124 22928 12152
rect 18003 12121 18015 12124
rect 17957 12115 18015 12121
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 1854 12084 1860 12096
rect 1811 12056 1860 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 7837 12087 7895 12093
rect 7837 12053 7849 12087
rect 7883 12084 7895 12087
rect 8018 12084 8024 12096
rect 7883 12056 8024 12084
rect 7883 12053 7895 12056
rect 7837 12047 7895 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 9493 12087 9551 12093
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 9582 12084 9588 12096
rect 9539 12056 9588 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10045 12087 10103 12093
rect 10045 12053 10057 12087
rect 10091 12084 10103 12087
rect 11054 12084 11060 12096
rect 10091 12056 11060 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 12434 12084 12440 12096
rect 11379 12056 12440 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12989 12087 13047 12093
rect 12989 12084 13001 12087
rect 12584 12056 13001 12084
rect 12584 12044 12590 12056
rect 12989 12053 13001 12056
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 15930 12084 15936 12096
rect 15528 12056 15936 12084
rect 15528 12044 15534 12056
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 18782 12084 18788 12096
rect 16080 12056 18788 12084
rect 16080 12044 16086 12056
rect 18782 12044 18788 12056
rect 18840 12044 18846 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 21266 12084 21272 12096
rect 19300 12056 21272 12084
rect 19300 12044 19306 12056
rect 21266 12044 21272 12056
rect 21324 12044 21330 12096
rect 22756 12084 22784 12124
rect 22922 12112 22928 12124
rect 22980 12112 22986 12164
rect 24581 12155 24639 12161
rect 24581 12152 24593 12155
rect 23492 12124 24593 12152
rect 23492 12084 23520 12124
rect 24581 12121 24593 12124
rect 24627 12152 24639 12155
rect 24762 12152 24768 12164
rect 24627 12124 24768 12152
rect 24627 12121 24639 12124
rect 24581 12115 24639 12121
rect 24762 12112 24768 12124
rect 24820 12112 24826 12164
rect 25133 12155 25191 12161
rect 25133 12121 25145 12155
rect 25179 12152 25191 12155
rect 25590 12152 25596 12164
rect 25179 12124 25596 12152
rect 25179 12121 25191 12124
rect 25133 12115 25191 12121
rect 25590 12112 25596 12124
rect 25648 12112 25654 12164
rect 25774 12152 25780 12164
rect 25735 12124 25780 12152
rect 25774 12112 25780 12124
rect 25832 12112 25838 12164
rect 25961 12155 26019 12161
rect 25961 12121 25973 12155
rect 26007 12121 26019 12155
rect 25961 12115 26019 12121
rect 23658 12084 23664 12096
rect 22756 12056 23520 12084
rect 23619 12056 23664 12084
rect 23658 12044 23664 12056
rect 23716 12044 23722 12096
rect 23750 12044 23756 12096
rect 23808 12084 23814 12096
rect 24026 12084 24032 12096
rect 23808 12056 24032 12084
rect 23808 12044 23814 12056
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 25976 12084 26004 12115
rect 26142 12112 26148 12164
rect 26200 12152 26206 12164
rect 26528 12152 26556 12183
rect 26602 12180 26608 12232
rect 26660 12220 26666 12232
rect 26660 12192 26705 12220
rect 26660 12180 26666 12192
rect 26200 12124 26556 12152
rect 26804 12152 26832 12328
rect 28736 12328 30472 12356
rect 27062 12248 27068 12300
rect 27120 12288 27126 12300
rect 28629 12291 28687 12297
rect 28629 12288 28641 12291
rect 27120 12260 28641 12288
rect 27120 12248 27126 12260
rect 28629 12257 28641 12260
rect 28675 12257 28687 12291
rect 28629 12251 28687 12257
rect 28736 12229 28764 12328
rect 30466 12316 30472 12328
rect 30524 12316 30530 12368
rect 29825 12291 29883 12297
rect 29825 12257 29837 12291
rect 29871 12288 29883 12291
rect 29871 12260 31754 12288
rect 29871 12257 29883 12260
rect 29825 12251 29883 12257
rect 28721 12223 28779 12229
rect 28721 12189 28733 12223
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 31726 12164 31754 12260
rect 27433 12155 27491 12161
rect 27433 12152 27445 12155
rect 26804 12124 27445 12152
rect 26200 12112 26206 12124
rect 27433 12121 27445 12124
rect 27479 12121 27491 12155
rect 27433 12115 27491 12121
rect 27525 12155 27583 12161
rect 27525 12121 27537 12155
rect 27571 12121 27583 12155
rect 27525 12115 27583 12121
rect 28077 12155 28135 12161
rect 28077 12121 28089 12155
rect 28123 12152 28135 12155
rect 29638 12152 29644 12164
rect 28123 12124 29644 12152
rect 28123 12121 28135 12124
rect 28077 12115 28135 12121
rect 27338 12084 27344 12096
rect 25976 12056 27344 12084
rect 27338 12044 27344 12056
rect 27396 12044 27402 12096
rect 27540 12084 27568 12115
rect 29638 12112 29644 12124
rect 29696 12112 29702 12164
rect 29822 12112 29828 12164
rect 29880 12152 29886 12164
rect 29917 12155 29975 12161
rect 29917 12152 29929 12155
rect 29880 12124 29929 12152
rect 29880 12112 29886 12124
rect 29917 12121 29929 12124
rect 29963 12121 29975 12155
rect 30466 12152 30472 12164
rect 30379 12124 30472 12152
rect 29917 12115 29975 12121
rect 30466 12112 30472 12124
rect 30524 12152 30530 12164
rect 30650 12152 30656 12164
rect 30524 12124 30656 12152
rect 30524 12112 30530 12124
rect 30650 12112 30656 12124
rect 30708 12112 30714 12164
rect 31726 12152 31760 12164
rect 31667 12124 31760 12152
rect 31754 12112 31760 12124
rect 31812 12152 31818 12164
rect 31812 12124 32168 12152
rect 31812 12112 31818 12124
rect 28442 12084 28448 12096
rect 27540 12056 28448 12084
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 32140 12093 32168 12124
rect 32125 12087 32183 12093
rect 32125 12053 32137 12087
rect 32171 12084 32183 12087
rect 32398 12084 32404 12096
rect 32171 12056 32404 12084
rect 32171 12053 32183 12056
rect 32125 12047 32183 12053
rect 32398 12044 32404 12056
rect 32456 12044 32462 12096
rect 1104 11994 36892 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 36892 11994
rect 1104 11920 36892 11942
rect 8662 11880 8668 11892
rect 8623 11852 8668 11880
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9217 11883 9275 11889
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 11146 11880 11152 11892
rect 9263 11852 11152 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12400 11852 15700 11880
rect 12400 11840 12406 11852
rect 11330 11812 11336 11824
rect 10520 11784 11336 11812
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 8754 11744 8760 11756
rect 1903 11716 8760 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 10520 11753 10548 11784
rect 11330 11772 11336 11784
rect 11388 11772 11394 11824
rect 11514 11772 11520 11824
rect 11572 11812 11578 11824
rect 11885 11815 11943 11821
rect 11885 11812 11897 11815
rect 11572 11784 11897 11812
rect 11572 11772 11578 11784
rect 11885 11781 11897 11784
rect 11931 11781 11943 11815
rect 11885 11775 11943 11781
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 13265 11815 13323 11821
rect 13265 11812 13277 11815
rect 12492 11784 13277 11812
rect 12492 11772 12498 11784
rect 13265 11781 13277 11784
rect 13311 11781 13323 11815
rect 13265 11775 13323 11781
rect 13630 11772 13636 11824
rect 13688 11812 13694 11824
rect 14553 11815 14611 11821
rect 14553 11812 14565 11815
rect 13688 11784 14565 11812
rect 13688 11772 13694 11784
rect 14553 11781 14565 11784
rect 14599 11781 14611 11815
rect 14553 11775 14611 11781
rect 14642 11772 14648 11824
rect 14700 11812 14706 11824
rect 15672 11812 15700 11852
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 15804 11852 16221 11880
rect 15804 11840 15810 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 16209 11843 16267 11849
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 16816 11852 17785 11880
rect 16816 11840 16822 11852
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 17773 11843 17831 11849
rect 17880 11852 19932 11880
rect 17880 11812 17908 11852
rect 19904 11821 19932 11852
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 21048 11852 21189 11880
rect 21048 11840 21054 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 22189 11883 22247 11889
rect 22189 11849 22201 11883
rect 22235 11880 22247 11883
rect 22278 11880 22284 11892
rect 22235 11852 22284 11880
rect 22235 11849 22247 11852
rect 22189 11843 22247 11849
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 22738 11840 22744 11892
rect 22796 11880 22802 11892
rect 23382 11880 23388 11892
rect 22796 11852 23388 11880
rect 22796 11840 22802 11852
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 25038 11840 25044 11892
rect 25096 11880 25102 11892
rect 25869 11883 25927 11889
rect 25869 11880 25881 11883
rect 25096 11852 25881 11880
rect 25096 11840 25102 11852
rect 25869 11849 25881 11852
rect 25915 11849 25927 11883
rect 25869 11843 25927 11849
rect 26418 11840 26424 11892
rect 26476 11880 26482 11892
rect 26513 11883 26571 11889
rect 26513 11880 26525 11883
rect 26476 11852 26525 11880
rect 26476 11840 26482 11852
rect 26513 11849 26525 11852
rect 26559 11849 26571 11883
rect 27246 11880 27252 11892
rect 27207 11852 27252 11880
rect 26513 11843 26571 11849
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27798 11840 27804 11892
rect 27856 11880 27862 11892
rect 27893 11883 27951 11889
rect 27893 11880 27905 11883
rect 27856 11852 27905 11880
rect 27856 11840 27862 11852
rect 27893 11849 27905 11852
rect 27939 11849 27951 11883
rect 27893 11843 27951 11849
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 29825 11883 29883 11889
rect 29825 11880 29837 11883
rect 28500 11852 29837 11880
rect 28500 11840 28506 11852
rect 29825 11849 29837 11852
rect 29871 11849 29883 11883
rect 29825 11843 29883 11849
rect 18601 11815 18659 11821
rect 18601 11812 18613 11815
rect 14700 11784 14745 11812
rect 15672 11784 17908 11812
rect 18064 11784 18613 11812
rect 14700 11772 14706 11784
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 9876 11676 9904 11707
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10744 11716 10977 11744
rect 10744 11704 10750 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 13817 11747 13875 11753
rect 11112 11716 11560 11744
rect 11112 11704 11118 11716
rect 11532 11676 11560 11716
rect 13817 11713 13829 11747
rect 13863 11744 13875 11747
rect 14366 11744 14372 11756
rect 13863 11716 14372 11744
rect 13863 11713 13875 11716
rect 13817 11707 13875 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 15838 11744 15844 11756
rect 15212 11716 15844 11744
rect 11790 11676 11796 11688
rect 9876 11648 11192 11676
rect 11532 11648 11796 11676
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 9769 11611 9827 11617
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 10870 11608 10876 11620
rect 9815 11580 10876 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 10870 11568 10876 11580
rect 10928 11568 10934 11620
rect 11164 11608 11192 11648
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 12066 11676 12072 11688
rect 12027 11648 12072 11676
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12268 11648 12434 11676
rect 12268 11608 12296 11648
rect 11164 11580 12296 11608
rect 12406 11608 12434 11648
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 12768 11648 13185 11676
rect 12768 11636 12774 11648
rect 13173 11645 13185 11648
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 13320 11648 14841 11676
rect 13320 11636 13326 11648
rect 14829 11645 14841 11648
rect 14875 11676 14887 11679
rect 15212 11676 15240 11716
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16206 11744 16212 11756
rect 16163 11716 16212 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11713 17279 11747
rect 17862 11744 17868 11756
rect 17823 11716 17868 11744
rect 17221 11707 17279 11713
rect 14875 11648 15240 11676
rect 14875 11645 14887 11648
rect 14829 11639 14887 11645
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 16850 11676 16856 11688
rect 15344 11648 16856 11676
rect 15344 11636 15350 11648
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17236 11676 17264 11707
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 17954 11676 17960 11688
rect 17236 11648 17960 11676
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 13630 11608 13636 11620
rect 12406 11580 13636 11608
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 18064 11608 18092 11784
rect 18601 11781 18613 11784
rect 18647 11781 18659 11815
rect 18601 11775 18659 11781
rect 19889 11815 19947 11821
rect 19889 11781 19901 11815
rect 19935 11781 19947 11815
rect 20438 11812 20444 11824
rect 20399 11784 20444 11812
rect 19889 11775 19947 11781
rect 20438 11772 20444 11784
rect 20496 11772 20502 11824
rect 20533 11815 20591 11821
rect 20533 11781 20545 11815
rect 20579 11812 20591 11815
rect 20714 11812 20720 11824
rect 20579 11784 20720 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 22554 11772 22560 11824
rect 22612 11812 22618 11824
rect 23106 11812 23112 11824
rect 22612 11784 23112 11812
rect 22612 11772 22618 11784
rect 23106 11772 23112 11784
rect 23164 11812 23170 11824
rect 23201 11815 23259 11821
rect 23201 11812 23213 11815
rect 23164 11784 23213 11812
rect 23164 11772 23170 11784
rect 23201 11781 23213 11784
rect 23247 11781 23259 11815
rect 28537 11815 28595 11821
rect 28537 11812 28549 11815
rect 24426 11784 28549 11812
rect 23201 11775 23259 11781
rect 28537 11781 28549 11784
rect 28583 11781 28595 11815
rect 28537 11775 28595 11781
rect 28810 11772 28816 11824
rect 28868 11812 28874 11824
rect 30377 11815 30435 11821
rect 30377 11812 30389 11815
rect 28868 11784 30389 11812
rect 28868 11772 28874 11784
rect 30377 11781 30389 11784
rect 30423 11781 30435 11815
rect 30377 11775 30435 11781
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21910 11744 21916 11756
rect 21315 11716 21916 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 25222 11704 25228 11756
rect 25280 11704 25286 11756
rect 25317 11747 25375 11753
rect 25317 11713 25329 11747
rect 25363 11744 25375 11747
rect 25682 11744 25688 11756
rect 25363 11716 25688 11744
rect 25363 11713 25375 11716
rect 25317 11707 25375 11713
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 18506 11676 18512 11688
rect 18467 11648 18512 11676
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18782 11676 18788 11688
rect 18743 11648 18788 11676
rect 18782 11636 18788 11648
rect 18840 11676 18846 11688
rect 22922 11676 22928 11688
rect 18840 11648 22094 11676
rect 22883 11648 22928 11676
rect 18840 11636 18846 11648
rect 15488 11580 18092 11608
rect 22066 11608 22094 11648
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 25240 11676 25268 11704
rect 23032 11648 25268 11676
rect 23032 11608 23060 11648
rect 25792 11608 25820 11707
rect 26234 11704 26240 11756
rect 26292 11744 26298 11756
rect 26605 11747 26663 11753
rect 26605 11744 26617 11747
rect 26292 11716 26617 11744
rect 26292 11704 26298 11716
rect 26605 11713 26617 11716
rect 26651 11713 26663 11747
rect 27338 11744 27344 11756
rect 27299 11716 27344 11744
rect 26605 11707 26663 11713
rect 26620 11676 26648 11707
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 27522 11704 27528 11756
rect 27580 11744 27586 11756
rect 27985 11747 28043 11753
rect 27985 11744 27997 11747
rect 27580 11716 27997 11744
rect 27580 11704 27586 11716
rect 27985 11713 27997 11716
rect 28031 11744 28043 11747
rect 28166 11744 28172 11756
rect 28031 11716 28172 11744
rect 28031 11713 28043 11716
rect 27985 11707 28043 11713
rect 28166 11704 28172 11716
rect 28224 11704 28230 11756
rect 28442 11704 28448 11756
rect 28500 11744 28506 11756
rect 28629 11747 28687 11753
rect 28629 11744 28641 11747
rect 28500 11716 28641 11744
rect 28500 11704 28506 11716
rect 28629 11713 28641 11716
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 29273 11747 29331 11753
rect 29273 11713 29285 11747
rect 29319 11744 29331 11747
rect 29546 11744 29552 11756
rect 29319 11716 29552 11744
rect 29319 11713 29331 11716
rect 29273 11707 29331 11713
rect 29546 11704 29552 11716
rect 29604 11704 29610 11756
rect 29730 11744 29736 11756
rect 29691 11716 29736 11744
rect 29730 11704 29736 11716
rect 29788 11704 29794 11756
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11744 35679 11747
rect 36262 11744 36268 11756
rect 35667 11716 36268 11744
rect 35667 11713 35679 11716
rect 35621 11707 35679 11713
rect 36262 11704 36268 11716
rect 36320 11704 36326 11756
rect 30929 11679 30987 11685
rect 30929 11676 30941 11679
rect 26620 11648 30941 11676
rect 28644 11620 28672 11648
rect 30929 11645 30941 11648
rect 30975 11645 30987 11679
rect 30929 11639 30987 11645
rect 22066 11580 23060 11608
rect 24228 11580 25820 11608
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8202 11540 8208 11552
rect 8159 11512 8208 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8202 11500 8208 11512
rect 8260 11540 8266 11552
rect 10042 11540 10048 11552
rect 8260 11512 10048 11540
rect 8260 11500 8266 11512
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10410 11540 10416 11552
rect 10371 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 15488 11540 15516 11580
rect 11103 11512 15516 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 17129 11543 17187 11549
rect 17129 11540 17141 11543
rect 15804 11512 17141 11540
rect 15804 11500 15810 11512
rect 17129 11509 17141 11512
rect 17175 11509 17187 11543
rect 17129 11503 17187 11509
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 20070 11540 20076 11552
rect 17920 11512 20076 11540
rect 17920 11500 17926 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 24228 11540 24256 11580
rect 28626 11568 28632 11620
rect 28684 11568 28690 11620
rect 28994 11568 29000 11620
rect 29052 11608 29058 11620
rect 29362 11608 29368 11620
rect 29052 11580 29368 11608
rect 29052 11568 29058 11580
rect 29362 11568 29368 11580
rect 29420 11568 29426 11620
rect 36078 11608 36084 11620
rect 36039 11580 36084 11608
rect 36078 11568 36084 11580
rect 36136 11568 36142 11620
rect 20864 11512 24256 11540
rect 24673 11543 24731 11549
rect 20864 11500 20870 11512
rect 24673 11509 24685 11543
rect 24719 11540 24731 11543
rect 25038 11540 25044 11552
rect 24719 11512 25044 11540
rect 24719 11509 24731 11512
rect 24673 11503 24731 11509
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 25222 11540 25228 11552
rect 25183 11512 25228 11540
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 25590 11500 25596 11552
rect 25648 11540 25654 11552
rect 29181 11543 29239 11549
rect 29181 11540 29193 11543
rect 25648 11512 29193 11540
rect 25648 11500 25654 11512
rect 29181 11509 29193 11512
rect 29227 11509 29239 11543
rect 29181 11503 29239 11509
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 31481 11543 31539 11549
rect 31481 11540 31493 11543
rect 30156 11512 31493 11540
rect 30156 11500 30162 11512
rect 31481 11509 31493 11512
rect 31527 11540 31539 11543
rect 31662 11540 31668 11552
rect 31527 11512 31668 11540
rect 31527 11509 31539 11512
rect 31481 11503 31539 11509
rect 31662 11500 31668 11512
rect 31720 11500 31726 11552
rect 1104 11450 36892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36892 11450
rect 1104 11376 36892 11398
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 2556 11308 9505 11336
rect 2556 11296 2562 11308
rect 9493 11305 9505 11308
rect 9539 11336 9551 11339
rect 9858 11336 9864 11348
rect 9539 11308 9864 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 13906 11336 13912 11348
rect 10468 11308 13912 11336
rect 10468 11296 10474 11308
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 14553 11339 14611 11345
rect 14553 11305 14565 11339
rect 14599 11336 14611 11339
rect 16574 11336 16580 11348
rect 14599 11308 16580 11336
rect 14599 11305 14611 11308
rect 14553 11299 14611 11305
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 18046 11336 18052 11348
rect 17236 11308 18052 11336
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 11054 11268 11060 11280
rect 10744 11240 11060 11268
rect 10744 11228 10750 11240
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11330 11268 11336 11280
rect 11291 11240 11336 11268
rect 11330 11228 11336 11240
rect 11388 11268 11394 11280
rect 12066 11268 12072 11280
rect 11388 11240 12072 11268
rect 11388 11228 11394 11240
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 12253 11271 12311 11277
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12299 11240 15332 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 10183 11172 10793 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 10781 11169 10793 11172
rect 10827 11200 10839 11203
rect 11882 11200 11888 11212
rect 10827 11172 11888 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 11882 11160 11888 11172
rect 11940 11200 11946 11212
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 11940 11172 12909 11200
rect 11940 11160 11946 11172
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 13262 11200 13268 11212
rect 13223 11172 13268 11200
rect 12897 11163 12955 11169
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 14182 11160 14188 11212
rect 14240 11200 14246 11212
rect 15194 11200 15200 11212
rect 14240 11172 15200 11200
rect 14240 11160 14246 11172
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15304 11200 15332 11240
rect 16574 11200 16580 11212
rect 15304 11172 16580 11200
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 17126 11200 17132 11212
rect 16715 11172 17132 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 10042 11132 10048 11144
rect 10003 11104 10048 11132
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11132 12403 11135
rect 12618 11132 12624 11144
rect 12391 11104 12624 11132
rect 12391 11101 12403 11104
rect 12345 11095 12403 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13688 11104 14473 11132
rect 13688 11092 13694 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 7926 11064 7932 11076
rect 7887 11036 7932 11064
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 8573 11067 8631 11073
rect 8076 11036 8121 11064
rect 8076 11024 8082 11036
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9674 11064 9680 11076
rect 8619 11036 9680 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 9674 11024 9680 11036
rect 9732 11064 9738 11076
rect 9732 11036 10824 11064
rect 9732 11024 9738 11036
rect 10796 10996 10824 11036
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 12250 11064 12256 11076
rect 10928 11036 10973 11064
rect 11072 11036 12256 11064
rect 10928 11024 10934 11036
rect 11072 10996 11100 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12986 11064 12992 11076
rect 12947 11036 12992 11064
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 14476 11064 14504 11095
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17000 11104 17045 11132
rect 17000 11092 17006 11104
rect 17236 11064 17264 11308
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 20438 11336 20444 11348
rect 18187 11308 20444 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 25317 11339 25375 11345
rect 25317 11336 25329 11339
rect 23256 11308 25329 11336
rect 23256 11296 23262 11308
rect 25317 11305 25329 11308
rect 25363 11305 25375 11339
rect 25317 11299 25375 11305
rect 25590 11296 25596 11348
rect 25648 11336 25654 11348
rect 26605 11339 26663 11345
rect 26605 11336 26617 11339
rect 25648 11308 26617 11336
rect 25648 11296 25654 11308
rect 26605 11305 26617 11308
rect 26651 11305 26663 11339
rect 27890 11336 27896 11348
rect 27851 11308 27896 11336
rect 26605 11299 26663 11305
rect 27890 11296 27896 11308
rect 27948 11296 27954 11348
rect 29822 11336 29828 11348
rect 28000 11308 29132 11336
rect 29783 11308 29828 11336
rect 17494 11228 17500 11280
rect 17552 11268 17558 11280
rect 17770 11268 17776 11280
rect 17552 11240 17776 11268
rect 17552 11228 17558 11240
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 18230 11228 18236 11280
rect 18288 11268 18294 11280
rect 18785 11271 18843 11277
rect 18785 11268 18797 11271
rect 18288 11240 18797 11268
rect 18288 11228 18294 11240
rect 18785 11237 18797 11240
rect 18831 11237 18843 11271
rect 18785 11231 18843 11237
rect 21453 11271 21511 11277
rect 21453 11237 21465 11271
rect 21499 11268 21511 11271
rect 21634 11268 21640 11280
rect 21499 11240 21640 11268
rect 21499 11237 21511 11240
rect 21453 11231 21511 11237
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 23290 11228 23296 11280
rect 23348 11268 23354 11280
rect 25961 11271 26019 11277
rect 25961 11268 25973 11271
rect 23348 11240 25973 11268
rect 23348 11228 23354 11240
rect 25961 11237 25973 11240
rect 26007 11237 26019 11271
rect 25961 11231 26019 11237
rect 27338 11228 27344 11280
rect 27396 11268 27402 11280
rect 28000 11268 28028 11308
rect 27396 11240 28028 11268
rect 27396 11228 27402 11240
rect 28718 11228 28724 11280
rect 28776 11268 28782 11280
rect 28994 11268 29000 11280
rect 28776 11240 29000 11268
rect 28776 11228 28782 11240
rect 28994 11228 29000 11240
rect 29052 11228 29058 11280
rect 29104 11268 29132 11308
rect 29822 11296 29828 11308
rect 29880 11296 29886 11348
rect 30377 11271 30435 11277
rect 30377 11268 30389 11271
rect 29104 11240 30389 11268
rect 30377 11237 30389 11240
rect 30423 11268 30435 11271
rect 30423 11240 31524 11268
rect 30423 11237 30435 11240
rect 30377 11231 30435 11237
rect 19426 11200 19432 11212
rect 18064 11172 19432 11200
rect 17494 11132 17500 11144
rect 17455 11104 17500 11132
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 18064 11141 18092 11172
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19978 11200 19984 11212
rect 19751 11172 19984 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20622 11160 20628 11212
rect 20680 11200 20686 11212
rect 23658 11200 23664 11212
rect 20680 11172 23664 11200
rect 20680 11160 20686 11172
rect 23658 11160 23664 11172
rect 23716 11160 23722 11212
rect 30929 11203 30987 11209
rect 30929 11200 30941 11203
rect 28276 11172 30941 11200
rect 28276 11144 28304 11172
rect 30929 11169 30941 11172
rect 30975 11169 30987 11203
rect 30929 11163 30987 11169
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11101 17647 11135
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17589 11095 17647 11101
rect 17696 11104 18061 11132
rect 14476 11036 15424 11064
rect 16238 11036 17264 11064
rect 10796 10968 11100 10996
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 13354 10996 13360 11008
rect 11756 10968 13360 10996
rect 11756 10956 11762 10968
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 14458 10996 14464 11008
rect 14240 10968 14464 10996
rect 14240 10956 14246 10968
rect 14458 10956 14464 10968
rect 14516 10956 14522 11008
rect 15194 10996 15200 11008
rect 15155 10968 15200 10996
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15396 10996 15424 11036
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17604 11064 17632 11095
rect 17368 11036 17632 11064
rect 17368 11024 17374 11036
rect 17696 10996 17724 11104
rect 18049 11101 18061 11104
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11132 22155 11135
rect 22462 11132 22468 11144
rect 22143 11104 22468 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 17954 11024 17960 11076
rect 18012 11064 18018 11076
rect 18782 11064 18788 11076
rect 18012 11036 18788 11064
rect 18012 11024 18018 11036
rect 18782 11024 18788 11036
rect 18840 11064 18846 11076
rect 18892 11064 18920 11095
rect 22462 11092 22468 11104
rect 22520 11092 22526 11144
rect 22646 11132 22652 11144
rect 22607 11104 22652 11132
rect 22646 11092 22652 11104
rect 22704 11092 22710 11144
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 23385 11135 23443 11141
rect 22796 11104 22841 11132
rect 22796 11092 22802 11104
rect 23385 11101 23397 11135
rect 23431 11132 23443 11135
rect 24029 11135 24087 11141
rect 23431 11104 23520 11132
rect 23431 11101 23443 11104
rect 23385 11095 23443 11101
rect 18840 11036 18920 11064
rect 19981 11067 20039 11073
rect 18840 11024 18846 11036
rect 19981 11033 19993 11067
rect 20027 11064 20039 11067
rect 20027 11036 20392 11064
rect 20027 11033 20039 11036
rect 19981 11027 20039 11033
rect 20364 11008 20392 11036
rect 20714 11024 20720 11076
rect 20772 11024 20778 11076
rect 23293 11067 23351 11073
rect 23293 11064 23305 11067
rect 21284 11036 23305 11064
rect 15396 10968 17724 10996
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 19518 10996 19524 11008
rect 18380 10968 19524 10996
rect 18380 10956 18386 10968
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 20346 10956 20352 11008
rect 20404 10956 20410 11008
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 21284 10996 21312 11036
rect 23293 11033 23305 11036
rect 23339 11033 23351 11067
rect 23293 11027 23351 11033
rect 21048 10968 21312 10996
rect 21048 10956 21054 10968
rect 21542 10956 21548 11008
rect 21600 10996 21606 11008
rect 22005 10999 22063 11005
rect 22005 10996 22017 10999
rect 21600 10968 22017 10996
rect 21600 10956 21606 10968
rect 22005 10965 22017 10968
rect 22051 10965 22063 10999
rect 23492 10996 23520 11104
rect 24029 11101 24041 11135
rect 24075 11132 24087 11135
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 24075 11104 24777 11132
rect 24075 11101 24087 11104
rect 24029 11095 24087 11101
rect 24765 11101 24777 11104
rect 24811 11132 24823 11135
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 24811 11104 25421 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 25409 11101 25421 11104
rect 25455 11132 25467 11135
rect 25774 11132 25780 11144
rect 25455 11104 25780 11132
rect 25455 11101 25467 11104
rect 25409 11095 25467 11101
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 26053 11135 26111 11141
rect 26053 11101 26065 11135
rect 26099 11101 26111 11135
rect 26694 11132 26700 11144
rect 26655 11104 26700 11132
rect 26053 11095 26111 11101
rect 23566 11024 23572 11076
rect 23624 11064 23630 11076
rect 23937 11067 23995 11073
rect 23937 11064 23949 11067
rect 23624 11036 23949 11064
rect 23624 11024 23630 11036
rect 23937 11033 23949 11036
rect 23983 11033 23995 11067
rect 24670 11064 24676 11076
rect 24631 11036 24676 11064
rect 23937 11027 23995 11033
rect 24670 11024 24676 11036
rect 24728 11024 24734 11076
rect 26068 11064 26096 11095
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 27338 11132 27344 11144
rect 27299 11104 27344 11132
rect 27338 11092 27344 11104
rect 27396 11092 27402 11144
rect 27801 11135 27859 11141
rect 27801 11101 27813 11135
rect 27847 11132 27859 11135
rect 28258 11132 28264 11144
rect 27847 11104 28264 11132
rect 27847 11101 27859 11104
rect 27801 11095 27859 11101
rect 28258 11092 28264 11104
rect 28316 11092 28322 11144
rect 28534 11132 28540 11144
rect 28495 11104 28540 11132
rect 28534 11092 28540 11104
rect 28592 11092 28598 11144
rect 28626 11092 28632 11144
rect 28684 11132 28690 11144
rect 29178 11132 29184 11144
rect 28684 11104 28729 11132
rect 29139 11104 29184 11132
rect 28684 11092 28690 11104
rect 29178 11092 29184 11104
rect 29236 11092 29242 11144
rect 29546 11092 29552 11144
rect 29604 11132 29610 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29604 11104 29745 11132
rect 29604 11092 29610 11104
rect 29733 11101 29745 11104
rect 29779 11132 29791 11135
rect 30098 11132 30104 11144
rect 29779 11104 30104 11132
rect 29779 11101 29791 11104
rect 29733 11095 29791 11101
rect 30098 11092 30104 11104
rect 30156 11092 30162 11144
rect 31496 11134 31524 11240
rect 31496 11106 31616 11134
rect 28442 11064 28448 11076
rect 24780 11036 28448 11064
rect 24210 10996 24216 11008
rect 23492 10968 24216 10996
rect 22005 10959 22063 10965
rect 24210 10956 24216 10968
rect 24268 10996 24274 11008
rect 24780 10996 24808 11036
rect 28442 11024 28448 11036
rect 28500 11024 28506 11076
rect 31481 11067 31539 11073
rect 31481 11064 31493 11067
rect 28966 11036 31493 11064
rect 24268 10968 24808 10996
rect 24268 10956 24274 10968
rect 24946 10956 24952 11008
rect 25004 10996 25010 11008
rect 26142 10996 26148 11008
rect 25004 10968 26148 10996
rect 25004 10956 25010 10968
rect 26142 10956 26148 10968
rect 26200 10956 26206 11008
rect 27246 10996 27252 11008
rect 27207 10968 27252 10996
rect 27246 10956 27252 10968
rect 27304 10956 27310 11008
rect 28626 10956 28632 11008
rect 28684 10996 28690 11008
rect 28966 10996 28994 11036
rect 31481 11033 31493 11036
rect 31527 11033 31539 11067
rect 31588 11064 31616 11106
rect 31662 11092 31668 11144
rect 31720 11132 31726 11144
rect 32033 11135 32091 11141
rect 32033 11132 32045 11135
rect 31720 11104 32045 11132
rect 31720 11092 31726 11104
rect 32033 11101 32045 11104
rect 32079 11101 32091 11135
rect 32033 11095 32091 11101
rect 35526 11064 35532 11076
rect 31588 11036 35532 11064
rect 31481 11027 31539 11033
rect 35526 11024 35532 11036
rect 35584 11024 35590 11076
rect 28684 10968 28994 10996
rect 28684 10956 28690 10968
rect 1104 10906 36892 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 36892 10906
rect 1104 10832 36892 10854
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 7984 10764 8033 10792
rect 7984 10752 7990 10764
rect 8021 10761 8033 10764
rect 8067 10761 8079 10795
rect 8754 10792 8760 10804
rect 8715 10764 8760 10792
rect 8021 10755 8079 10761
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 13078 10792 13084 10804
rect 11164 10764 13084 10792
rect 10502 10724 10508 10736
rect 10463 10696 10508 10724
rect 10502 10684 10508 10696
rect 10560 10684 10566 10736
rect 1854 10656 1860 10668
rect 1815 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 10134 10656 10140 10668
rect 8895 10628 10140 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 11164 10665 11192 10764
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 13173 10795 13231 10801
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 16298 10792 16304 10804
rect 13219 10764 16304 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 19334 10792 19340 10804
rect 16991 10764 19340 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 21266 10792 21272 10804
rect 20220 10764 21272 10792
rect 20220 10752 20226 10764
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 21358 10752 21364 10804
rect 21416 10792 21422 10804
rect 24946 10792 24952 10804
rect 21416 10764 24952 10792
rect 21416 10752 21422 10764
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 25133 10795 25191 10801
rect 25133 10761 25145 10795
rect 25179 10792 25191 10795
rect 25498 10792 25504 10804
rect 25179 10764 25504 10792
rect 25179 10761 25191 10764
rect 25133 10755 25191 10761
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 26050 10752 26056 10804
rect 26108 10792 26114 10804
rect 26421 10795 26479 10801
rect 26421 10792 26433 10795
rect 26108 10764 26433 10792
rect 26108 10752 26114 10764
rect 26421 10761 26433 10764
rect 26467 10761 26479 10795
rect 26421 10755 26479 10761
rect 27249 10795 27307 10801
rect 27249 10761 27261 10795
rect 27295 10792 27307 10795
rect 27982 10792 27988 10804
rect 27295 10764 27988 10792
rect 27295 10761 27307 10764
rect 27249 10755 27307 10761
rect 27982 10752 27988 10764
rect 28040 10752 28046 10804
rect 35526 10792 35532 10804
rect 35487 10764 35532 10792
rect 35526 10752 35532 10764
rect 35584 10752 35590 10804
rect 11882 10684 11888 10736
rect 11940 10724 11946 10736
rect 14737 10727 14795 10733
rect 14737 10724 14749 10727
rect 11940 10696 14749 10724
rect 11940 10684 11946 10696
rect 14737 10693 14749 10696
rect 14783 10693 14795 10727
rect 14737 10687 14795 10693
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 14884 10696 15226 10724
rect 14884 10684 14890 10696
rect 17218 10684 17224 10736
rect 17276 10724 17282 10736
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 17276 10696 17785 10724
rect 17276 10684 17282 10696
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 19242 10724 19248 10736
rect 18998 10696 19248 10724
rect 17773 10687 17831 10693
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 19720 10696 19993 10724
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 11149 10619 11207 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12952 10628 13093 10656
rect 12952 10616 12958 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10625 13875 10659
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 13817 10619 13875 10625
rect 15948 10628 16865 10656
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11238 10588 11244 10600
rect 11103 10560 11244 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 11974 10588 11980 10600
rect 11935 10560 11980 10588
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 9858 10480 9864 10532
rect 9916 10520 9922 10532
rect 9953 10523 10011 10529
rect 9953 10520 9965 10523
rect 9916 10492 9965 10520
rect 9916 10480 9922 10492
rect 9953 10489 9965 10492
rect 9999 10520 10011 10523
rect 13832 10520 13860 10619
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14458 10588 14464 10600
rect 14056 10560 14101 10588
rect 14419 10560 14464 10588
rect 14056 10548 14062 10560
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 9999 10492 13860 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 9398 10452 9404 10464
rect 9359 10424 9404 10452
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12526 10452 12532 10464
rect 12483 10424 12532 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 15948 10452 15976 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 19720 10656 19748 10696
rect 19981 10693 19993 10696
rect 20027 10724 20039 10727
rect 20254 10724 20260 10736
rect 20027 10696 20260 10724
rect 20027 10693 20039 10696
rect 19981 10687 20039 10693
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 22002 10724 22008 10736
rect 21206 10696 22008 10724
rect 22002 10684 22008 10696
rect 22060 10684 22066 10736
rect 22738 10684 22744 10736
rect 22796 10724 22802 10736
rect 22796 10696 22876 10724
rect 22796 10684 22802 10696
rect 17000 10628 17540 10656
rect 17000 10616 17006 10628
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16960 10588 16988 10616
rect 17512 10597 17540 10628
rect 19260 10628 19748 10656
rect 19260 10597 19288 10628
rect 21266 10616 21272 10668
rect 21324 10656 21330 10668
rect 22848 10665 22876 10696
rect 23106 10684 23112 10736
rect 23164 10724 23170 10736
rect 23658 10724 23664 10736
rect 23164 10696 23664 10724
rect 23164 10684 23170 10696
rect 23658 10684 23664 10696
rect 23716 10684 23722 10736
rect 25406 10724 25412 10736
rect 24886 10696 25412 10724
rect 25406 10684 25412 10696
rect 25464 10684 25470 10736
rect 26694 10724 26700 10736
rect 25884 10696 26700 10724
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 21324 10628 22201 10656
rect 21324 10616 21330 10628
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 22922 10616 22928 10668
rect 22980 10656 22986 10668
rect 25884 10665 25912 10696
rect 26694 10684 26700 10696
rect 26752 10684 26758 10736
rect 28074 10724 28080 10736
rect 28035 10696 28080 10724
rect 28074 10684 28080 10696
rect 28132 10684 28138 10736
rect 28629 10727 28687 10733
rect 28629 10693 28641 10727
rect 28675 10724 28687 10727
rect 30285 10727 30343 10733
rect 30285 10724 30297 10727
rect 28675 10696 30297 10724
rect 28675 10693 28687 10696
rect 28629 10687 28687 10693
rect 30285 10693 30297 10696
rect 30331 10693 30343 10727
rect 35544 10724 35572 10752
rect 35544 10696 36124 10724
rect 30285 10687 30343 10693
rect 23385 10659 23443 10665
rect 23385 10656 23397 10659
rect 22980 10628 23397 10656
rect 22980 10616 22986 10628
rect 23385 10625 23397 10628
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 25869 10659 25927 10665
rect 25869 10625 25881 10659
rect 25915 10625 25927 10659
rect 25869 10619 25927 10625
rect 26329 10659 26387 10665
rect 26329 10625 26341 10659
rect 26375 10656 26387 10659
rect 26418 10656 26424 10668
rect 26375 10628 26424 10656
rect 26375 10625 26387 10628
rect 26329 10619 26387 10625
rect 26418 10616 26424 10628
rect 26476 10616 26482 10668
rect 26878 10616 26884 10668
rect 26936 10656 26942 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 26936 10628 27169 10656
rect 26936 10616 26942 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 29178 10616 29184 10668
rect 29236 10656 29242 10668
rect 29733 10659 29791 10665
rect 29733 10656 29745 10659
rect 29236 10628 29745 10656
rect 29236 10616 29242 10628
rect 29733 10625 29745 10628
rect 29779 10656 29791 10659
rect 30006 10656 30012 10668
rect 29779 10628 30012 10656
rect 29779 10625 29791 10628
rect 29733 10619 29791 10625
rect 30006 10616 30012 10628
rect 30064 10616 30070 10668
rect 30190 10616 30196 10668
rect 30248 10656 30254 10668
rect 30377 10659 30435 10665
rect 30377 10656 30389 10659
rect 30248 10628 30389 10656
rect 30248 10616 30254 10628
rect 30377 10625 30389 10628
rect 30423 10625 30435 10659
rect 30377 10619 30435 10625
rect 31021 10659 31079 10665
rect 31021 10625 31033 10659
rect 31067 10656 31079 10659
rect 35986 10656 35992 10668
rect 31067 10628 35992 10656
rect 31067 10625 31079 10628
rect 31021 10619 31079 10625
rect 16632 10560 16988 10588
rect 17497 10591 17555 10597
rect 16632 10548 16638 10560
rect 17497 10557 17509 10591
rect 17543 10557 17555 10591
rect 19245 10591 19303 10597
rect 17497 10551 17555 10557
rect 17604 10560 18828 10588
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 17604 10520 17632 10560
rect 17184 10492 17632 10520
rect 18800 10520 18828 10560
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 19610 10520 19616 10532
rect 18800 10492 19616 10520
rect 17184 10480 17190 10492
rect 19610 10480 19616 10492
rect 19668 10480 19674 10532
rect 13688 10424 15976 10452
rect 13688 10412 13694 10424
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 16080 10424 16221 10452
rect 16080 10412 16086 10424
rect 16209 10421 16221 10424
rect 16255 10421 16267 10455
rect 16209 10415 16267 10421
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 17954 10452 17960 10464
rect 16356 10424 17960 10452
rect 16356 10412 16362 10424
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 19720 10452 19748 10551
rect 20438 10548 20444 10600
rect 20496 10588 20502 10600
rect 22741 10591 22799 10597
rect 22741 10588 22753 10591
rect 20496 10560 22753 10588
rect 20496 10548 20502 10560
rect 22741 10557 22753 10560
rect 22787 10557 22799 10591
rect 27246 10588 27252 10600
rect 22741 10551 22799 10557
rect 23492 10560 27252 10588
rect 21082 10480 21088 10532
rect 21140 10520 21146 10532
rect 23492 10520 23520 10560
rect 27246 10548 27252 10560
rect 27304 10548 27310 10600
rect 28718 10588 28724 10600
rect 28679 10560 28724 10588
rect 28718 10548 28724 10560
rect 28776 10548 28782 10600
rect 29457 10591 29515 10597
rect 29457 10557 29469 10591
rect 29503 10557 29515 10591
rect 30392 10588 30420 10619
rect 35986 10616 35992 10628
rect 36044 10616 36050 10668
rect 36096 10665 36124 10696
rect 36081 10659 36139 10665
rect 36081 10625 36093 10659
rect 36127 10625 36139 10659
rect 36081 10619 36139 10625
rect 31481 10591 31539 10597
rect 31481 10588 31493 10591
rect 30392 10560 31493 10588
rect 29457 10551 29515 10557
rect 31481 10557 31493 10560
rect 31527 10557 31539 10591
rect 31481 10551 31539 10557
rect 25777 10523 25835 10529
rect 25777 10520 25789 10523
rect 21140 10492 23520 10520
rect 24688 10492 25789 10520
rect 21140 10480 21146 10492
rect 19978 10452 19984 10464
rect 19720 10424 19984 10452
rect 19978 10412 19984 10424
rect 20036 10452 20042 10464
rect 20530 10452 20536 10464
rect 20036 10424 20536 10452
rect 20036 10412 20042 10424
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 21358 10412 21364 10464
rect 21416 10452 21422 10464
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 21416 10424 21465 10452
rect 21416 10412 21422 10424
rect 21453 10421 21465 10424
rect 21499 10421 21511 10455
rect 21453 10415 21511 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22152 10424 22197 10452
rect 22152 10412 22158 10424
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 24688 10452 24716 10492
rect 25777 10489 25789 10492
rect 25823 10489 25835 10523
rect 25777 10483 25835 10489
rect 26694 10480 26700 10532
rect 26752 10520 26758 10532
rect 27154 10520 27160 10532
rect 26752 10492 27160 10520
rect 26752 10480 26758 10492
rect 27154 10480 27160 10492
rect 27212 10480 27218 10532
rect 23440 10424 24716 10452
rect 23440 10412 23446 10424
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 29472 10452 29500 10551
rect 24820 10424 29500 10452
rect 24820 10412 24826 10424
rect 30374 10412 30380 10464
rect 30432 10452 30438 10464
rect 30929 10455 30987 10461
rect 30929 10452 30941 10455
rect 30432 10424 30941 10452
rect 30432 10412 30438 10424
rect 30929 10421 30941 10424
rect 30975 10421 30987 10455
rect 36262 10452 36268 10464
rect 36223 10424 36268 10452
rect 30929 10415 30987 10421
rect 36262 10412 36268 10424
rect 36320 10412 36326 10464
rect 1104 10362 36892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36892 10362
rect 1104 10288 36892 10310
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 9456 10220 10333 10248
rect 9456 10208 9462 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10321 10211 10379 10217
rect 11701 10251 11759 10257
rect 11701 10217 11713 10251
rect 11747 10248 11759 10251
rect 11974 10248 11980 10260
rect 11747 10220 11980 10248
rect 11747 10217 11759 10220
rect 11701 10211 11759 10217
rect 10336 10180 10364 10211
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 12986 10248 12992 10260
rect 12391 10220 12992 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 15562 10248 15568 10260
rect 13679 10220 15568 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 18322 10248 18328 10260
rect 16080 10220 18328 10248
rect 16080 10208 16086 10220
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10217 18843 10251
rect 18785 10211 18843 10217
rect 12894 10180 12900 10192
rect 10336 10152 12900 10180
rect 12894 10140 12900 10152
rect 12952 10180 12958 10192
rect 13538 10180 13544 10192
rect 12952 10152 13544 10180
rect 12952 10140 12958 10152
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 16758 10140 16764 10192
rect 16816 10180 16822 10192
rect 17678 10180 17684 10192
rect 16816 10152 17684 10180
rect 16816 10140 16822 10152
rect 17678 10140 17684 10152
rect 17736 10140 17742 10192
rect 18046 10140 18052 10192
rect 18104 10180 18110 10192
rect 18800 10180 18828 10211
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 21450 10248 21456 10260
rect 18932 10220 21456 10248
rect 18932 10208 18938 10220
rect 21450 10208 21456 10220
rect 21508 10208 21514 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 21876 10220 23121 10248
rect 21876 10208 21882 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 25682 10248 25688 10260
rect 23109 10211 23167 10217
rect 23400 10220 25688 10248
rect 18104 10152 18828 10180
rect 18104 10140 18110 10152
rect 19334 10140 19340 10192
rect 19392 10180 19398 10192
rect 20254 10180 20260 10192
rect 19392 10152 20260 10180
rect 19392 10140 19398 10152
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 21910 10140 21916 10192
rect 21968 10180 21974 10192
rect 21968 10152 22094 10180
rect 21968 10140 21974 10152
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 13556 10112 13584 10140
rect 9824 10084 12296 10112
rect 13556 10084 14504 10112
rect 9824 10072 9830 10084
rect 12268 10056 12296 10084
rect 10873 10047 10931 10053
rect 10873 10044 10885 10047
rect 8496 10016 10885 10044
rect 1762 9936 1768 9988
rect 1820 9976 1826 9988
rect 2682 9976 2688 9988
rect 1820 9948 2688 9976
rect 1820 9936 1826 9948
rect 2682 9936 2688 9948
rect 2740 9976 2746 9988
rect 8496 9985 8524 10016
rect 10873 10013 10885 10016
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11882 10044 11888 10056
rect 11655 10016 11888 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 12250 10044 12256 10056
rect 12163 10016 12256 10044
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10044 12955 10047
rect 13446 10044 13452 10056
rect 12943 10016 13452 10044
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 8481 9979 8539 9985
rect 8481 9976 8493 9979
rect 2740 9948 8493 9976
rect 2740 9936 2746 9948
rect 8481 9945 8493 9948
rect 8527 9945 8539 9979
rect 8481 9939 8539 9945
rect 9861 9979 9919 9985
rect 9861 9945 9873 9979
rect 9907 9976 9919 9979
rect 9907 9948 12434 9976
rect 9907 9945 9919 9948
rect 9861 9939 9919 9945
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9766 9908 9772 9920
rect 9355 9880 9772 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10965 9911 11023 9917
rect 10965 9877 10977 9911
rect 11011 9908 11023 9911
rect 12158 9908 12164 9920
rect 11011 9880 12164 9908
rect 11011 9877 11023 9880
rect 10965 9871 11023 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12406 9908 12434 9948
rect 12912 9908 12940 10007
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14366 10044 14372 10056
rect 13771 10016 14372 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14476 10053 14504 10084
rect 14642 10072 14648 10124
rect 14700 10072 14706 10124
rect 15105 10115 15163 10121
rect 15105 10081 15117 10115
rect 15151 10112 15163 10115
rect 16574 10112 16580 10124
rect 15151 10084 16580 10112
rect 15151 10081 15163 10084
rect 15105 10075 15163 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 17586 10112 17592 10124
rect 17175 10084 17592 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 21542 10112 21548 10124
rect 17972 10084 21548 10112
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9976 13047 9979
rect 14660 9976 14688 10072
rect 17972 10044 18000 10084
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 22066 10112 22094 10152
rect 22738 10140 22744 10192
rect 22796 10180 22802 10192
rect 23400 10180 23428 10220
rect 25682 10208 25688 10220
rect 25740 10208 25746 10260
rect 27157 10251 27215 10257
rect 27157 10217 27169 10251
rect 27203 10248 27215 10251
rect 27614 10248 27620 10260
rect 27203 10220 27620 10248
rect 27203 10217 27215 10220
rect 27157 10211 27215 10217
rect 27614 10208 27620 10220
rect 27672 10208 27678 10260
rect 22796 10152 23428 10180
rect 22796 10140 22802 10152
rect 23934 10140 23940 10192
rect 23992 10180 23998 10192
rect 24854 10180 24860 10192
rect 23992 10152 24860 10180
rect 23992 10140 23998 10152
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 28718 10140 28724 10192
rect 28776 10180 28782 10192
rect 30374 10180 30380 10192
rect 28776 10152 30380 10180
rect 28776 10140 28782 10152
rect 30374 10140 30380 10152
rect 30432 10140 30438 10192
rect 30190 10112 30196 10124
rect 22066 10084 30196 10112
rect 30190 10072 30196 10084
rect 30248 10072 30254 10124
rect 16514 10016 18000 10044
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 18104 10016 18149 10044
rect 18104 10004 18110 10016
rect 18782 10004 18788 10056
rect 18840 10044 18846 10056
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 18840 10016 18889 10044
rect 18840 10004 18846 10016
rect 18877 10013 18889 10016
rect 18923 10044 18935 10047
rect 19889 10047 19947 10053
rect 19889 10044 19901 10047
rect 18923 10016 19901 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19889 10013 19901 10016
rect 19935 10044 19947 10047
rect 20162 10044 20168 10056
rect 19935 10016 20168 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 20530 10044 20536 10056
rect 20491 10016 20536 10044
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 21910 10004 21916 10056
rect 21968 10004 21974 10056
rect 23201 10047 23259 10053
rect 23201 10013 23213 10047
rect 23247 10044 23259 10047
rect 23845 10047 23903 10053
rect 23845 10044 23857 10047
rect 23247 10016 23857 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 23845 10013 23857 10016
rect 23891 10044 23903 10047
rect 24210 10044 24216 10056
rect 23891 10016 24216 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24210 10004 24216 10016
rect 24268 10004 24274 10056
rect 24670 10044 24676 10056
rect 24504 10016 24676 10044
rect 15378 9976 15384 9988
rect 13035 9948 14688 9976
rect 15339 9948 15384 9976
rect 13035 9945 13047 9948
rect 12989 9939 13047 9945
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17310 9976 17316 9988
rect 16908 9948 17316 9976
rect 16908 9936 16914 9948
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 18322 9936 18328 9988
rect 18380 9976 18386 9988
rect 20714 9976 20720 9988
rect 18380 9948 20720 9976
rect 18380 9936 18386 9948
rect 20714 9936 20720 9948
rect 20772 9936 20778 9988
rect 20806 9936 20812 9988
rect 20864 9976 20870 9988
rect 22557 9979 22615 9985
rect 20864 9948 20909 9976
rect 20864 9936 20870 9948
rect 22557 9945 22569 9979
rect 22603 9976 22615 9979
rect 24504 9976 24532 10016
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 26602 10004 26608 10056
rect 26660 10044 26666 10056
rect 27062 10044 27068 10056
rect 26660 10016 26705 10044
rect 27023 10016 27068 10044
rect 26660 10004 26666 10016
rect 27062 10004 27068 10016
rect 27120 10004 27126 10056
rect 27890 10044 27896 10056
rect 27851 10016 27896 10044
rect 27890 10004 27896 10016
rect 27948 10004 27954 10056
rect 29178 10044 29184 10056
rect 29139 10016 29184 10044
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 30926 10004 30932 10056
rect 30984 10044 30990 10056
rect 31113 10047 31171 10053
rect 31113 10044 31125 10047
rect 30984 10016 31125 10044
rect 30984 10004 30990 10016
rect 31113 10013 31125 10016
rect 31159 10044 31171 10047
rect 31573 10047 31631 10053
rect 31573 10044 31585 10047
rect 31159 10016 31585 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 31573 10013 31585 10016
rect 31619 10013 31631 10047
rect 31573 10007 31631 10013
rect 22603 9948 24532 9976
rect 24581 9979 24639 9985
rect 22603 9945 22615 9948
rect 22557 9939 22615 9945
rect 24581 9945 24593 9979
rect 24627 9976 24639 9979
rect 24854 9976 24860 9988
rect 24627 9948 24860 9976
rect 24627 9945 24639 9948
rect 24581 9939 24639 9945
rect 14550 9908 14556 9920
rect 12406 9880 12940 9908
rect 14511 9880 14556 9908
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 18046 9908 18052 9920
rect 17644 9880 18052 9908
rect 17644 9868 17650 9880
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 18966 9908 18972 9920
rect 18187 9880 18972 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 19981 9911 20039 9917
rect 19981 9877 19993 9911
rect 20027 9908 20039 9911
rect 21082 9908 21088 9920
rect 20027 9880 21088 9908
rect 20027 9877 20039 9880
rect 19981 9871 20039 9877
rect 21082 9868 21088 9880
rect 21140 9868 21146 9920
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 22572 9908 22600 9939
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 26329 9979 26387 9985
rect 25898 9948 26280 9976
rect 23750 9908 23756 9920
rect 21508 9880 22600 9908
rect 23711 9880 23756 9908
rect 21508 9868 21514 9880
rect 23750 9868 23756 9880
rect 23808 9868 23814 9920
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24762 9908 24768 9920
rect 24084 9880 24768 9908
rect 24084 9868 24090 9880
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 26252 9908 26280 9948
rect 26329 9945 26341 9979
rect 26375 9976 26387 9979
rect 27614 9976 27620 9988
rect 26375 9948 27620 9976
rect 26375 9945 26387 9948
rect 26329 9939 26387 9945
rect 27614 9936 27620 9948
rect 27672 9976 27678 9988
rect 28350 9976 28356 9988
rect 27672 9948 28356 9976
rect 27672 9936 27678 9948
rect 28350 9936 28356 9948
rect 28408 9936 28414 9988
rect 28718 9936 28724 9988
rect 28776 9976 28782 9988
rect 28905 9979 28963 9985
rect 28905 9976 28917 9979
rect 28776 9948 28917 9976
rect 28776 9936 28782 9948
rect 28905 9945 28917 9948
rect 28951 9945 28963 9979
rect 28905 9939 28963 9945
rect 29086 9936 29092 9988
rect 29144 9976 29150 9988
rect 29733 9979 29791 9985
rect 29733 9976 29745 9979
rect 29144 9948 29745 9976
rect 29144 9936 29150 9948
rect 29733 9945 29745 9948
rect 29779 9976 29791 9979
rect 30190 9976 30196 9988
rect 29779 9948 30196 9976
rect 29779 9945 29791 9948
rect 29733 9939 29791 9945
rect 30190 9936 30196 9948
rect 30248 9936 30254 9988
rect 30285 9979 30343 9985
rect 30285 9945 30297 9979
rect 30331 9945 30343 9979
rect 30285 9939 30343 9945
rect 27706 9908 27712 9920
rect 26252 9880 27712 9908
rect 27706 9868 27712 9880
rect 27764 9868 27770 9920
rect 27801 9911 27859 9917
rect 27801 9877 27813 9911
rect 27847 9908 27859 9911
rect 27982 9908 27988 9920
rect 27847 9880 27988 9908
rect 27847 9877 27859 9880
rect 27801 9871 27859 9877
rect 27982 9868 27988 9880
rect 28040 9868 28046 9920
rect 30300 9908 30328 9939
rect 30374 9936 30380 9988
rect 30432 9976 30438 9988
rect 30432 9948 30477 9976
rect 30432 9936 30438 9948
rect 31021 9911 31079 9917
rect 31021 9908 31033 9911
rect 30300 9880 31033 9908
rect 31021 9877 31033 9880
rect 31067 9877 31079 9911
rect 31021 9871 31079 9877
rect 1104 9818 36892 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 36892 9818
rect 1104 9744 36892 9766
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 15654 9704 15660 9716
rect 13136 9676 15660 9704
rect 13136 9664 13142 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 32030 9704 32036 9716
rect 15896 9676 32036 9704
rect 15896 9664 15902 9676
rect 32030 9664 32036 9676
rect 32088 9664 32094 9716
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 11422 9636 11428 9648
rect 10643 9608 11428 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 12253 9639 12311 9645
rect 12253 9636 12265 9639
rect 12032 9608 12265 9636
rect 12032 9596 12038 9608
rect 12253 9605 12265 9608
rect 12299 9605 12311 9639
rect 12253 9599 12311 9605
rect 12345 9639 12403 9645
rect 12345 9605 12357 9639
rect 12391 9636 12403 9639
rect 12526 9636 12532 9648
rect 12391 9608 12532 9636
rect 12391 9605 12403 9608
rect 12345 9599 12403 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 13265 9639 13323 9645
rect 13265 9605 13277 9639
rect 13311 9636 13323 9639
rect 14734 9636 14740 9648
rect 13311 9608 14740 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 16945 9639 17003 9645
rect 15594 9608 16896 9636
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11698 9568 11704 9580
rect 11195 9540 11704 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9568 13875 9571
rect 13998 9568 14004 9580
rect 13863 9540 14004 9568
rect 13863 9537 13875 9540
rect 13817 9531 13875 9537
rect 10502 9500 10508 9512
rect 10415 9472 10508 9500
rect 10502 9460 10508 9472
rect 10560 9500 10566 9512
rect 12069 9503 12127 9509
rect 10560 9472 11928 9500
rect 10560 9460 10566 9472
rect 11900 9432 11928 9472
rect 12069 9469 12081 9503
rect 12115 9500 12127 9503
rect 12158 9500 12164 9512
rect 12115 9472 12164 9500
rect 12115 9469 12127 9472
rect 12069 9463 12127 9469
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 13188 9500 13216 9531
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 16868 9568 16896 9608
rect 16945 9605 16957 9639
rect 16991 9636 17003 9639
rect 17034 9636 17040 9648
rect 16991 9608 17040 9636
rect 16991 9605 17003 9608
rect 16945 9599 17003 9605
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 18138 9596 18144 9648
rect 18196 9596 18202 9648
rect 19429 9639 19487 9645
rect 19429 9605 19441 9639
rect 19475 9636 19487 9639
rect 20346 9636 20352 9648
rect 19475 9608 20352 9636
rect 19475 9605 19487 9608
rect 19429 9599 19487 9605
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 25222 9636 25228 9648
rect 23782 9608 25228 9636
rect 25222 9596 25228 9608
rect 25280 9596 25286 9648
rect 25406 9636 25412 9648
rect 25367 9608 25412 9636
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 25682 9596 25688 9648
rect 25740 9636 25746 9648
rect 29546 9636 29552 9648
rect 25740 9608 25912 9636
rect 25740 9596 25746 9608
rect 17310 9568 17316 9580
rect 16868 9540 17316 9568
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 20162 9528 20168 9580
rect 20220 9568 20226 9580
rect 20441 9571 20499 9577
rect 20441 9568 20453 9571
rect 20220 9540 20453 9568
rect 20220 9528 20226 9540
rect 20441 9537 20453 9540
rect 20487 9537 20499 9571
rect 21085 9571 21143 9577
rect 21085 9568 21097 9571
rect 20441 9531 20499 9537
rect 20732 9540 21097 9568
rect 12308 9472 13216 9500
rect 12308 9460 12314 9472
rect 12710 9432 12716 9444
rect 11900 9404 12716 9432
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 13188 9432 13216 9472
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9500 13967 9503
rect 15286 9500 15292 9512
rect 13955 9472 15292 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15712 9472 16037 9500
rect 15712 9460 15718 9472
rect 16025 9469 16037 9472
rect 16071 9500 16083 9503
rect 16301 9503 16359 9509
rect 16071 9472 16252 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16224 9432 16252 9472
rect 16301 9469 16313 9503
rect 16347 9500 16359 9503
rect 16574 9500 16580 9512
rect 16347 9472 16580 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 16574 9460 16580 9472
rect 16632 9500 16638 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16632 9472 17417 9500
rect 16632 9460 16638 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 17828 9472 20361 9500
rect 17828 9460 17834 9472
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 17034 9432 17040 9444
rect 13188 9404 15056 9432
rect 16224 9404 17040 9432
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10962 9364 10968 9376
rect 9999 9336 10968 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 14553 9367 14611 9373
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 14642 9364 14648 9376
rect 14599 9336 14648 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15028 9364 15056 9404
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 20732 9432 20760 9540
rect 21085 9537 21097 9540
rect 21131 9568 21143 9571
rect 21450 9568 21456 9580
rect 21131 9540 21456 9568
rect 21131 9537 21143 9540
rect 21085 9531 21143 9537
rect 21450 9528 21456 9540
rect 21508 9568 21514 9580
rect 21508 9540 22094 9568
rect 21508 9528 21514 9540
rect 19300 9404 20760 9432
rect 19300 9392 19306 9404
rect 15562 9364 15568 9376
rect 15028 9336 15568 9364
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 17402 9364 17408 9376
rect 15896 9336 17408 9364
rect 15896 9324 15902 9336
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17668 9367 17726 9373
rect 17668 9333 17680 9367
rect 17714 9364 17726 9367
rect 18046 9364 18052 9376
rect 17714 9336 18052 9364
rect 17714 9333 17726 9336
rect 17668 9327 17726 9333
rect 18046 9324 18052 9336
rect 18104 9364 18110 9376
rect 18690 9364 18696 9376
rect 18104 9336 18696 9364
rect 18104 9324 18110 9336
rect 18690 9324 18696 9336
rect 18748 9324 18754 9376
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19978 9364 19984 9376
rect 18932 9336 19984 9364
rect 18932 9324 18938 9336
rect 19978 9324 19984 9336
rect 20036 9364 20042 9376
rect 20346 9364 20352 9376
rect 20036 9336 20352 9364
rect 20036 9324 20042 9336
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20714 9324 20720 9376
rect 20772 9364 20778 9376
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 20772 9336 21005 9364
rect 20772 9324 20778 9336
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 22066 9364 22094 9540
rect 24486 9528 24492 9580
rect 24544 9568 24550 9580
rect 25501 9571 25559 9577
rect 24544 9540 24589 9568
rect 24544 9528 24550 9540
rect 25501 9537 25513 9571
rect 25547 9568 25559 9571
rect 25774 9568 25780 9580
rect 25547 9540 25780 9568
rect 25547 9537 25559 9540
rect 25501 9531 25559 9537
rect 25774 9528 25780 9540
rect 25832 9528 25838 9580
rect 25884 9568 25912 9608
rect 28000 9608 29552 9636
rect 26121 9569 26179 9575
rect 25884 9566 26004 9568
rect 26121 9566 26133 9569
rect 25884 9540 26133 9566
rect 25976 9538 26133 9540
rect 26121 9535 26133 9538
rect 26167 9535 26179 9569
rect 27338 9568 27344 9580
rect 27299 9540 27344 9568
rect 26121 9529 26179 9535
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 27798 9528 27804 9580
rect 27856 9568 27862 9580
rect 28000 9577 28028 9608
rect 29546 9596 29552 9608
rect 29604 9596 29610 9648
rect 29638 9596 29644 9648
rect 29696 9636 29702 9648
rect 30009 9639 30067 9645
rect 30009 9636 30021 9639
rect 29696 9608 30021 9636
rect 29696 9596 29702 9608
rect 30009 9605 30021 9608
rect 30055 9605 30067 9639
rect 30558 9636 30564 9648
rect 30519 9608 30564 9636
rect 30009 9599 30067 9605
rect 30558 9596 30564 9608
rect 30616 9596 30622 9648
rect 30650 9596 30656 9648
rect 30708 9636 30714 9648
rect 30708 9608 30753 9636
rect 30708 9596 30714 9608
rect 27985 9571 28043 9577
rect 27985 9568 27997 9571
rect 27856 9540 27997 9568
rect 27856 9528 27862 9540
rect 27985 9537 27997 9540
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 28629 9571 28687 9577
rect 28629 9537 28641 9571
rect 28675 9537 28687 9571
rect 28629 9531 28687 9537
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 23842 9500 23848 9512
rect 22511 9472 23848 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 23842 9460 23848 9472
rect 23900 9460 23906 9512
rect 24213 9503 24271 9509
rect 24213 9469 24225 9503
rect 24259 9500 24271 9503
rect 24504 9500 24532 9528
rect 26602 9500 26608 9512
rect 24259 9472 24440 9500
rect 24504 9472 26608 9500
rect 24259 9469 24271 9472
rect 24213 9463 24271 9469
rect 24412 9432 24440 9472
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27890 9460 27896 9512
rect 27948 9500 27954 9512
rect 28644 9500 28672 9531
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 29273 9571 29331 9577
rect 29273 9568 29285 9571
rect 29052 9540 29285 9568
rect 29052 9528 29058 9540
rect 29273 9537 29285 9540
rect 29319 9537 29331 9571
rect 29273 9531 29331 9537
rect 35897 9571 35955 9577
rect 35897 9537 35909 9571
rect 35943 9568 35955 9571
rect 35986 9568 35992 9580
rect 35943 9540 35992 9568
rect 35943 9537 35955 9540
rect 35897 9531 35955 9537
rect 35986 9528 35992 9540
rect 36044 9528 36050 9580
rect 27948 9472 28672 9500
rect 27948 9460 27954 9472
rect 26510 9432 26516 9444
rect 24412 9404 26516 9432
rect 26510 9392 26516 9404
rect 26568 9392 26574 9444
rect 27154 9392 27160 9444
rect 27212 9432 27218 9444
rect 29181 9435 29239 9441
rect 29181 9432 29193 9435
rect 27212 9404 29193 9432
rect 27212 9392 27218 9404
rect 29181 9401 29193 9404
rect 29227 9401 29239 9435
rect 29181 9395 29239 9401
rect 24026 9364 24032 9376
rect 22066 9336 24032 9364
rect 20993 9327 21051 9333
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 24210 9324 24216 9376
rect 24268 9364 24274 9376
rect 26053 9367 26111 9373
rect 26053 9364 26065 9367
rect 24268 9336 26065 9364
rect 24268 9324 24274 9336
rect 26053 9333 26065 9336
rect 26099 9333 26111 9367
rect 26053 9327 26111 9333
rect 26234 9324 26240 9376
rect 26292 9364 26298 9376
rect 27249 9367 27307 9373
rect 27249 9364 27261 9367
rect 26292 9336 27261 9364
rect 26292 9324 26298 9336
rect 27249 9333 27261 9336
rect 27295 9333 27307 9367
rect 27249 9327 27307 9333
rect 27798 9324 27804 9376
rect 27856 9364 27862 9376
rect 27893 9367 27951 9373
rect 27893 9364 27905 9367
rect 27856 9336 27905 9364
rect 27856 9324 27862 9336
rect 27893 9333 27905 9336
rect 27939 9333 27951 9367
rect 28534 9364 28540 9376
rect 28495 9336 28540 9364
rect 27893 9327 27951 9333
rect 28534 9324 28540 9336
rect 28592 9324 28598 9376
rect 36078 9364 36084 9376
rect 36039 9336 36084 9364
rect 36078 9324 36084 9336
rect 36136 9324 36142 9376
rect 1104 9274 36892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36892 9274
rect 1104 9200 36892 9222
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 9824 9132 9873 9160
rect 9824 9120 9830 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 10502 9160 10508 9172
rect 10463 9132 10508 9160
rect 9861 9123 9919 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 11422 9160 11428 9172
rect 11383 9132 11428 9160
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 14274 9160 14280 9172
rect 12216 9132 14280 9160
rect 12216 9120 12222 9132
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 15473 9163 15531 9169
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 15930 9160 15936 9172
rect 15519 9132 15936 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 18138 9160 18144 9172
rect 16132 9132 18144 9160
rect 11054 9052 11060 9104
rect 11112 9092 11118 9104
rect 13262 9092 13268 9104
rect 11112 9064 11836 9092
rect 13223 9064 13268 9092
rect 11112 9052 11118 9064
rect 9398 9024 9404 9036
rect 9311 8996 9404 9024
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 9456 8996 11560 9024
rect 9456 8984 9462 8996
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 11532 8965 11560 8996
rect 11808 8968 11836 9064
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 14829 9095 14887 9101
rect 14829 9061 14841 9095
rect 14875 9092 14887 9095
rect 16132 9092 16160 9132
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 19521 9163 19579 9169
rect 19521 9129 19533 9163
rect 19567 9160 19579 9163
rect 20070 9160 20076 9172
rect 19567 9132 20076 9160
rect 19567 9129 19579 9132
rect 19521 9123 19579 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 23385 9163 23443 9169
rect 23385 9160 23397 9163
rect 22428 9132 23397 9160
rect 22428 9120 22434 9132
rect 23385 9129 23397 9132
rect 23431 9129 23443 9163
rect 23385 9123 23443 9129
rect 25222 9120 25228 9172
rect 25280 9160 25286 9172
rect 30745 9163 30803 9169
rect 30745 9160 30757 9163
rect 25280 9132 30757 9160
rect 25280 9120 25286 9132
rect 30745 9129 30757 9132
rect 30791 9129 30803 9163
rect 30745 9123 30803 9129
rect 14875 9064 16160 9092
rect 14875 9061 14887 9064
rect 14829 9055 14887 9061
rect 17310 9052 17316 9104
rect 17368 9092 17374 9104
rect 20165 9095 20223 9101
rect 20165 9092 20177 9095
rect 17368 9064 20177 9092
rect 17368 9052 17374 9064
rect 20165 9061 20177 9064
rect 20211 9061 20223 9095
rect 20165 9055 20223 9061
rect 26050 9052 26056 9104
rect 26108 9092 26114 9104
rect 26108 9064 27200 9092
rect 26108 9052 26114 9064
rect 12710 9024 12716 9036
rect 12671 8996 12716 9024
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 16301 9027 16359 9033
rect 16301 9024 16313 9027
rect 15528 8996 16313 9024
rect 15528 8984 15534 8996
rect 16301 8993 16313 8996
rect 16347 9024 16359 9027
rect 18322 9024 18328 9036
rect 16347 8996 18328 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 18506 9024 18512 9036
rect 18467 8996 18512 9024
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 20438 9024 20444 9036
rect 19444 8996 20444 9024
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 9732 8928 10425 8956
rect 9732 8916 9738 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 11698 8956 11704 8968
rect 11563 8928 11704 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11848 8928 11989 8956
rect 11848 8916 11854 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 14734 8956 14740 8968
rect 13596 8928 14740 8956
rect 13596 8916 13602 8928
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 15381 8959 15439 8965
rect 15381 8958 15393 8959
rect 15304 8956 15393 8958
rect 15068 8930 15393 8956
rect 15068 8928 15332 8930
rect 15068 8916 15074 8928
rect 15381 8925 15393 8930
rect 15427 8925 15439 8959
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 15381 8919 15439 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 19444 8956 19472 8996
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 20809 9027 20867 9033
rect 20809 8993 20821 9027
rect 20855 9024 20867 9027
rect 20898 9024 20904 9036
rect 20855 8996 20904 9024
rect 20855 8993 20867 8996
rect 20809 8987 20867 8993
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 9024 22891 9027
rect 22922 9024 22928 9036
rect 22879 8996 22928 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 22922 8984 22928 8996
rect 22980 9024 22986 9036
rect 24486 9024 24492 9036
rect 22980 8996 24492 9024
rect 22980 8984 22986 8996
rect 24486 8984 24492 8996
rect 24544 9024 24550 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 24544 8996 24593 9024
rect 24544 8984 24550 8996
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24581 8987 24639 8993
rect 24857 9027 24915 9033
rect 24857 8993 24869 9027
rect 24903 9024 24915 9027
rect 25498 9024 25504 9036
rect 24903 8996 25504 9024
rect 24903 8993 24915 8996
rect 24857 8987 24915 8993
rect 25498 8984 25504 8996
rect 25556 8984 25562 9036
rect 26142 8984 26148 9036
rect 26200 9024 26206 9036
rect 26200 8996 26372 9024
rect 26200 8984 26206 8996
rect 17434 8928 19472 8956
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8956 19671 8959
rect 19978 8956 19984 8968
rect 19659 8928 19984 8956
rect 19659 8925 19671 8928
rect 19613 8919 19671 8925
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20254 8956 20260 8968
rect 20215 8928 20260 8956
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 23106 8916 23112 8968
rect 23164 8956 23170 8968
rect 23477 8959 23535 8965
rect 23477 8956 23489 8959
rect 23164 8928 23489 8956
rect 23164 8916 23170 8928
rect 23477 8925 23489 8928
rect 23523 8925 23535 8959
rect 26234 8956 26240 8968
rect 25990 8928 26240 8956
rect 23477 8919 23535 8925
rect 26234 8916 26240 8928
rect 26292 8916 26298 8968
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 12710 8888 12716 8900
rect 10008 8860 12716 8888
rect 10008 8848 10014 8860
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 12805 8891 12863 8897
rect 12805 8857 12817 8891
rect 12851 8857 12863 8891
rect 12805 8851 12863 8857
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12820 8820 12848 8851
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 18046 8888 18052 8900
rect 14976 8860 16712 8888
rect 18007 8860 18052 8888
rect 14976 8848 14982 8860
rect 12115 8792 12848 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 15654 8820 15660 8832
rect 13412 8792 15660 8820
rect 13412 8780 13418 8792
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16574 8820 16580 8832
rect 16080 8792 16580 8820
rect 16080 8780 16086 8792
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 16684 8820 16712 8860
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 18138 8848 18144 8900
rect 18196 8888 18202 8900
rect 20438 8888 20444 8900
rect 18196 8860 20444 8888
rect 18196 8848 18202 8860
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 22094 8848 22100 8900
rect 22152 8848 22158 8900
rect 22557 8891 22615 8897
rect 22557 8857 22569 8891
rect 22603 8857 22615 8891
rect 24026 8888 24032 8900
rect 23987 8860 24032 8888
rect 22557 8851 22615 8857
rect 22370 8820 22376 8832
rect 16684 8792 22376 8820
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 22572 8820 22600 8851
rect 24026 8848 24032 8860
rect 24084 8848 24090 8900
rect 26344 8888 26372 8996
rect 26602 8984 26608 9036
rect 26660 9024 26666 9036
rect 27065 9027 27123 9033
rect 27065 9024 27077 9027
rect 26660 8996 27077 9024
rect 26660 8984 26666 8996
rect 27065 8993 27077 8996
rect 27111 8993 27123 9027
rect 27172 9024 27200 9064
rect 29546 9052 29552 9104
rect 29604 9092 29610 9104
rect 29604 9064 29960 9092
rect 29604 9052 29610 9064
rect 27798 9024 27804 9036
rect 27172 8996 27804 9024
rect 27065 8987 27123 8993
rect 27798 8984 27804 8996
rect 27856 8984 27862 9036
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 29932 9033 29960 9064
rect 29917 9027 29975 9033
rect 29236 8996 29776 9024
rect 29236 8984 29242 8996
rect 29748 8965 29776 8996
rect 29917 8993 29929 9027
rect 29963 8993 29975 9027
rect 29917 8987 29975 8993
rect 30190 8984 30196 9036
rect 30248 9024 30254 9036
rect 31481 9027 31539 9033
rect 31481 9024 31493 9027
rect 30248 8996 31493 9024
rect 30248 8984 30254 8996
rect 31481 8993 31493 8996
rect 31527 8993 31539 9027
rect 31481 8987 31539 8993
rect 29733 8959 29791 8965
rect 29733 8925 29745 8959
rect 29779 8956 29791 8959
rect 29822 8956 29828 8968
rect 29779 8928 29828 8956
rect 29779 8925 29791 8928
rect 29733 8919 29791 8925
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 30282 8916 30288 8968
rect 30340 8956 30346 8968
rect 30653 8959 30711 8965
rect 30653 8956 30665 8959
rect 30340 8928 30665 8956
rect 30340 8916 30346 8928
rect 30653 8925 30665 8928
rect 30699 8925 30711 8959
rect 30653 8919 30711 8925
rect 26602 8888 26608 8900
rect 26344 8860 26608 8888
rect 26602 8848 26608 8860
rect 26660 8848 26666 8900
rect 26970 8848 26976 8900
rect 27028 8888 27034 8900
rect 27341 8891 27399 8897
rect 27341 8888 27353 8891
rect 27028 8860 27353 8888
rect 27028 8848 27034 8860
rect 27341 8857 27353 8860
rect 27387 8857 27399 8891
rect 29178 8888 29184 8900
rect 28566 8860 29184 8888
rect 27341 8851 27399 8857
rect 29178 8848 29184 8860
rect 29236 8848 29242 8900
rect 31573 8891 31631 8897
rect 31573 8857 31585 8891
rect 31619 8888 31631 8891
rect 31754 8888 31760 8900
rect 31619 8860 31760 8888
rect 31619 8857 31631 8860
rect 31573 8851 31631 8857
rect 31754 8848 31760 8860
rect 31812 8848 31818 8900
rect 32125 8891 32183 8897
rect 32125 8857 32137 8891
rect 32171 8857 32183 8891
rect 32125 8851 32183 8857
rect 28813 8823 28871 8829
rect 28813 8820 28825 8823
rect 22572 8792 28825 8820
rect 28813 8789 28825 8792
rect 28859 8820 28871 8823
rect 29270 8820 29276 8832
rect 28859 8792 29276 8820
rect 28859 8789 28871 8792
rect 28813 8783 28871 8789
rect 29270 8780 29276 8792
rect 29328 8780 29334 8832
rect 29638 8780 29644 8832
rect 29696 8820 29702 8832
rect 29914 8820 29920 8832
rect 29696 8792 29920 8820
rect 29696 8780 29702 8792
rect 29914 8780 29920 8792
rect 29972 8820 29978 8832
rect 32140 8820 32168 8851
rect 29972 8792 32168 8820
rect 29972 8780 29978 8792
rect 1104 8730 36892 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 36892 8730
rect 1104 8656 36892 8678
rect 11974 8616 11980 8628
rect 11935 8588 11980 8616
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 13354 8616 13360 8628
rect 13315 8588 13360 8616
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 13909 8619 13967 8625
rect 13909 8616 13921 8619
rect 13872 8588 13921 8616
rect 13872 8576 13878 8588
rect 13909 8585 13921 8588
rect 13955 8585 13967 8619
rect 13909 8579 13967 8585
rect 14553 8619 14611 8625
rect 14553 8585 14565 8619
rect 14599 8616 14611 8619
rect 15378 8616 15384 8628
rect 14599 8588 15384 8616
rect 14599 8585 14611 8588
rect 14553 8579 14611 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15930 8576 15936 8628
rect 15988 8576 15994 8628
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 20622 8616 20628 8628
rect 17828 8588 20628 8616
rect 17828 8576 17834 8588
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21542 8616 21548 8628
rect 21315 8588 21548 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 21542 8576 21548 8588
rect 21600 8616 21606 8628
rect 21818 8616 21824 8628
rect 21600 8588 21824 8616
rect 21600 8576 21606 8588
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22664 8588 24532 8616
rect 10134 8548 10140 8560
rect 10095 8520 10140 8548
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 10686 8548 10692 8560
rect 10647 8520 10692 8548
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 10778 8508 10784 8560
rect 10836 8548 10842 8560
rect 12805 8551 12863 8557
rect 10836 8520 10881 8548
rect 10836 8508 10842 8520
rect 12805 8517 12817 8551
rect 12851 8548 12863 8551
rect 13538 8548 13544 8560
rect 12851 8520 13544 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 15948 8548 15976 8576
rect 15594 8520 15976 8548
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16850 8548 16856 8560
rect 16080 8520 16125 8548
rect 16811 8520 16856 8548
rect 16080 8508 16086 8520
rect 16850 8508 16856 8520
rect 16908 8548 16914 8560
rect 17586 8548 17592 8560
rect 16908 8520 17592 8548
rect 16908 8508 16914 8520
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1673 8483 1731 8489
rect 1673 8480 1685 8483
rect 1636 8452 1685 8480
rect 1636 8440 1642 8452
rect 1673 8449 1685 8452
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 13814 8480 13820 8492
rect 12115 8452 13820 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 13998 8480 14004 8492
rect 13959 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 17420 8489 17448 8520
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 18012 8520 18630 8548
rect 18012 8508 18018 8520
rect 21174 8508 21180 8560
rect 21232 8548 21238 8560
rect 22664 8548 22692 8588
rect 21232 8520 22692 8548
rect 21232 8508 21238 8520
rect 22738 8508 22744 8560
rect 22796 8548 22802 8560
rect 23201 8551 23259 8557
rect 23201 8548 23213 8551
rect 22796 8520 23213 8548
rect 22796 8508 22802 8520
rect 23201 8517 23213 8520
rect 23247 8517 23259 8551
rect 23201 8511 23259 8517
rect 24210 8508 24216 8560
rect 24268 8508 24274 8560
rect 24504 8548 24532 8588
rect 24670 8576 24676 8628
rect 24728 8616 24734 8628
rect 26602 8616 26608 8628
rect 24728 8588 26608 8616
rect 24728 8576 24734 8588
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 28261 8619 28319 8625
rect 28261 8616 28273 8619
rect 27764 8588 28273 8616
rect 27764 8576 27770 8588
rect 28261 8585 28273 8588
rect 28307 8585 28319 8619
rect 28261 8579 28319 8585
rect 24949 8551 25007 8557
rect 24949 8548 24961 8551
rect 24504 8520 24961 8548
rect 24949 8517 24961 8520
rect 24995 8517 25007 8551
rect 24949 8511 25007 8517
rect 26510 8508 26516 8560
rect 26568 8548 26574 8560
rect 30006 8548 30012 8560
rect 26568 8520 30012 8548
rect 26568 8508 26574 8520
rect 30006 8508 30012 8520
rect 30064 8508 30070 8560
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 20254 8440 20260 8492
rect 20312 8480 20318 8492
rect 20717 8483 20775 8489
rect 20717 8480 20729 8483
rect 20312 8452 20729 8480
rect 20312 8440 20318 8452
rect 20717 8449 20729 8452
rect 20763 8480 20775 8483
rect 21818 8480 21824 8492
rect 20763 8452 21824 8480
rect 20763 8449 20775 8452
rect 20717 8443 20775 8449
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 22922 8480 22928 8492
rect 22883 8452 22928 8480
rect 22922 8440 22928 8452
rect 22980 8440 22986 8492
rect 27338 8440 27344 8492
rect 27396 8480 27402 8492
rect 27433 8483 27491 8489
rect 27433 8480 27445 8483
rect 27396 8452 27445 8480
rect 27396 8440 27402 8452
rect 27433 8449 27445 8452
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 12710 8372 12716 8424
rect 12768 8412 12774 8424
rect 16301 8415 16359 8421
rect 12768 8384 16252 8412
rect 12768 8372 12774 8384
rect 1854 8344 1860 8356
rect 1815 8316 1860 8344
rect 1854 8304 1860 8316
rect 1912 8304 1918 8356
rect 9674 8344 9680 8356
rect 9635 8316 9680 8344
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 11606 8304 11612 8356
rect 11664 8344 11670 8356
rect 16224 8344 16252 8384
rect 16301 8381 16313 8415
rect 16347 8412 16359 8415
rect 16574 8412 16580 8424
rect 16347 8384 16580 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 17954 8412 17960 8424
rect 17543 8384 17960 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18138 8412 18144 8424
rect 18095 8384 18144 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18064 8344 18092 8375
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 19484 8384 19809 8412
rect 19484 8372 19490 8384
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 19797 8375 19855 8381
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20530 8412 20536 8424
rect 20119 8384 20536 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 22370 8372 22376 8424
rect 22428 8412 22434 8424
rect 22428 8384 23060 8412
rect 22428 8372 22434 8384
rect 11664 8316 15056 8344
rect 16224 8316 18092 8344
rect 11664 8304 11670 8316
rect 15028 8276 15056 8316
rect 20254 8304 20260 8356
rect 20312 8344 20318 8356
rect 20625 8347 20683 8353
rect 20625 8344 20637 8347
rect 20312 8316 20637 8344
rect 20312 8304 20318 8316
rect 20625 8313 20637 8316
rect 20671 8313 20683 8347
rect 21266 8344 21272 8356
rect 20625 8307 20683 8313
rect 21100 8316 21272 8344
rect 15470 8276 15476 8288
rect 15028 8248 15476 8276
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 21100 8276 21128 8316
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 22278 8344 22284 8356
rect 22239 8316 22284 8344
rect 22278 8304 22284 8316
rect 22336 8344 22342 8356
rect 22830 8344 22836 8356
rect 22336 8316 22836 8344
rect 22336 8304 22342 8316
rect 22830 8304 22836 8316
rect 22888 8304 22894 8356
rect 16080 8248 21128 8276
rect 23032 8276 23060 8384
rect 23658 8372 23664 8424
rect 23716 8412 23722 8424
rect 26234 8412 26240 8424
rect 23716 8384 24440 8412
rect 26195 8384 26240 8412
rect 23716 8372 23722 8384
rect 24412 8356 24440 8384
rect 26234 8372 26240 8384
rect 26292 8412 26298 8424
rect 26418 8412 26424 8424
rect 26292 8384 26424 8412
rect 26292 8372 26298 8384
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 27448 8412 27476 8443
rect 27706 8440 27712 8492
rect 27764 8480 27770 8492
rect 28350 8480 28356 8492
rect 27764 8452 28356 8480
rect 27764 8440 27770 8452
rect 28350 8440 28356 8452
rect 28408 8480 28414 8492
rect 28718 8480 28724 8492
rect 28408 8452 28724 8480
rect 28408 8440 28414 8452
rect 28718 8440 28724 8452
rect 28776 8440 28782 8492
rect 29822 8480 29828 8492
rect 29783 8452 29828 8480
rect 29822 8440 29828 8452
rect 29880 8480 29886 8492
rect 30285 8483 30343 8489
rect 30285 8480 30297 8483
rect 29880 8452 30297 8480
rect 29880 8440 29886 8452
rect 30285 8449 30297 8452
rect 30331 8449 30343 8483
rect 31205 8483 31263 8489
rect 31205 8480 31217 8483
rect 30285 8443 30343 8449
rect 30484 8452 31217 8480
rect 28810 8412 28816 8424
rect 27448 8384 28816 8412
rect 28810 8372 28816 8384
rect 28868 8412 28874 8424
rect 30484 8421 30512 8452
rect 31205 8449 31217 8452
rect 31251 8449 31263 8483
rect 36078 8480 36084 8492
rect 36039 8452 36084 8480
rect 31205 8443 31263 8449
rect 36078 8440 36084 8452
rect 36136 8440 36142 8492
rect 29549 8415 29607 8421
rect 29549 8412 29561 8415
rect 28868 8384 29561 8412
rect 28868 8372 28874 8384
rect 29549 8381 29561 8384
rect 29595 8381 29607 8415
rect 29549 8375 29607 8381
rect 30469 8415 30527 8421
rect 30469 8381 30481 8415
rect 30515 8381 30527 8415
rect 30469 8375 30527 8381
rect 24394 8304 24400 8356
rect 24452 8344 24458 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 24452 8316 25421 8344
rect 24452 8304 24458 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 25409 8307 25467 8313
rect 25682 8304 25688 8356
rect 25740 8344 25746 8356
rect 27341 8347 27399 8353
rect 27341 8344 27353 8347
rect 25740 8316 27353 8344
rect 25740 8304 25746 8316
rect 27341 8313 27353 8316
rect 27387 8313 27399 8347
rect 27341 8307 27399 8313
rect 27448 8316 28396 8344
rect 24670 8276 24676 8288
rect 23032 8248 24676 8276
rect 16080 8236 16086 8248
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 24854 8236 24860 8288
rect 24912 8276 24918 8288
rect 26694 8276 26700 8288
rect 24912 8248 26700 8276
rect 24912 8236 24918 8248
rect 26694 8236 26700 8248
rect 26752 8276 26758 8288
rect 27448 8276 27476 8316
rect 26752 8248 27476 8276
rect 28368 8276 28396 8316
rect 28442 8304 28448 8356
rect 28500 8344 28506 8356
rect 30484 8344 30512 8375
rect 36262 8344 36268 8356
rect 28500 8316 30512 8344
rect 36223 8316 36268 8344
rect 28500 8304 28506 8316
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 28813 8279 28871 8285
rect 28813 8276 28825 8279
rect 28368 8248 28825 8276
rect 26752 8236 26758 8248
rect 28813 8245 28825 8248
rect 28859 8245 28871 8279
rect 31294 8276 31300 8288
rect 31255 8248 31300 8276
rect 28813 8239 28871 8245
rect 31294 8236 31300 8248
rect 31352 8236 31358 8288
rect 1104 8186 36892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36892 8186
rect 1104 8112 36892 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 10686 8032 10692 8084
rect 10744 8072 10750 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10744 8044 10977 8072
rect 10744 8032 10750 8044
rect 10965 8041 10977 8044
rect 11011 8041 11023 8075
rect 10965 8035 11023 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13538 8072 13544 8084
rect 12676 8044 13544 8072
rect 12676 8032 12682 8044
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 18509 8075 18567 8081
rect 14016 8044 16436 8072
rect 10778 7964 10784 8016
rect 10836 8004 10842 8016
rect 10836 7976 12434 8004
rect 10836 7964 10842 7976
rect 10502 7896 10508 7948
rect 10560 7936 10566 7948
rect 10560 7908 12112 7936
rect 10560 7896 10566 7908
rect 6362 7868 6368 7880
rect 6323 7840 6368 7868
rect 6362 7828 6368 7840
rect 6420 7868 6426 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6420 7840 7021 7868
rect 6420 7828 6426 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11882 7868 11888 7880
rect 11103 7840 11888 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 10413 7803 10471 7809
rect 10413 7769 10425 7803
rect 10459 7800 10471 7803
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 10459 7772 11989 7800
rect 10459 7769 10471 7772
rect 10413 7763 10471 7769
rect 11072 7744 11100 7772
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 12084 7800 12112 7908
rect 12406 7868 12434 7976
rect 14016 7868 14044 8044
rect 16408 8004 16436 8044
rect 18509 8041 18521 8075
rect 18555 8072 18567 8075
rect 21174 8072 21180 8084
rect 18555 8044 21180 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 23382 8032 23388 8084
rect 23440 8072 23446 8084
rect 31294 8072 31300 8084
rect 23440 8044 31300 8072
rect 23440 8032 23446 8044
rect 31294 8032 31300 8044
rect 31352 8032 31358 8084
rect 19058 8004 19064 8016
rect 16408 7976 19064 8004
rect 19058 7964 19064 7976
rect 19116 7964 19122 8016
rect 19426 7964 19432 8016
rect 19484 8004 19490 8016
rect 19705 8007 19763 8013
rect 19705 8004 19717 8007
rect 19484 7976 19717 8004
rect 19484 7964 19490 7976
rect 19705 7973 19717 7976
rect 19751 7973 19763 8007
rect 24302 8004 24308 8016
rect 19705 7967 19763 7973
rect 23216 7976 24308 8004
rect 16574 7936 16580 7948
rect 15120 7908 16580 7936
rect 12406 7840 14044 7868
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 15120 7877 15148 7908
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 17129 7939 17187 7945
rect 17129 7905 17141 7939
rect 17175 7936 17187 7939
rect 17218 7936 17224 7948
rect 17175 7908 17224 7936
rect 17175 7905 17187 7908
rect 17129 7899 17187 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 20622 7896 20628 7948
rect 20680 7936 20686 7948
rect 21453 7939 21511 7945
rect 21453 7936 21465 7939
rect 20680 7908 21465 7936
rect 20680 7896 20686 7908
rect 21453 7905 21465 7908
rect 21499 7936 21511 7939
rect 21913 7939 21971 7945
rect 21913 7936 21925 7939
rect 21499 7908 21925 7936
rect 21499 7905 21511 7908
rect 21453 7899 21511 7905
rect 21913 7905 21925 7908
rect 21959 7905 21971 7939
rect 22186 7936 22192 7948
rect 22099 7908 22192 7936
rect 21913 7899 21971 7905
rect 22186 7896 22192 7908
rect 22244 7936 22250 7948
rect 23216 7936 23244 7976
rect 24302 7964 24308 7976
rect 24360 7964 24366 8016
rect 28074 7964 28080 8016
rect 28132 8004 28138 8016
rect 28353 8007 28411 8013
rect 28353 8004 28365 8007
rect 28132 7976 28365 8004
rect 28132 7964 28138 7976
rect 28353 7973 28365 7976
rect 28399 7973 28411 8007
rect 28353 7967 28411 7973
rect 22244 7908 23244 7936
rect 22244 7896 22250 7908
rect 23658 7896 23664 7948
rect 23716 7936 23722 7948
rect 24486 7936 24492 7948
rect 23716 7908 24492 7936
rect 23716 7896 23722 7908
rect 24486 7896 24492 7908
rect 24544 7936 24550 7948
rect 24581 7939 24639 7945
rect 24581 7936 24593 7939
rect 24544 7908 24593 7936
rect 24544 7896 24550 7908
rect 24581 7905 24593 7908
rect 24627 7905 24639 7939
rect 24854 7936 24860 7948
rect 24815 7908 24860 7936
rect 24581 7899 24639 7905
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 25866 7896 25872 7948
rect 25924 7936 25930 7948
rect 27433 7939 27491 7945
rect 27433 7936 27445 7939
rect 25924 7908 27445 7936
rect 25924 7896 25930 7908
rect 27433 7905 27445 7908
rect 27479 7905 27491 7939
rect 28994 7936 29000 7948
rect 27433 7899 27491 7905
rect 27540 7908 29000 7936
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14148 7840 14473 7868
rect 14148 7828 14154 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 13722 7800 13728 7812
rect 12084 7772 12434 7800
rect 13683 7772 13728 7800
rect 11977 7763 12035 7769
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 11054 7692 11060 7744
rect 11112 7692 11118 7744
rect 12406 7732 12434 7772
rect 13722 7760 13728 7772
rect 13780 7800 13786 7812
rect 15120 7800 15148 7831
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17644 7840 17785 7868
rect 17644 7828 17650 7840
rect 17773 7837 17785 7840
rect 17819 7868 17831 7871
rect 18417 7871 18475 7877
rect 18417 7868 18429 7871
rect 17819 7840 18429 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 18417 7837 18429 7840
rect 18463 7868 18475 7871
rect 18506 7868 18512 7880
rect 18463 7840 18512 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 18506 7828 18512 7840
rect 18564 7868 18570 7880
rect 19242 7868 19248 7880
rect 18564 7840 19248 7868
rect 18564 7828 18570 7840
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 26142 7828 26148 7880
rect 26200 7868 26206 7880
rect 27540 7877 27568 7908
rect 28994 7896 29000 7908
rect 29052 7936 29058 7948
rect 30009 7939 30067 7945
rect 30009 7936 30021 7939
rect 29052 7908 30021 7936
rect 29052 7896 29058 7908
rect 30009 7905 30021 7908
rect 30055 7936 30067 7939
rect 30282 7936 30288 7948
rect 30055 7908 30288 7936
rect 30055 7905 30067 7908
rect 30009 7899 30067 7905
rect 30282 7896 30288 7908
rect 30340 7896 30346 7948
rect 27525 7871 27583 7877
rect 26200 7840 27292 7868
rect 26200 7828 26206 7840
rect 13780 7772 15148 7800
rect 15381 7803 15439 7809
rect 13780 7760 13786 7772
rect 15381 7769 15393 7803
rect 15427 7769 15439 7803
rect 17678 7800 17684 7812
rect 16606 7772 17684 7800
rect 15381 7763 15439 7769
rect 14277 7735 14335 7741
rect 14277 7732 14289 7735
rect 12406 7704 14289 7732
rect 14277 7701 14289 7704
rect 14323 7701 14335 7735
rect 15396 7732 15424 7763
rect 17678 7760 17684 7772
rect 17736 7760 17742 7812
rect 17865 7803 17923 7809
rect 17865 7769 17877 7803
rect 17911 7800 17923 7803
rect 17911 7772 20010 7800
rect 17911 7769 17923 7772
rect 17865 7763 17923 7769
rect 20898 7760 20904 7812
rect 20956 7800 20962 7812
rect 21177 7803 21235 7809
rect 21177 7800 21189 7803
rect 20956 7772 21189 7800
rect 20956 7760 20962 7772
rect 21177 7769 21189 7772
rect 21223 7800 21235 7803
rect 21818 7800 21824 7812
rect 21223 7772 21824 7800
rect 21223 7769 21235 7772
rect 21177 7763 21235 7769
rect 21818 7760 21824 7772
rect 21876 7760 21882 7812
rect 23750 7800 23756 7812
rect 23414 7772 23756 7800
rect 23750 7760 23756 7772
rect 23808 7760 23814 7812
rect 27154 7800 27160 7812
rect 26082 7772 27160 7800
rect 27154 7760 27160 7772
rect 27212 7760 27218 7812
rect 27264 7800 27292 7840
rect 27525 7837 27537 7871
rect 27571 7837 27583 7871
rect 27525 7831 27583 7837
rect 28350 7828 28356 7880
rect 28408 7868 28414 7880
rect 28445 7871 28503 7877
rect 28445 7868 28457 7871
rect 28408 7840 28457 7868
rect 28408 7828 28414 7840
rect 28445 7837 28457 7840
rect 28491 7837 28503 7871
rect 28445 7831 28503 7837
rect 28534 7828 28540 7880
rect 28592 7868 28598 7880
rect 29089 7871 29147 7877
rect 29089 7868 29101 7871
rect 28592 7840 29101 7868
rect 28592 7828 28598 7840
rect 29089 7837 29101 7840
rect 29135 7837 29147 7871
rect 29822 7868 29828 7880
rect 29783 7840 29828 7868
rect 29089 7831 29147 7837
rect 29822 7828 29828 7840
rect 29880 7868 29886 7880
rect 32490 7868 32496 7880
rect 29880 7840 32496 7868
rect 29880 7828 29886 7840
rect 32490 7828 32496 7840
rect 32548 7828 32554 7880
rect 29362 7800 29368 7812
rect 27264 7772 29368 7800
rect 29362 7760 29368 7772
rect 29420 7760 29426 7812
rect 16114 7732 16120 7744
rect 15396 7704 16120 7732
rect 14277 7695 14335 7701
rect 16114 7692 16120 7704
rect 16172 7692 16178 7744
rect 20162 7692 20168 7744
rect 20220 7732 20226 7744
rect 22186 7732 22192 7744
rect 20220 7704 22192 7732
rect 20220 7692 20226 7704
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 23661 7735 23719 7741
rect 23661 7701 23673 7735
rect 23707 7732 23719 7735
rect 24946 7732 24952 7744
rect 23707 7704 24952 7732
rect 23707 7701 23719 7704
rect 23661 7695 23719 7701
rect 24946 7692 24952 7704
rect 25004 7732 25010 7744
rect 26142 7732 26148 7744
rect 25004 7704 26148 7732
rect 25004 7692 25010 7704
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 26329 7735 26387 7741
rect 26329 7701 26341 7735
rect 26375 7732 26387 7735
rect 26510 7732 26516 7744
rect 26375 7704 26516 7732
rect 26375 7701 26387 7704
rect 26329 7695 26387 7701
rect 26510 7692 26516 7704
rect 26568 7692 26574 7744
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 28997 7735 29055 7741
rect 28997 7732 29009 7735
rect 26752 7704 29009 7732
rect 26752 7692 26758 7704
rect 28997 7701 29009 7704
rect 29043 7701 29055 7735
rect 28997 7695 29055 7701
rect 1104 7642 36892 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 36892 7642
rect 1104 7568 36892 7590
rect 12066 7488 12072 7540
rect 12124 7488 12130 7540
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 13630 7528 13636 7540
rect 12584 7500 13636 7528
rect 12584 7488 12590 7500
rect 13630 7488 13636 7500
rect 13688 7528 13694 7540
rect 13725 7531 13783 7537
rect 13725 7528 13737 7531
rect 13688 7500 13737 7528
rect 13688 7488 13694 7500
rect 13725 7497 13737 7500
rect 13771 7497 13783 7531
rect 20162 7528 20168 7540
rect 13725 7491 13783 7497
rect 13832 7500 15884 7528
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2130 7460 2136 7472
rect 1903 7432 2136 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 10134 7420 10140 7472
rect 10192 7460 10198 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 10192 7432 10425 7460
rect 10192 7420 10198 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10962 7460 10968 7472
rect 10923 7432 10968 7460
rect 10413 7423 10471 7429
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 11330 7460 11336 7472
rect 11103 7432 11336 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11330 7420 11336 7432
rect 11388 7420 11394 7472
rect 12084 7460 12112 7488
rect 12253 7463 12311 7469
rect 12253 7460 12265 7463
rect 12084 7432 12265 7460
rect 12253 7429 12265 7432
rect 12299 7429 12311 7463
rect 12253 7423 12311 7429
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 13832 7460 13860 7500
rect 13596 7432 13860 7460
rect 13596 7420 13602 7432
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 11974 7324 11980 7336
rect 11935 7296 11980 7324
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 13372 7256 13400 7378
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13780 7364 14289 7392
rect 13780 7352 13786 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 15856 7392 15884 7500
rect 16316 7500 20168 7528
rect 16316 7469 16344 7500
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 23382 7528 23388 7540
rect 20272 7500 23388 7528
rect 16301 7463 16359 7469
rect 16301 7429 16313 7463
rect 16347 7429 16359 7463
rect 16301 7423 16359 7429
rect 17218 7420 17224 7472
rect 17276 7460 17282 7472
rect 17313 7463 17371 7469
rect 17313 7460 17325 7463
rect 17276 7432 17325 7460
rect 17276 7420 17282 7432
rect 17313 7429 17325 7432
rect 17359 7429 17371 7463
rect 17313 7423 17371 7429
rect 17862 7420 17868 7472
rect 17920 7460 17926 7472
rect 17957 7463 18015 7469
rect 17957 7460 17969 7463
rect 17920 7432 17969 7460
rect 17920 7420 17926 7432
rect 17957 7429 17969 7432
rect 18003 7429 18015 7463
rect 20272 7460 20300 7500
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 29178 7528 29184 7540
rect 23492 7500 25728 7528
rect 29139 7500 29184 7528
rect 19918 7432 20300 7460
rect 20349 7463 20407 7469
rect 17957 7423 18015 7429
rect 20349 7429 20361 7463
rect 20395 7460 20407 7463
rect 20395 7432 21220 7460
rect 20395 7429 20407 7432
rect 20349 7423 20407 7429
rect 19058 7392 19064 7404
rect 14277 7355 14335 7361
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14550 7324 14556 7336
rect 14240 7296 14556 7324
rect 14240 7284 14246 7296
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 15672 7324 15700 7378
rect 15856 7364 19064 7392
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 15672 7296 20576 7324
rect 20548 7256 20576 7296
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 21192 7324 21220 7432
rect 21818 7420 21824 7472
rect 21876 7460 21882 7472
rect 22005 7463 22063 7469
rect 22005 7460 22017 7463
rect 21876 7432 22017 7460
rect 21876 7420 21882 7432
rect 22005 7429 22017 7432
rect 22051 7429 22063 7463
rect 22005 7423 22063 7429
rect 22649 7463 22707 7469
rect 22649 7429 22661 7463
rect 22695 7460 22707 7463
rect 22738 7460 22744 7472
rect 22695 7432 22744 7460
rect 22695 7429 22707 7432
rect 22649 7423 22707 7429
rect 22738 7420 22744 7432
rect 22796 7420 22802 7472
rect 21266 7352 21272 7404
rect 21324 7392 21330 7404
rect 23492 7392 23520 7500
rect 24210 7460 24216 7472
rect 21324 7364 23520 7392
rect 23584 7432 24216 7460
rect 21324 7352 21330 7364
rect 22738 7324 22744 7336
rect 20680 7296 20725 7324
rect 21192 7296 22744 7324
rect 20680 7284 20686 7296
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 23201 7327 23259 7333
rect 23201 7293 23213 7327
rect 23247 7324 23259 7327
rect 23584 7324 23612 7432
rect 24210 7420 24216 7432
rect 24268 7420 24274 7472
rect 25590 7460 25596 7472
rect 25162 7432 25596 7460
rect 25590 7420 25596 7432
rect 25648 7420 25654 7472
rect 25700 7469 25728 7500
rect 29178 7488 29184 7500
rect 29236 7488 29242 7540
rect 25685 7463 25743 7469
rect 25685 7429 25697 7463
rect 25731 7429 25743 7463
rect 26694 7460 26700 7472
rect 25685 7423 25743 7429
rect 25792 7432 26700 7460
rect 25498 7352 25504 7404
rect 25556 7392 25562 7404
rect 25792 7392 25820 7432
rect 26694 7420 26700 7432
rect 26752 7420 26758 7472
rect 35894 7420 35900 7472
rect 35952 7460 35958 7472
rect 36081 7463 36139 7469
rect 36081 7460 36093 7463
rect 35952 7432 36093 7460
rect 35952 7420 35958 7432
rect 36081 7429 36093 7432
rect 36127 7429 36139 7463
rect 36081 7423 36139 7429
rect 25556 7364 25820 7392
rect 26605 7395 26663 7401
rect 25556 7352 25562 7364
rect 26605 7361 26617 7395
rect 26651 7392 26663 7395
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 26651 7364 27353 7392
rect 26651 7361 26663 7364
rect 26605 7355 26663 7361
rect 27341 7361 27353 7364
rect 27387 7392 27399 7395
rect 27890 7392 27896 7404
rect 27387 7364 27896 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 27890 7352 27896 7364
rect 27948 7352 27954 7404
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7392 28043 7395
rect 28074 7392 28080 7404
rect 28031 7364 28080 7392
rect 28031 7361 28043 7364
rect 27985 7355 28043 7361
rect 28074 7352 28080 7364
rect 28132 7392 28138 7404
rect 28534 7392 28540 7404
rect 28132 7364 28540 7392
rect 28132 7352 28138 7364
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 28629 7395 28687 7401
rect 28629 7361 28641 7395
rect 28675 7392 28687 7395
rect 28994 7392 29000 7404
rect 28675 7364 29000 7392
rect 28675 7361 28687 7364
rect 28629 7355 28687 7361
rect 28994 7352 29000 7364
rect 29052 7352 29058 7404
rect 29273 7395 29331 7401
rect 29273 7361 29285 7395
rect 29319 7361 29331 7395
rect 29273 7355 29331 7361
rect 23247 7296 23612 7324
rect 23247 7293 23259 7296
rect 23201 7287 23259 7293
rect 23658 7284 23664 7336
rect 23716 7324 23722 7336
rect 23934 7324 23940 7336
rect 23716 7296 23761 7324
rect 23895 7296 23940 7324
rect 23716 7284 23722 7296
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 24026 7284 24032 7336
rect 24084 7324 24090 7336
rect 26513 7327 26571 7333
rect 26513 7324 26525 7327
rect 24084 7296 26525 7324
rect 24084 7284 24090 7296
rect 26513 7293 26525 7296
rect 26559 7293 26571 7327
rect 28552 7324 28580 7352
rect 29288 7324 29316 7355
rect 29546 7352 29552 7404
rect 29604 7392 29610 7404
rect 29917 7395 29975 7401
rect 29917 7392 29929 7395
rect 29604 7364 29929 7392
rect 29604 7352 29610 7364
rect 29917 7361 29929 7364
rect 29963 7392 29975 7395
rect 30377 7395 30435 7401
rect 30377 7392 30389 7395
rect 29963 7364 30389 7392
rect 29963 7361 29975 7364
rect 29917 7355 29975 7361
rect 30377 7361 30389 7364
rect 30423 7361 30435 7395
rect 30377 7355 30435 7361
rect 35621 7395 35679 7401
rect 35621 7361 35633 7395
rect 35667 7392 35679 7395
rect 35802 7392 35808 7404
rect 35667 7364 35808 7392
rect 35667 7361 35679 7364
rect 35621 7355 35679 7361
rect 35802 7352 35808 7364
rect 35860 7392 35866 7404
rect 36265 7395 36323 7401
rect 36265 7392 36277 7395
rect 35860 7364 36277 7392
rect 35860 7352 35866 7364
rect 36265 7361 36277 7364
rect 36311 7361 36323 7395
rect 36265 7355 36323 7361
rect 28552 7296 29316 7324
rect 26513 7287 26571 7293
rect 20990 7256 20996 7268
rect 13372 7228 14412 7256
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 9674 7188 9680 7200
rect 2188 7160 9680 7188
rect 2188 7148 2194 7160
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 14274 7188 14280 7200
rect 12124 7160 14280 7188
rect 12124 7148 12130 7160
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14384 7188 14412 7228
rect 17236 7228 19012 7256
rect 20548 7228 20996 7256
rect 17236 7188 17264 7228
rect 14384 7160 17264 7188
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 18874 7188 18880 7200
rect 18472 7160 18880 7188
rect 18472 7148 18478 7160
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 18984 7188 19012 7228
rect 20990 7216 20996 7228
rect 21048 7216 21054 7268
rect 21100 7228 22094 7256
rect 21100 7188 21128 7228
rect 18984 7160 21128 7188
rect 21269 7191 21327 7197
rect 21269 7157 21281 7191
rect 21315 7188 21327 7191
rect 21450 7188 21456 7200
rect 21315 7160 21456 7188
rect 21315 7157 21327 7160
rect 21269 7151 21327 7157
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 22066 7188 22094 7228
rect 22186 7216 22192 7268
rect 22244 7256 22250 7268
rect 29825 7259 29883 7265
rect 29825 7256 29837 7259
rect 22244 7228 23796 7256
rect 22244 7216 22250 7228
rect 23566 7188 23572 7200
rect 22066 7160 23572 7188
rect 23566 7148 23572 7160
rect 23624 7148 23630 7200
rect 23768 7188 23796 7228
rect 25976 7228 29837 7256
rect 25976 7188 26004 7228
rect 29825 7225 29837 7228
rect 29871 7225 29883 7259
rect 29825 7219 29883 7225
rect 27246 7188 27252 7200
rect 23768 7160 26004 7188
rect 27207 7160 27252 7188
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 27522 7148 27528 7200
rect 27580 7188 27586 7200
rect 27893 7191 27951 7197
rect 27893 7188 27905 7191
rect 27580 7160 27905 7188
rect 27580 7148 27586 7160
rect 27893 7157 27905 7160
rect 27939 7157 27951 7191
rect 28534 7188 28540 7200
rect 28495 7160 28540 7188
rect 27893 7151 27951 7157
rect 28534 7148 28540 7160
rect 28592 7148 28598 7200
rect 30374 7148 30380 7200
rect 30432 7188 30438 7200
rect 30469 7191 30527 7197
rect 30469 7188 30481 7191
rect 30432 7160 30481 7188
rect 30432 7148 30438 7160
rect 30469 7157 30481 7160
rect 30515 7157 30527 7191
rect 30469 7151 30527 7157
rect 1104 7098 36892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36892 7098
rect 1104 7024 36892 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 10505 6987 10563 6993
rect 10505 6953 10517 6987
rect 10551 6984 10563 6987
rect 10962 6984 10968 6996
rect 10551 6956 10968 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12066 6984 12072 6996
rect 11572 6956 12072 6984
rect 11572 6944 11578 6956
rect 12066 6944 12072 6956
rect 12124 6984 12130 6996
rect 12234 6987 12292 6993
rect 12234 6984 12246 6987
rect 12124 6956 12246 6984
rect 12124 6944 12130 6956
rect 12234 6953 12246 6956
rect 12280 6953 12292 6987
rect 12234 6947 12292 6953
rect 14274 6944 14280 6996
rect 14332 6984 14338 6996
rect 14918 6984 14924 6996
rect 14332 6956 14924 6984
rect 14332 6944 14338 6956
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 15194 6993 15200 6996
rect 15184 6987 15200 6993
rect 15184 6953 15196 6987
rect 15184 6947 15200 6953
rect 15194 6944 15200 6947
rect 15252 6944 15258 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 20898 6984 20904 6996
rect 15620 6956 20904 6984
rect 15620 6944 15626 6956
rect 20898 6944 20904 6956
rect 20956 6944 20962 6996
rect 21818 6944 21824 6996
rect 21876 6984 21882 6996
rect 27246 6984 27252 6996
rect 21876 6956 27252 6984
rect 21876 6944 21882 6956
rect 27246 6944 27252 6956
rect 27304 6944 27310 6996
rect 14182 6876 14188 6928
rect 14240 6916 14246 6928
rect 14240 6888 15056 6916
rect 14240 6876 14246 6888
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9766 6848 9772 6860
rect 9355 6820 9772 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6848 10011 6851
rect 10134 6848 10140 6860
rect 9999 6820 10140 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13596 6820 13737 6848
rect 13596 6808 13602 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 14516 6820 14933 6848
rect 14516 6808 14522 6820
rect 14921 6817 14933 6820
rect 14967 6817 14979 6851
rect 15028 6848 15056 6888
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 19426 6916 19432 6928
rect 17920 6888 19432 6916
rect 17920 6876 17926 6888
rect 19426 6876 19432 6888
rect 19484 6876 19490 6928
rect 21910 6876 21916 6928
rect 21968 6916 21974 6928
rect 28534 6916 28540 6928
rect 21968 6888 28540 6916
rect 21968 6876 21974 6888
rect 28534 6876 28540 6888
rect 28592 6876 28598 6928
rect 17494 6848 17500 6860
rect 15028 6820 17500 6848
rect 14921 6811 14979 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 18104 6820 19533 6848
rect 18104 6808 18110 6820
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 20257 6851 20315 6857
rect 20257 6817 20269 6851
rect 20303 6848 20315 6851
rect 22094 6848 22100 6860
rect 20303 6820 22100 6848
rect 20303 6817 20315 6820
rect 20257 6811 20315 6817
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22281 6851 22339 6857
rect 22281 6817 22293 6851
rect 22327 6848 22339 6851
rect 24394 6848 24400 6860
rect 22327 6820 24400 6848
rect 22327 6817 22339 6820
rect 22281 6811 22339 6817
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 24581 6851 24639 6857
rect 24581 6848 24593 6851
rect 24544 6820 24593 6848
rect 24544 6808 24550 6820
rect 24581 6817 24593 6820
rect 24627 6817 24639 6851
rect 24581 6811 24639 6817
rect 24762 6808 24768 6860
rect 24820 6848 24826 6860
rect 29825 6851 29883 6857
rect 29825 6848 29837 6851
rect 24820 6820 29837 6848
rect 24820 6808 24826 6820
rect 29825 6817 29837 6820
rect 29871 6817 29883 6851
rect 29825 6811 29883 6817
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6780 10471 6783
rect 19334 6780 19340 6792
rect 10459 6752 11192 6780
rect 13386 6752 14872 6780
rect 16330 6752 19340 6780
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 9398 6672 9404 6724
rect 9456 6712 9462 6724
rect 9456 6684 9501 6712
rect 9456 6672 9462 6684
rect 11164 6653 11192 6752
rect 14844 6712 14872 6752
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 23198 6780 23204 6792
rect 21666 6752 23204 6780
rect 23198 6740 23204 6752
rect 23256 6740 23262 6792
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6780 26387 6783
rect 26375 6752 26464 6780
rect 26375 6749 26387 6752
rect 26329 6743 26387 6749
rect 16942 6712 16948 6724
rect 14844 6684 15608 6712
rect 16903 6684 16948 6712
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 11238 6644 11244 6656
rect 11195 6616 11244 6644
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 13906 6644 13912 6656
rect 12492 6616 13912 6644
rect 12492 6604 12498 6616
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14461 6647 14519 6653
rect 14461 6613 14473 6647
rect 14507 6644 14519 6647
rect 14550 6644 14556 6656
rect 14507 6616 14556 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15580 6644 15608 6684
rect 16942 6672 16948 6684
rect 17000 6672 17006 6724
rect 18230 6712 18236 6724
rect 17052 6684 18236 6712
rect 17052 6644 17080 6684
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 18417 6715 18475 6721
rect 18417 6681 18429 6715
rect 18463 6712 18475 6715
rect 18506 6712 18512 6724
rect 18463 6684 18512 6712
rect 18463 6681 18475 6684
rect 18417 6675 18475 6681
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 19058 6672 19064 6724
rect 19116 6712 19122 6724
rect 20533 6715 20591 6721
rect 20533 6712 20545 6715
rect 19116 6684 20545 6712
rect 19116 6672 19122 6684
rect 20533 6681 20545 6684
rect 20579 6681 20591 6715
rect 20533 6675 20591 6681
rect 21910 6672 21916 6724
rect 21968 6712 21974 6724
rect 23934 6712 23940 6724
rect 21968 6684 23940 6712
rect 21968 6672 21974 6684
rect 23934 6672 23940 6684
rect 23992 6672 23998 6724
rect 15580 6616 17080 6644
rect 17126 6604 17132 6656
rect 17184 6644 17190 6656
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 17184 6616 17509 6644
rect 17184 6604 17190 6616
rect 17497 6613 17509 6616
rect 17543 6644 17555 6647
rect 20806 6644 20812 6656
rect 17543 6616 20812 6644
rect 17543 6613 17555 6616
rect 17497 6607 17555 6613
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 21450 6604 21456 6656
rect 21508 6644 21514 6656
rect 23014 6644 23020 6656
rect 21508 6616 23020 6644
rect 21508 6604 21514 6616
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23198 6644 23204 6656
rect 23159 6616 23204 6644
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 23658 6644 23664 6656
rect 23619 6616 23664 6644
rect 23658 6604 23664 6616
rect 23716 6604 23722 6656
rect 26436 6644 26464 6752
rect 26602 6740 26608 6792
rect 26660 6780 26666 6792
rect 27433 6783 27491 6789
rect 27433 6780 27445 6783
rect 26660 6752 27445 6780
rect 26660 6740 26666 6752
rect 27433 6749 27445 6752
rect 27479 6749 27491 6783
rect 27433 6743 27491 6749
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6780 27583 6783
rect 28074 6780 28080 6792
rect 27571 6752 28080 6780
rect 27571 6749 27583 6752
rect 27525 6743 27583 6749
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 28169 6783 28227 6789
rect 28169 6749 28181 6783
rect 28215 6780 28227 6783
rect 28810 6780 28816 6792
rect 28215 6752 28816 6780
rect 28215 6749 28227 6752
rect 28169 6743 28227 6749
rect 28810 6740 28816 6752
rect 28868 6740 28874 6792
rect 28994 6740 29000 6792
rect 29052 6780 29058 6792
rect 29917 6783 29975 6789
rect 29917 6780 29929 6783
rect 29052 6752 29929 6780
rect 29052 6740 29058 6752
rect 29917 6749 29929 6752
rect 29963 6780 29975 6783
rect 30282 6780 30288 6792
rect 29963 6752 30288 6780
rect 29963 6749 29975 6752
rect 29917 6743 29975 6749
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 32490 6780 32496 6792
rect 32451 6752 32496 6780
rect 32490 6740 32496 6752
rect 32548 6740 32554 6792
rect 26694 6672 26700 6724
rect 26752 6712 26758 6724
rect 26789 6715 26847 6721
rect 26789 6712 26801 6715
rect 26752 6684 26801 6712
rect 26752 6672 26758 6684
rect 26789 6681 26801 6684
rect 26835 6681 26847 6715
rect 26789 6675 26847 6681
rect 31846 6672 31852 6724
rect 31904 6712 31910 6724
rect 32769 6715 32827 6721
rect 32769 6712 32781 6715
rect 31904 6684 32781 6712
rect 31904 6672 31910 6684
rect 32769 6681 32781 6684
rect 32815 6681 32827 6715
rect 32769 6675 32827 6681
rect 27246 6644 27252 6656
rect 26436 6616 27252 6644
rect 27246 6604 27252 6616
rect 27304 6604 27310 6656
rect 28074 6644 28080 6656
rect 28035 6616 28080 6644
rect 28074 6604 28080 6616
rect 28132 6604 28138 6656
rect 28718 6644 28724 6656
rect 28679 6616 28724 6644
rect 28718 6604 28724 6616
rect 28776 6604 28782 6656
rect 1104 6554 36892 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 36892 6554
rect 1104 6480 36892 6502
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8260 6412 8493 6440
rect 8260 6400 8266 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9824 6412 9873 6440
rect 9824 6400 9830 6412
rect 9861 6409 9873 6412
rect 9907 6409 9919 6443
rect 9861 6403 9919 6409
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 14458 6440 14464 6452
rect 12032 6412 14464 6440
rect 12032 6400 12038 6412
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6304 8079 6307
rect 8220 6304 8248 6400
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 11422 6372 11428 6384
rect 10643 6344 11428 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 12360 6313 12388 6412
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 17126 6440 17132 6452
rect 14568 6412 17132 6440
rect 13906 6332 13912 6384
rect 13964 6372 13970 6384
rect 14568 6372 14596 6412
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 20254 6440 20260 6452
rect 17788 6412 20260 6440
rect 17788 6372 17816 6412
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 22094 6440 22100 6452
rect 22066 6400 22100 6440
rect 22152 6400 22158 6452
rect 23658 6440 23664 6452
rect 22296 6412 23664 6440
rect 13964 6344 14596 6372
rect 15594 6344 17816 6372
rect 19153 6375 19211 6381
rect 13964 6332 13970 6344
rect 19153 6341 19165 6375
rect 19199 6372 19211 6375
rect 20622 6372 20628 6384
rect 19199 6344 20628 6372
rect 19199 6341 19211 6344
rect 19153 6335 19211 6341
rect 20622 6332 20628 6344
rect 20680 6332 20686 6384
rect 22066 6372 22094 6400
rect 22296 6384 22324 6412
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 23842 6400 23848 6452
rect 23900 6440 23906 6452
rect 26234 6440 26240 6452
rect 23900 6412 26240 6440
rect 23900 6400 23906 6412
rect 26234 6400 26240 6412
rect 26292 6400 26298 6452
rect 22278 6372 22284 6384
rect 22020 6344 22094 6372
rect 22191 6344 22284 6372
rect 8067 6276 8248 6304
rect 12345 6307 12403 6313
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 12345 6273 12357 6307
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 17402 6304 17408 6316
rect 17363 6276 17408 6304
rect 17402 6264 17408 6276
rect 17460 6304 17466 6316
rect 17460 6276 19334 6304
rect 17460 6264 17466 6276
rect 19306 6248 19334 6276
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 22020 6313 22048 6344
rect 22278 6332 22284 6344
rect 22336 6332 22342 6384
rect 23290 6332 23296 6384
rect 23348 6332 23354 6384
rect 24857 6375 24915 6381
rect 24857 6341 24869 6375
rect 24903 6372 24915 6375
rect 24946 6372 24952 6384
rect 24903 6344 24952 6372
rect 24903 6341 24915 6344
rect 24857 6335 24915 6341
rect 24946 6332 24952 6344
rect 25004 6332 25010 6384
rect 27798 6372 27804 6384
rect 27759 6344 27804 6372
rect 27798 6332 27804 6344
rect 27856 6332 27862 6384
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21324 6276 21373 6304
rect 21324 6264 21330 6276
rect 21361 6273 21373 6276
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6273 22063 6307
rect 27890 6304 27896 6316
rect 22005 6267 22063 6273
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9732 6208 10517 6236
rect 9732 6196 9738 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 13814 6236 13820 6248
rect 12667 6208 13820 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14424 6208 14565 6236
rect 14424 6196 14430 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 14700 6208 16037 6236
rect 14700 6196 14706 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 16850 6236 16856 6248
rect 16347 6208 16856 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 17586 6236 17592 6248
rect 16908 6208 17592 6236
rect 16908 6196 16914 6208
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 19242 6196 19248 6248
rect 19300 6236 19334 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19300 6208 19625 6236
rect 19300 6196 19306 6208
rect 19613 6205 19625 6208
rect 19659 6205 19671 6239
rect 22278 6236 22284 6248
rect 19613 6199 19671 6205
rect 22066 6208 22284 6236
rect 11057 6171 11115 6177
rect 11057 6137 11069 6171
rect 11103 6168 11115 6171
rect 11103 6140 12480 6168
rect 11103 6137 11115 6140
rect 11057 6131 11115 6137
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11698 6100 11704 6112
rect 11572 6072 11704 6100
rect 11572 6060 11578 6072
rect 11698 6060 11704 6072
rect 11756 6100 11762 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11756 6072 11805 6100
rect 11756 6060 11762 6072
rect 11793 6069 11805 6072
rect 11839 6100 11851 6103
rect 12342 6100 12348 6112
rect 11839 6072 12348 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 12452 6100 12480 6140
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 13964 6140 14105 6168
rect 13964 6128 13970 6140
rect 14093 6137 14105 6140
rect 14139 6168 14151 6171
rect 15010 6168 15016 6180
rect 14139 6140 15016 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 18506 6168 18512 6180
rect 16868 6140 18512 6168
rect 13998 6100 14004 6112
rect 12452 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 16868 6109 16896 6140
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 18874 6128 18880 6180
rect 18932 6168 18938 6180
rect 22066 6168 22094 6208
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 23014 6196 23020 6248
rect 23072 6236 23078 6248
rect 24029 6239 24087 6245
rect 24029 6236 24041 6239
rect 23072 6208 24041 6236
rect 23072 6196 23078 6208
rect 24029 6205 24041 6208
rect 24075 6205 24087 6239
rect 24578 6236 24584 6248
rect 24539 6208 24584 6236
rect 24029 6199 24087 6205
rect 24578 6196 24584 6208
rect 24636 6196 24642 6248
rect 25976 6236 26004 6290
rect 27851 6276 27896 6304
rect 27890 6264 27896 6276
rect 27948 6264 27954 6316
rect 29089 6307 29147 6313
rect 29089 6273 29101 6307
rect 29135 6304 29147 6307
rect 29546 6304 29552 6316
rect 29135 6276 29552 6304
rect 29135 6273 29147 6276
rect 29089 6267 29147 6273
rect 29546 6264 29552 6276
rect 29604 6304 29610 6316
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29604 6276 29745 6304
rect 29604 6264 29610 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 30282 6264 30288 6316
rect 30340 6304 30346 6316
rect 30377 6307 30435 6313
rect 30377 6304 30389 6307
rect 30340 6276 30389 6304
rect 30340 6264 30346 6276
rect 30377 6273 30389 6276
rect 30423 6273 30435 6307
rect 30377 6267 30435 6273
rect 27522 6236 27528 6248
rect 25976 6208 27528 6236
rect 27522 6196 27528 6208
rect 27580 6196 27586 6248
rect 30285 6171 30343 6177
rect 30285 6168 30297 6171
rect 18932 6140 22094 6168
rect 25884 6140 30297 6168
rect 18932 6128 18938 6140
rect 16853 6103 16911 6109
rect 16853 6069 16865 6103
rect 16899 6069 16911 6103
rect 16853 6063 16911 6069
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 22922 6100 22928 6112
rect 17000 6072 22928 6100
rect 17000 6060 17006 6072
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 23474 6060 23480 6112
rect 23532 6100 23538 6112
rect 25884 6100 25912 6140
rect 30285 6137 30297 6140
rect 30331 6137 30343 6171
rect 30285 6131 30343 6137
rect 23532 6072 25912 6100
rect 26329 6103 26387 6109
rect 23532 6060 23538 6072
rect 26329 6069 26341 6103
rect 26375 6100 26387 6103
rect 26970 6100 26976 6112
rect 26375 6072 26976 6100
rect 26375 6069 26387 6072
rect 26329 6063 26387 6069
rect 26970 6060 26976 6072
rect 27028 6060 27034 6112
rect 27246 6100 27252 6112
rect 27207 6072 27252 6100
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 28997 6103 29055 6109
rect 28997 6069 29009 6103
rect 29043 6100 29055 6103
rect 29086 6100 29092 6112
rect 29043 6072 29092 6100
rect 29043 6069 29055 6072
rect 28997 6063 29055 6069
rect 29086 6060 29092 6072
rect 29144 6060 29150 6112
rect 29638 6100 29644 6112
rect 29599 6072 29644 6100
rect 29638 6060 29644 6072
rect 29696 6060 29702 6112
rect 1104 6010 36892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36892 6010
rect 1104 5936 36892 5958
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 9398 5896 9404 5908
rect 9263 5868 9404 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 11422 5896 11428 5908
rect 11383 5868 11428 5896
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 13906 5896 13912 5908
rect 12308 5868 13912 5896
rect 12308 5856 12314 5868
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 22186 5896 22192 5908
rect 14056 5868 22192 5896
rect 14056 5856 14062 5868
rect 22186 5856 22192 5868
rect 22244 5856 22250 5908
rect 24581 5899 24639 5905
rect 24581 5865 24593 5899
rect 24627 5896 24639 5899
rect 24854 5896 24860 5908
rect 24627 5868 24860 5896
rect 24627 5865 24639 5868
rect 24581 5859 24639 5865
rect 24854 5856 24860 5868
rect 24912 5896 24918 5908
rect 25958 5896 25964 5908
rect 24912 5868 25964 5896
rect 24912 5856 24918 5868
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 26234 5856 26240 5908
rect 26292 5896 26298 5908
rect 26789 5899 26847 5905
rect 26789 5896 26801 5899
rect 26292 5868 26801 5896
rect 26292 5856 26298 5868
rect 26789 5865 26801 5868
rect 26835 5865 26847 5899
rect 31754 5896 31760 5908
rect 31715 5868 31760 5896
rect 26789 5859 26847 5865
rect 31754 5856 31760 5868
rect 31812 5856 31818 5908
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 9180 5800 12112 5828
rect 9180 5788 9186 5800
rect 11974 5760 11980 5772
rect 11935 5732 11980 5760
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12084 5760 12112 5800
rect 14090 5788 14096 5840
rect 14148 5828 14154 5840
rect 14277 5831 14335 5837
rect 14277 5828 14289 5831
rect 14148 5800 14289 5828
rect 14148 5788 14154 5800
rect 14277 5797 14289 5800
rect 14323 5797 14335 5831
rect 14918 5828 14924 5840
rect 14879 5800 14924 5828
rect 14277 5791 14335 5797
rect 14918 5788 14924 5800
rect 14976 5788 14982 5840
rect 18233 5831 18291 5837
rect 18233 5797 18245 5831
rect 18279 5828 18291 5831
rect 18322 5828 18328 5840
rect 18279 5800 18328 5828
rect 18279 5797 18291 5800
rect 18233 5791 18291 5797
rect 18322 5788 18328 5800
rect 18380 5788 18386 5840
rect 18506 5788 18512 5840
rect 18564 5828 18570 5840
rect 18693 5831 18751 5837
rect 18693 5828 18705 5831
rect 18564 5800 18705 5828
rect 18564 5788 18570 5800
rect 18693 5797 18705 5800
rect 18739 5797 18751 5831
rect 21542 5828 21548 5840
rect 18693 5791 18751 5797
rect 18892 5800 21548 5828
rect 15562 5760 15568 5772
rect 12084 5732 15568 5760
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 17586 5760 17592 5772
rect 17547 5732 17592 5760
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 18892 5760 18920 5800
rect 21542 5788 21548 5800
rect 21600 5788 21606 5840
rect 17920 5732 18920 5760
rect 17920 5720 17926 5732
rect 20346 5720 20352 5772
rect 20404 5760 20410 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20404 5732 21005 5760
rect 20404 5720 20410 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5760 22799 5763
rect 23842 5760 23848 5772
rect 22787 5732 23848 5760
rect 22787 5729 22799 5732
rect 22741 5723 22799 5729
rect 23842 5720 23848 5732
rect 23900 5720 23906 5772
rect 24578 5720 24584 5772
rect 24636 5760 24642 5772
rect 26329 5763 26387 5769
rect 26329 5760 26341 5763
rect 24636 5732 26341 5760
rect 24636 5720 24642 5732
rect 26329 5729 26341 5732
rect 26375 5729 26387 5763
rect 26329 5723 26387 5729
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 11146 5692 11152 5704
rect 9355 5664 11152 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11514 5692 11520 5704
rect 11475 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 15838 5692 15844 5704
rect 13596 5664 15844 5692
rect 13596 5652 13602 5664
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 21450 5692 21456 5704
rect 18156 5664 21456 5692
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 11974 5624 11980 5636
rect 11848 5596 11980 5624
rect 11848 5584 11854 5596
rect 11974 5584 11980 5596
rect 12032 5624 12038 5636
rect 12253 5627 12311 5633
rect 12253 5624 12265 5627
rect 12032 5596 12265 5624
rect 12032 5584 12038 5596
rect 12253 5593 12265 5596
rect 12299 5593 12311 5627
rect 13630 5624 13636 5636
rect 13478 5596 13636 5624
rect 12253 5587 12311 5593
rect 13630 5584 13636 5596
rect 13688 5584 13694 5636
rect 16298 5584 16304 5636
rect 16356 5584 16362 5636
rect 17313 5627 17371 5633
rect 17313 5593 17325 5627
rect 17359 5624 17371 5627
rect 18046 5624 18052 5636
rect 17359 5596 18052 5624
rect 17359 5593 17371 5596
rect 17313 5587 17371 5593
rect 18046 5584 18052 5596
rect 18104 5584 18110 5636
rect 13722 5556 13728 5568
rect 13683 5528 13728 5556
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 18156 5556 18184 5664
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 23017 5695 23075 5701
rect 23017 5661 23029 5695
rect 23063 5692 23075 5695
rect 23382 5692 23388 5704
rect 23063 5664 23388 5692
rect 23063 5661 23075 5664
rect 23017 5655 23075 5661
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 23750 5692 23756 5704
rect 23711 5664 23756 5692
rect 23750 5652 23756 5664
rect 23808 5652 23814 5704
rect 30009 5695 30067 5701
rect 30009 5661 30021 5695
rect 30055 5692 30067 5695
rect 30282 5692 30288 5704
rect 30055 5664 30288 5692
rect 30055 5661 30067 5664
rect 30009 5655 30067 5661
rect 30282 5652 30288 5664
rect 30340 5652 30346 5704
rect 31202 5652 31208 5704
rect 31260 5692 31266 5704
rect 31665 5695 31723 5701
rect 31665 5692 31677 5695
rect 31260 5664 31677 5692
rect 31260 5652 31266 5664
rect 31665 5661 31677 5664
rect 31711 5661 31723 5695
rect 31665 5655 31723 5661
rect 21082 5584 21088 5636
rect 21140 5624 21146 5636
rect 24762 5624 24768 5636
rect 21140 5596 21574 5624
rect 23400 5596 24768 5624
rect 21140 5584 21146 5596
rect 14608 5528 18184 5556
rect 14608 5516 14614 5528
rect 19242 5516 19248 5568
rect 19300 5556 19306 5568
rect 19429 5559 19487 5565
rect 19429 5556 19441 5559
rect 19300 5528 19441 5556
rect 19300 5516 19306 5528
rect 19429 5525 19441 5528
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 20533 5559 20591 5565
rect 20533 5525 20545 5559
rect 20579 5556 20591 5559
rect 21266 5556 21272 5568
rect 20579 5528 21272 5556
rect 20579 5525 20591 5528
rect 20533 5519 20591 5525
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 21726 5516 21732 5568
rect 21784 5556 21790 5568
rect 23400 5556 23428 5596
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 25498 5584 25504 5636
rect 25556 5584 25562 5636
rect 25958 5584 25964 5636
rect 26016 5624 26022 5636
rect 26053 5627 26111 5633
rect 26053 5624 26065 5627
rect 26016 5596 26065 5624
rect 26016 5584 26022 5596
rect 26053 5593 26065 5596
rect 26099 5593 26111 5627
rect 26053 5587 26111 5593
rect 23566 5556 23572 5568
rect 21784 5528 23428 5556
rect 23527 5528 23572 5556
rect 21784 5516 21790 5528
rect 23566 5516 23572 5528
rect 23624 5516 23630 5568
rect 27338 5556 27344 5568
rect 27299 5528 27344 5556
rect 27338 5516 27344 5528
rect 27396 5516 27402 5568
rect 29178 5516 29184 5568
rect 29236 5556 29242 5568
rect 29917 5559 29975 5565
rect 29917 5556 29929 5559
rect 29236 5528 29929 5556
rect 29236 5516 29242 5528
rect 29917 5525 29929 5528
rect 29963 5525 29975 5559
rect 29917 5519 29975 5525
rect 1104 5466 36892 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 36892 5466
rect 1104 5392 36892 5414
rect 1762 5352 1768 5364
rect 1723 5324 1768 5352
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11698 5352 11704 5364
rect 11112 5324 11704 5352
rect 11112 5312 11118 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 12066 5312 12072 5364
rect 12124 5352 12130 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 12124 5324 12265 5352
rect 12124 5312 12130 5324
rect 12253 5321 12265 5324
rect 12299 5321 12311 5355
rect 15746 5352 15752 5364
rect 12253 5315 12311 5321
rect 13648 5324 15752 5352
rect 9766 5284 9772 5296
rect 9727 5256 9772 5284
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 13648 5284 13676 5324
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16206 5352 16212 5364
rect 16167 5324 16212 5352
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 26329 5355 26387 5361
rect 18012 5324 22094 5352
rect 18012 5312 18018 5324
rect 13294 5256 13676 5284
rect 13725 5287 13783 5293
rect 13725 5253 13737 5287
rect 13771 5284 13783 5287
rect 14366 5284 14372 5296
rect 13771 5256 14372 5284
rect 13771 5253 13783 5256
rect 13725 5247 13783 5253
rect 14366 5244 14372 5256
rect 14424 5244 14430 5296
rect 14458 5244 14464 5296
rect 14516 5244 14522 5296
rect 14737 5287 14795 5293
rect 14737 5253 14749 5287
rect 14783 5284 14795 5287
rect 14826 5284 14832 5296
rect 14783 5256 14832 5284
rect 14783 5253 14795 5256
rect 14737 5247 14795 5253
rect 14826 5244 14832 5256
rect 14884 5244 14890 5296
rect 16482 5284 16488 5296
rect 15962 5256 16488 5284
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 18141 5287 18199 5293
rect 18141 5253 18153 5287
rect 18187 5284 18199 5287
rect 18506 5284 18512 5296
rect 18187 5256 18512 5284
rect 18187 5253 18199 5256
rect 18141 5247 18199 5253
rect 18506 5244 18512 5256
rect 18564 5244 18570 5296
rect 21726 5284 21732 5296
rect 20470 5256 21732 5284
rect 21726 5244 21732 5256
rect 21784 5244 21790 5296
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1636 5188 1685 5216
rect 1636 5176 1642 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14476 5216 14504 5244
rect 14056 5188 14504 5216
rect 14056 5176 14062 5188
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 16172 5188 17233 5216
rect 16172 5176 16178 5188
rect 17221 5185 17233 5188
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 17586 5176 17592 5228
rect 17644 5216 17650 5228
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 17644 5188 18981 5216
rect 17644 5176 17650 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 20993 5219 21051 5225
rect 20993 5185 21005 5219
rect 21039 5216 21051 5219
rect 21910 5216 21916 5228
rect 21039 5188 21916 5216
rect 21039 5185 21051 5188
rect 20993 5179 21051 5185
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 22066 5216 22094 5324
rect 24872 5324 26188 5352
rect 23198 5244 23204 5296
rect 23256 5284 23262 5296
rect 24872 5284 24900 5324
rect 23256 5256 24900 5284
rect 23256 5244 23262 5256
rect 25866 5244 25872 5296
rect 25924 5244 25930 5296
rect 26160 5284 26188 5324
rect 26329 5321 26341 5355
rect 26375 5352 26387 5355
rect 26418 5352 26424 5364
rect 26375 5324 26424 5352
rect 26375 5321 26387 5324
rect 26329 5315 26387 5321
rect 26418 5312 26424 5324
rect 26476 5352 26482 5364
rect 27062 5352 27068 5364
rect 26476 5324 27068 5352
rect 26476 5312 26482 5324
rect 27062 5312 27068 5324
rect 27120 5312 27126 5364
rect 26878 5284 26884 5296
rect 26160 5256 26884 5284
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 30098 5284 30104 5296
rect 27816 5256 30104 5284
rect 24578 5216 24584 5228
rect 22066 5188 22402 5216
rect 24539 5188 24584 5216
rect 24578 5176 24584 5188
rect 24636 5176 24642 5228
rect 26234 5176 26240 5228
rect 26292 5216 26298 5228
rect 27816 5216 27844 5256
rect 30098 5244 30104 5256
rect 30156 5244 30162 5296
rect 26292 5188 27844 5216
rect 26292 5176 26298 5188
rect 27890 5176 27896 5228
rect 27948 5216 27954 5228
rect 29089 5219 29147 5225
rect 29089 5216 29101 5219
rect 27948 5188 29101 5216
rect 27948 5176 27954 5188
rect 29089 5185 29101 5188
rect 29135 5216 29147 5219
rect 30006 5216 30012 5228
rect 29135 5188 30012 5216
rect 29135 5185 29147 5188
rect 29089 5179 29147 5185
rect 30006 5176 30012 5188
rect 30064 5176 30070 5228
rect 36081 5219 36139 5225
rect 36081 5185 36093 5219
rect 36127 5216 36139 5219
rect 36170 5216 36176 5228
rect 36127 5188 36176 5216
rect 36127 5185 36139 5188
rect 36081 5179 36139 5185
rect 36170 5176 36176 5188
rect 36228 5176 36234 5228
rect 9674 5148 9680 5160
rect 9635 5120 9680 5148
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9916 5120 9965 5148
rect 9916 5108 9922 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 19291 5120 20668 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 11149 5083 11207 5089
rect 11149 5049 11161 5083
rect 11195 5080 11207 5083
rect 11195 5052 12434 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 12406 5012 12434 5052
rect 13538 5012 13544 5024
rect 12406 4984 13544 5012
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 14476 5012 14504 5111
rect 15838 5040 15844 5092
rect 15896 5080 15902 5092
rect 16390 5080 16396 5092
rect 15896 5052 16396 5080
rect 15896 5040 15902 5052
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 16666 5040 16672 5092
rect 16724 5080 16730 5092
rect 20640 5080 20668 5120
rect 21634 5108 21640 5160
rect 21692 5148 21698 5160
rect 23477 5151 23535 5157
rect 23477 5148 23489 5151
rect 21692 5120 23489 5148
rect 21692 5108 21698 5120
rect 23477 5117 23489 5120
rect 23523 5117 23535 5151
rect 23753 5151 23811 5157
rect 23753 5148 23765 5151
rect 23477 5111 23535 5117
rect 23676 5120 23765 5148
rect 16724 5052 18644 5080
rect 20640 5052 22508 5080
rect 16724 5040 16730 5052
rect 15746 5012 15752 5024
rect 14476 4984 15752 5012
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 18616 5012 18644 5052
rect 21450 5012 21456 5024
rect 18616 4984 21456 5012
rect 21450 4972 21456 4984
rect 21508 5012 21514 5024
rect 22005 5015 22063 5021
rect 22005 5012 22017 5015
rect 21508 4984 22017 5012
rect 21508 4972 21514 4984
rect 22005 4981 22017 4984
rect 22051 4981 22063 5015
rect 22480 5012 22508 5052
rect 23106 5012 23112 5024
rect 22480 4984 23112 5012
rect 22005 4975 22063 4981
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 23382 4972 23388 5024
rect 23440 5012 23446 5024
rect 23676 5012 23704 5120
rect 23753 5117 23765 5120
rect 23799 5117 23811 5151
rect 23753 5111 23811 5117
rect 24857 5151 24915 5157
rect 24857 5117 24869 5151
rect 24903 5148 24915 5151
rect 26786 5148 26792 5160
rect 24903 5120 26792 5148
rect 24903 5117 24915 5120
rect 24857 5111 24915 5117
rect 26786 5108 26792 5120
rect 26844 5148 26850 5160
rect 27157 5151 27215 5157
rect 27157 5148 27169 5151
rect 26844 5120 27169 5148
rect 26844 5108 26850 5120
rect 27157 5117 27169 5120
rect 27203 5117 27215 5151
rect 27157 5111 27215 5117
rect 27246 5108 27252 5160
rect 27304 5148 27310 5160
rect 27801 5151 27859 5157
rect 27801 5148 27813 5151
rect 27304 5120 27813 5148
rect 27304 5108 27310 5120
rect 27801 5117 27813 5120
rect 27847 5148 27859 5151
rect 28810 5148 28816 5160
rect 27847 5120 28816 5148
rect 27847 5117 27859 5120
rect 27801 5111 27859 5117
rect 28810 5108 28816 5120
rect 28868 5108 28874 5160
rect 36354 5148 36360 5160
rect 36315 5120 36360 5148
rect 36354 5108 36360 5120
rect 36412 5108 36418 5160
rect 28718 5080 28724 5092
rect 25884 5052 28724 5080
rect 23440 4984 23704 5012
rect 23440 4972 23446 4984
rect 24302 4972 24308 5024
rect 24360 5012 24366 5024
rect 25884 5012 25912 5052
rect 28718 5040 28724 5052
rect 28776 5040 28782 5092
rect 29454 5080 29460 5092
rect 28828 5052 29460 5080
rect 24360 4984 25912 5012
rect 24360 4972 24366 4984
rect 25958 4972 25964 5024
rect 26016 5012 26022 5024
rect 28828 5012 28856 5052
rect 29454 5040 29460 5052
rect 29512 5040 29518 5092
rect 28994 5012 29000 5024
rect 26016 4984 28856 5012
rect 28955 4984 29000 5012
rect 26016 4972 26022 4984
rect 28994 4972 29000 4984
rect 29052 4972 29058 5024
rect 1104 4922 36892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36892 4922
rect 1104 4848 36892 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 9122 4808 9128 4820
rect 9083 4780 9128 4808
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9766 4808 9772 4820
rect 9727 4780 9772 4808
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10413 4811 10471 4817
rect 10413 4777 10425 4811
rect 10459 4808 10471 4811
rect 11330 4808 11336 4820
rect 10459 4780 11336 4808
rect 10459 4777 10471 4780
rect 10413 4771 10471 4777
rect 11330 4768 11336 4780
rect 11388 4808 11394 4820
rect 12158 4808 12164 4820
rect 11388 4780 12164 4808
rect 11388 4768 11394 4780
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12437 4811 12495 4817
rect 12437 4777 12449 4811
rect 12483 4808 12495 4811
rect 13998 4808 14004 4820
rect 12483 4780 14004 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 17402 4808 17408 4820
rect 14568 4780 17408 4808
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 14568 4681 14596 4780
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 18782 4808 18788 4820
rect 18743 4780 18788 4808
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 20714 4808 20720 4820
rect 19812 4780 20720 4808
rect 15197 4743 15255 4749
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 15470 4740 15476 4752
rect 15243 4712 15476 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18141 4743 18199 4749
rect 18141 4740 18153 4743
rect 18104 4712 18153 4740
rect 18104 4700 18110 4712
rect 18141 4709 18153 4712
rect 18187 4709 18199 4743
rect 18141 4703 18199 4709
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 11756 4644 14565 4672
rect 11756 4632 11762 4644
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 13740 4613 13768 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9180 4576 9873 4604
rect 9180 4564 9186 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 13725 4607 13783 4613
rect 11471 4576 11836 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 10965 4539 11023 4545
rect 10965 4505 10977 4539
rect 11011 4536 11023 4539
rect 11808 4536 11836 4576
rect 13725 4573 13737 4607
rect 13771 4573 13783 4607
rect 15488 4604 15516 4700
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 16448 4644 17693 4672
rect 16448 4632 16454 4644
rect 17681 4641 17693 4644
rect 17727 4672 17739 4675
rect 17862 4672 17868 4684
rect 17727 4644 17868 4672
rect 17727 4641 17739 4644
rect 17681 4635 17739 4641
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 15488 4576 15700 4604
rect 13725 4567 13783 4573
rect 15562 4536 15568 4548
rect 11011 4508 11652 4536
rect 11808 4508 15568 4536
rect 11011 4505 11023 4508
rect 10965 4499 11023 4505
rect 11624 4468 11652 4508
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 15672 4536 15700 4576
rect 17034 4564 17040 4616
rect 17092 4564 17098 4616
rect 15930 4536 15936 4548
rect 15672 4508 15936 4536
rect 15930 4496 15936 4508
rect 15988 4496 15994 4548
rect 18156 4536 18184 4703
rect 18230 4700 18236 4752
rect 18288 4740 18294 4752
rect 19812 4740 19840 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 24302 4808 24308 4820
rect 21100 4780 24308 4808
rect 18288 4712 19840 4740
rect 18288 4700 18294 4712
rect 18782 4632 18788 4684
rect 18840 4672 18846 4684
rect 19610 4672 19616 4684
rect 18840 4644 19616 4672
rect 18840 4632 18846 4644
rect 19610 4632 19616 4644
rect 19668 4632 19674 4684
rect 19981 4675 20039 4681
rect 19981 4641 19993 4675
rect 20027 4672 20039 4675
rect 20070 4672 20076 4684
rect 20027 4644 20076 4672
rect 20027 4641 20039 4644
rect 19981 4635 20039 4641
rect 20070 4632 20076 4644
rect 20128 4672 20134 4684
rect 20714 4672 20720 4684
rect 20128 4644 20720 4672
rect 20128 4632 20134 4644
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 19058 4564 19064 4616
rect 19116 4604 19122 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19116 4576 19717 4604
rect 19116 4564 19122 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 21100 4590 21128 4780
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 28994 4808 29000 4820
rect 24412 4780 29000 4808
rect 21468 4712 22094 4740
rect 19705 4567 19763 4573
rect 18156 4508 19748 4536
rect 14918 4468 14924 4480
rect 11624 4440 14924 4468
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15838 4428 15844 4480
rect 15896 4468 15902 4480
rect 18690 4468 18696 4480
rect 15896 4440 18696 4468
rect 15896 4428 15902 4440
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 19720 4468 19748 4508
rect 21468 4477 21496 4712
rect 22066 4672 22094 4712
rect 24302 4672 24308 4684
rect 22066 4644 24308 4672
rect 24302 4632 24308 4644
rect 24360 4632 24366 4684
rect 22094 4564 22100 4616
rect 22152 4604 22158 4616
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 22152 4576 22293 4604
rect 22152 4564 22158 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 24412 4604 24440 4780
rect 28994 4768 29000 4780
rect 29052 4768 29058 4820
rect 30558 4768 30564 4820
rect 30616 4808 30622 4820
rect 30837 4811 30895 4817
rect 30837 4808 30849 4811
rect 30616 4780 30849 4808
rect 30616 4768 30622 4780
rect 30837 4777 30849 4780
rect 30883 4777 30895 4811
rect 36354 4808 36360 4820
rect 36315 4780 36360 4808
rect 30837 4771 30895 4777
rect 36354 4768 36360 4780
rect 36412 4768 36418 4820
rect 26789 4743 26847 4749
rect 26789 4709 26801 4743
rect 26835 4709 26847 4743
rect 26789 4703 26847 4709
rect 24578 4672 24584 4684
rect 24539 4644 24584 4672
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 24854 4672 24860 4684
rect 24815 4644 24860 4672
rect 24854 4632 24860 4644
rect 24912 4632 24918 4684
rect 26602 4672 26608 4684
rect 25976 4644 26608 4672
rect 23690 4576 24440 4604
rect 25976 4590 26004 4644
rect 26602 4632 26608 4644
rect 26660 4632 26666 4684
rect 26694 4632 26700 4684
rect 26752 4672 26758 4684
rect 26804 4672 26832 4703
rect 26752 4644 26832 4672
rect 26752 4632 26758 4644
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 27028 4644 30788 4672
rect 27028 4632 27034 4644
rect 22281 4567 22339 4573
rect 26510 4564 26516 4616
rect 26568 4604 26574 4616
rect 27525 4607 27583 4613
rect 27525 4604 27537 4607
rect 26568 4576 27537 4604
rect 26568 4564 26574 4576
rect 27525 4573 27537 4576
rect 27571 4573 27583 4607
rect 27525 4567 27583 4573
rect 27614 4564 27620 4616
rect 27672 4564 27678 4616
rect 27798 4564 27804 4616
rect 27856 4604 27862 4616
rect 28353 4607 28411 4613
rect 28353 4604 28365 4607
rect 27856 4576 28365 4604
rect 27856 4564 27862 4576
rect 28353 4573 28365 4576
rect 28399 4604 28411 4607
rect 28626 4604 28632 4616
rect 28399 4576 28632 4604
rect 28399 4573 28411 4576
rect 28353 4567 28411 4573
rect 28626 4564 28632 4576
rect 28684 4564 28690 4616
rect 30760 4613 30788 4644
rect 30745 4607 30803 4613
rect 30745 4573 30757 4607
rect 30791 4573 30803 4607
rect 30745 4567 30803 4573
rect 22557 4539 22615 4545
rect 22557 4536 22569 4539
rect 22066 4508 22569 4536
rect 21453 4471 21511 4477
rect 21453 4468 21465 4471
rect 19720 4440 21465 4468
rect 21453 4437 21465 4440
rect 21499 4437 21511 4471
rect 21453 4431 21511 4437
rect 21542 4428 21548 4480
rect 21600 4468 21606 4480
rect 22066 4468 22094 4508
rect 22557 4505 22569 4508
rect 22603 4536 22615 4539
rect 22830 4536 22836 4548
rect 22603 4508 22836 4536
rect 22603 4505 22615 4508
rect 22557 4499 22615 4505
rect 22830 4496 22836 4508
rect 22888 4496 22894 4548
rect 26234 4496 26240 4548
rect 26292 4536 26298 4548
rect 26973 4539 27031 4545
rect 26973 4536 26985 4539
rect 26292 4508 26985 4536
rect 26292 4496 26298 4508
rect 26973 4505 26985 4508
rect 27019 4536 27031 4539
rect 27338 4536 27344 4548
rect 27019 4508 27344 4536
rect 27019 4505 27031 4508
rect 26973 4499 27031 4505
rect 27338 4496 27344 4508
rect 27396 4496 27402 4548
rect 27632 4536 27660 4564
rect 27540 4508 27660 4536
rect 21600 4440 22094 4468
rect 24029 4471 24087 4477
rect 21600 4428 21606 4440
rect 24029 4437 24041 4471
rect 24075 4468 24087 4471
rect 24118 4468 24124 4480
rect 24075 4440 24124 4468
rect 24075 4437 24087 4440
rect 24029 4431 24087 4437
rect 24118 4428 24124 4440
rect 24176 4428 24182 4480
rect 26329 4471 26387 4477
rect 26329 4437 26341 4471
rect 26375 4468 26387 4471
rect 27540 4468 27568 4508
rect 26375 4440 27568 4468
rect 26375 4437 26387 4440
rect 26329 4431 26387 4437
rect 27614 4428 27620 4480
rect 27672 4468 27678 4480
rect 27709 4471 27767 4477
rect 27709 4468 27721 4471
rect 27672 4440 27721 4468
rect 27672 4428 27678 4440
rect 27709 4437 27721 4440
rect 27755 4437 27767 4471
rect 27709 4431 27767 4437
rect 28718 4428 28724 4480
rect 28776 4468 28782 4480
rect 28813 4471 28871 4477
rect 28813 4468 28825 4471
rect 28776 4440 28825 4468
rect 28776 4428 28782 4440
rect 28813 4437 28825 4440
rect 28859 4437 28871 4471
rect 28813 4431 28871 4437
rect 1104 4378 36892 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 36892 4378
rect 1104 4304 36892 4326
rect 13262 4264 13268 4276
rect 12084 4236 13268 4264
rect 12084 4196 12112 4236
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 15838 4264 15844 4276
rect 14752 4236 15844 4264
rect 11992 4168 12112 4196
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 10778 4128 10784 4140
rect 9447 4100 10784 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 11330 4128 11336 4140
rect 11011 4100 11336 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11992 4128 12020 4168
rect 12231 4156 12237 4208
rect 12289 4205 12295 4208
rect 12289 4196 12298 4205
rect 13538 4196 13544 4208
rect 12289 4168 12334 4196
rect 13451 4168 13544 4196
rect 12289 4159 12298 4168
rect 12289 4156 12295 4159
rect 13538 4156 13544 4168
rect 13596 4196 13602 4208
rect 14752 4196 14780 4236
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16206 4264 16212 4276
rect 16040 4236 16212 4264
rect 13596 4168 14780 4196
rect 13596 4156 13602 4168
rect 15562 4156 15568 4208
rect 15620 4156 15626 4208
rect 16040 4205 16068 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 16908 4236 18644 4264
rect 16908 4224 16914 4236
rect 16025 4199 16083 4205
rect 16025 4165 16037 4199
rect 16071 4165 16083 4199
rect 18506 4196 18512 4208
rect 18354 4168 18512 4196
rect 16025 4159 16083 4165
rect 18506 4156 18512 4168
rect 18564 4156 18570 4208
rect 11440 4100 12020 4128
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 11440 4060 11468 4100
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16850 4128 16856 4140
rect 16356 4100 16401 4128
rect 16811 4100 16856 4128
rect 16356 4088 16362 4100
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 18616 4128 18644 4236
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 21910 4264 21916 4276
rect 18748 4236 21916 4264
rect 18748 4224 18754 4236
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 23382 4264 23388 4276
rect 22520 4236 23388 4264
rect 22520 4224 22526 4236
rect 23382 4224 23388 4236
rect 23440 4264 23446 4276
rect 26510 4264 26516 4276
rect 23440 4236 23796 4264
rect 26471 4236 26516 4264
rect 23440 4224 23446 4236
rect 19337 4199 19395 4205
rect 19337 4165 19349 4199
rect 19383 4196 19395 4199
rect 19426 4196 19432 4208
rect 19383 4168 19432 4196
rect 19383 4165 19395 4168
rect 19337 4159 19395 4165
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 21818 4196 21824 4208
rect 20562 4168 21824 4196
rect 21818 4156 21824 4168
rect 21876 4156 21882 4208
rect 23474 4196 23480 4208
rect 23046 4168 23480 4196
rect 23474 4156 23480 4168
rect 23532 4156 23538 4208
rect 19058 4128 19064 4140
rect 18616 4100 19064 4128
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 20990 4088 20996 4140
rect 21048 4128 21054 4140
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 21048 4100 21097 4128
rect 21048 4088 21054 4100
rect 21085 4097 21097 4100
rect 21131 4128 21143 4131
rect 21542 4128 21548 4140
rect 21131 4100 21548 4128
rect 21131 4097 21143 4100
rect 21085 4091 21143 4097
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 23768 4137 23796 4236
rect 26510 4224 26516 4236
rect 26568 4224 26574 4276
rect 26602 4224 26608 4276
rect 26660 4264 26666 4276
rect 31386 4264 31392 4276
rect 26660 4236 31392 4264
rect 26660 4224 26666 4236
rect 31386 4224 31392 4236
rect 31444 4224 31450 4276
rect 26050 4196 26056 4208
rect 25714 4168 26056 4196
rect 26050 4156 26056 4168
rect 26108 4156 26114 4208
rect 29638 4196 29644 4208
rect 28198 4168 29644 4196
rect 29638 4156 29644 4168
rect 29696 4156 29702 4208
rect 31754 4196 31760 4208
rect 30116 4168 31760 4196
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23799 4100 24225 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 26326 4088 26332 4140
rect 26384 4128 26390 4140
rect 26421 4131 26479 4137
rect 26421 4128 26433 4131
rect 26384 4100 26433 4128
rect 26384 4088 26390 4100
rect 26421 4097 26433 4100
rect 26467 4097 26479 4131
rect 26421 4091 26479 4097
rect 28905 4131 28963 4137
rect 28905 4097 28917 4131
rect 28951 4128 28963 4131
rect 28994 4128 29000 4140
rect 28951 4100 29000 4128
rect 28951 4097 28963 4100
rect 28905 4091 28963 4097
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 30006 4128 30012 4140
rect 29919 4100 30012 4128
rect 30006 4088 30012 4100
rect 30064 4128 30070 4140
rect 30116 4128 30144 4168
rect 31754 4156 31760 4168
rect 31812 4156 31818 4208
rect 30742 4128 30748 4140
rect 30064 4100 30144 4128
rect 30655 4100 30748 4128
rect 30064 4088 30070 4100
rect 30742 4088 30748 4100
rect 30800 4128 30806 4140
rect 31389 4131 31447 4137
rect 31389 4128 31401 4131
rect 30800 4100 31401 4128
rect 30800 4088 30806 4100
rect 31389 4097 31401 4100
rect 31435 4097 31447 4131
rect 31389 4091 31447 4097
rect 11974 4060 11980 4072
rect 10551 4032 11468 4060
rect 11935 4032 11980 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 13446 4060 13452 4072
rect 12084 4032 13452 4060
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 11238 3992 11244 4004
rect 9999 3964 11244 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 11238 3952 11244 3964
rect 11296 3992 11302 4004
rect 12084 3992 12112 4032
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 13872 4032 14565 4060
rect 13872 4020 13878 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 17126 4060 17132 4072
rect 14553 4023 14611 4029
rect 15028 4032 16988 4060
rect 17087 4032 17132 4060
rect 11296 3964 12112 3992
rect 11296 3952 11302 3964
rect 14458 3952 14464 4004
rect 14516 3992 14522 4004
rect 15028 3992 15056 4032
rect 14516 3964 15056 3992
rect 14516 3952 14522 3964
rect 11057 3927 11115 3933
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 13630 3924 13636 3936
rect 11103 3896 13636 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 13780 3896 13825 3924
rect 13780 3884 13786 3896
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 16758 3924 16764 3936
rect 14608 3896 16764 3924
rect 14608 3884 14614 3896
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 16960 3924 16988 4032
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4060 18659 4063
rect 20898 4060 20904 4072
rect 18647 4032 20904 4060
rect 18647 4029 18659 4032
rect 18601 4023 18659 4029
rect 20898 4020 20904 4032
rect 20956 4020 20962 4072
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4060 23535 4063
rect 23523 4032 23704 4060
rect 23523 4029 23535 4032
rect 23477 4023 23535 4029
rect 18524 3964 18736 3992
rect 18524 3924 18552 3964
rect 16960 3896 18552 3924
rect 18708 3924 18736 3964
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 21818 3992 21824 4004
rect 20772 3964 21824 3992
rect 20772 3952 20778 3964
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 23676 3992 23704 4032
rect 23842 4020 23848 4072
rect 23900 4060 23906 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 23900 4032 24501 4060
rect 23900 4020 23906 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 25038 4020 25044 4072
rect 25096 4060 25102 4072
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25096 4032 25973 4060
rect 25096 4020 25102 4032
rect 25961 4029 25973 4032
rect 26007 4060 26019 4063
rect 26050 4060 26056 4072
rect 26007 4032 26056 4060
rect 26007 4029 26019 4032
rect 25961 4023 26019 4029
rect 26050 4020 26056 4032
rect 26108 4020 26114 4072
rect 26878 4020 26884 4072
rect 26936 4060 26942 4072
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 26936 4032 27169 4060
rect 26936 4020 26942 4032
rect 27157 4029 27169 4032
rect 27203 4029 27215 4063
rect 28534 4060 28540 4072
rect 27157 4023 27215 4029
rect 27632 4032 28540 4060
rect 23676 3964 24348 3992
rect 22005 3927 22063 3933
rect 22005 3924 22017 3927
rect 18708 3896 22017 3924
rect 22005 3893 22017 3896
rect 22051 3924 22063 3927
rect 23382 3924 23388 3936
rect 22051 3896 23388 3924
rect 22051 3893 22063 3896
rect 22005 3887 22063 3893
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 24320 3924 24348 3964
rect 25866 3952 25872 4004
rect 25924 3992 25930 4004
rect 27632 3992 27660 4032
rect 28534 4020 28540 4032
rect 28592 4020 28598 4072
rect 28626 4020 28632 4072
rect 28684 4060 28690 4072
rect 28684 4032 28948 4060
rect 28684 4020 28690 4032
rect 25924 3964 27660 3992
rect 28920 3992 28948 4032
rect 30466 3992 30472 4004
rect 28920 3964 30472 3992
rect 25924 3952 25930 3964
rect 30466 3952 30472 3964
rect 30524 3952 30530 4004
rect 35894 3952 35900 4004
rect 35952 3992 35958 4004
rect 35952 3964 35997 3992
rect 35952 3952 35958 3964
rect 26418 3924 26424 3936
rect 24320 3896 26424 3924
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 26786 3884 26792 3936
rect 26844 3924 26850 3936
rect 28994 3924 29000 3936
rect 26844 3896 29000 3924
rect 26844 3884 26850 3896
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 29546 3884 29552 3936
rect 29604 3924 29610 3936
rect 29917 3927 29975 3933
rect 29917 3924 29929 3927
rect 29604 3896 29929 3924
rect 29604 3884 29610 3896
rect 29917 3893 29929 3896
rect 29963 3893 29975 3927
rect 29917 3887 29975 3893
rect 31205 3927 31263 3933
rect 31205 3893 31217 3927
rect 31251 3924 31263 3927
rect 31294 3924 31300 3936
rect 31251 3896 31300 3924
rect 31251 3893 31263 3896
rect 31205 3887 31263 3893
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 1104 3834 36892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36892 3834
rect 1104 3760 36892 3782
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 11606 3720 11612 3732
rect 9815 3692 11612 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12434 3720 12440 3732
rect 11808 3692 12440 3720
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 11808 3584 11836 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 13780 3692 18460 3720
rect 13780 3680 13786 3692
rect 13630 3612 13636 3664
rect 13688 3652 13694 3664
rect 13688 3624 15056 3652
rect 13688 3612 13694 3624
rect 11287 3556 11836 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 11940 3556 12265 3584
rect 11940 3544 11946 3556
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3584 14427 3587
rect 14550 3584 14556 3596
rect 14415 3556 14556 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 7834 3516 7840 3528
rect 1903 3488 7840 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 9324 3448 9352 3479
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11974 3516 11980 3528
rect 11572 3488 11980 3516
rect 11572 3476 11578 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 14182 3516 14188 3528
rect 13386 3488 14188 3516
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14921 3519 14979 3525
rect 14332 3488 14377 3516
rect 14332 3476 14338 3488
rect 14921 3485 14933 3519
rect 14967 3516 14979 3519
rect 15028 3516 15056 3624
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 16850 3584 16856 3596
rect 15160 3556 16856 3584
rect 15160 3544 15166 3556
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18322 3584 18328 3596
rect 18095 3556 18328 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 14967 3488 15056 3516
rect 14967 3485 14979 3488
rect 14921 3479 14979 3485
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15896 3488 16037 3516
rect 15896 3476 15902 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16025 3479 16083 3485
rect 5592 3420 9352 3448
rect 5592 3408 5598 3420
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 2406 3380 2412 3392
rect 2367 3352 2412 3380
rect 2406 3340 2412 3352
rect 2464 3340 2470 3392
rect 8570 3380 8576 3392
rect 8531 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9122 3380 9128 3392
rect 9083 3352 9128 3380
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9324 3380 9352 3420
rect 10778 3408 10784 3460
rect 10836 3408 10842 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 15010 3448 15016 3460
rect 11204 3420 12296 3448
rect 11204 3408 11210 3420
rect 11790 3380 11796 3392
rect 9324 3352 11796 3380
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 12268 3380 12296 3420
rect 13740 3420 15016 3448
rect 13740 3389 13768 3420
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 15286 3408 15292 3460
rect 15344 3448 15350 3460
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 15344 3420 16313 3448
rect 15344 3408 15350 3420
rect 16301 3417 16313 3420
rect 16347 3417 16359 3451
rect 18432 3448 18460 3692
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 22186 3720 22192 3732
rect 19116 3692 22192 3720
rect 19116 3680 19122 3692
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 22554 3680 22560 3732
rect 22612 3720 22618 3732
rect 23566 3720 23572 3732
rect 22612 3692 23572 3720
rect 22612 3680 22618 3692
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 26326 3720 26332 3732
rect 24636 3692 26332 3720
rect 24636 3680 24642 3692
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 26418 3680 26424 3732
rect 26476 3720 26482 3732
rect 27614 3720 27620 3732
rect 26476 3692 27620 3720
rect 26476 3680 26482 3692
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 27706 3680 27712 3732
rect 27764 3720 27770 3732
rect 28534 3720 28540 3732
rect 27764 3692 28120 3720
rect 28495 3692 28540 3720
rect 27764 3680 27770 3692
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 18748 3624 19441 3652
rect 18748 3612 18754 3624
rect 19429 3621 19441 3624
rect 19475 3652 19487 3655
rect 19794 3652 19800 3664
rect 19475 3624 19800 3652
rect 19475 3621 19487 3624
rect 19429 3615 19487 3621
rect 19794 3612 19800 3624
rect 19852 3612 19858 3664
rect 19978 3652 19984 3664
rect 19939 3624 19984 3652
rect 19978 3612 19984 3624
rect 20036 3612 20042 3664
rect 28092 3652 28120 3692
rect 28534 3680 28540 3692
rect 28592 3720 28598 3732
rect 31202 3720 31208 3732
rect 28592 3692 31208 3720
rect 28592 3680 28598 3692
rect 31202 3680 31208 3692
rect 31260 3680 31266 3732
rect 31386 3720 31392 3732
rect 31347 3692 31392 3720
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 32030 3720 32036 3732
rect 31991 3692 32036 3720
rect 32030 3680 32036 3692
rect 32088 3680 32094 3732
rect 29730 3652 29736 3664
rect 28092 3624 29736 3652
rect 29730 3612 29736 3624
rect 29788 3612 29794 3664
rect 29917 3655 29975 3661
rect 29917 3621 29929 3655
rect 29963 3652 29975 3655
rect 35342 3652 35348 3664
rect 29963 3624 35348 3652
rect 29963 3621 29975 3624
rect 29917 3615 29975 3621
rect 35342 3612 35348 3624
rect 35400 3612 35406 3664
rect 21082 3584 21088 3596
rect 19260 3556 21088 3584
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3510 18935 3519
rect 19260 3516 19288 3556
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3584 21787 3587
rect 22094 3584 22100 3596
rect 21775 3556 22100 3584
rect 21775 3553 21787 3556
rect 21729 3547 21787 3553
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 24578 3584 24584 3596
rect 22244 3556 22289 3584
rect 24539 3556 24584 3584
rect 22244 3544 22250 3556
rect 24578 3544 24584 3556
rect 24636 3544 24642 3596
rect 24854 3584 24860 3596
rect 24815 3556 24860 3584
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 25222 3544 25228 3596
rect 25280 3584 25286 3596
rect 25866 3584 25872 3596
rect 25280 3556 25872 3584
rect 25280 3544 25286 3556
rect 25866 3544 25872 3556
rect 25924 3544 25930 3596
rect 32490 3584 32496 3596
rect 25976 3556 31156 3584
rect 18984 3510 19288 3516
rect 18923 3488 19288 3510
rect 18923 3485 19012 3488
rect 18877 3482 19012 3485
rect 18877 3479 18935 3482
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19392 3488 20378 3516
rect 19392 3476 19398 3488
rect 21818 3476 21824 3528
rect 21876 3516 21882 3528
rect 21876 3488 22094 3516
rect 25976 3502 26004 3556
rect 21876 3476 21882 3488
rect 21450 3448 21456 3460
rect 17526 3420 18000 3448
rect 18432 3420 20208 3448
rect 21411 3420 21456 3448
rect 16301 3411 16359 3417
rect 13725 3383 13783 3389
rect 13725 3380 13737 3383
rect 12268 3352 13737 3380
rect 13725 3349 13737 3352
rect 13771 3349 13783 3383
rect 13725 3343 13783 3349
rect 14826 3340 14832 3392
rect 14884 3380 14890 3392
rect 15105 3383 15163 3389
rect 15105 3380 15117 3383
rect 14884 3352 15117 3380
rect 14884 3340 14890 3352
rect 15105 3349 15117 3352
rect 15151 3349 15163 3383
rect 17972 3380 18000 3420
rect 18598 3380 18604 3392
rect 17972 3352 18604 3380
rect 15105 3343 15163 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 18693 3383 18751 3389
rect 18693 3349 18705 3383
rect 18739 3380 18751 3383
rect 19334 3380 19340 3392
rect 18739 3352 19340 3380
rect 18739 3349 18751 3352
rect 18693 3343 18751 3349
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 20180 3380 20208 3420
rect 21450 3408 21456 3420
rect 21508 3408 21514 3460
rect 21726 3380 21732 3392
rect 20180 3352 21732 3380
rect 21726 3340 21732 3352
rect 21784 3340 21790 3392
rect 22066 3380 22094 3488
rect 26326 3476 26332 3528
rect 26384 3516 26390 3528
rect 26786 3516 26792 3528
rect 26384 3488 26792 3516
rect 26384 3476 26390 3488
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 28442 3476 28448 3528
rect 28500 3516 28506 3528
rect 29730 3516 29736 3528
rect 28500 3488 29736 3516
rect 28500 3476 28506 3488
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 29825 3519 29883 3525
rect 29825 3485 29837 3519
rect 29871 3516 29883 3519
rect 29914 3516 29920 3528
rect 29871 3488 29920 3516
rect 29871 3485 29883 3488
rect 29825 3479 29883 3485
rect 29914 3476 29920 3488
rect 29972 3476 29978 3528
rect 22462 3448 22468 3460
rect 22423 3420 22468 3448
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 24394 3448 24400 3460
rect 23690 3420 24400 3448
rect 24394 3408 24400 3420
rect 24452 3408 24458 3460
rect 25130 3448 25136 3460
rect 24688 3420 25136 3448
rect 23937 3383 23995 3389
rect 23937 3380 23949 3383
rect 22066 3352 23949 3380
rect 23937 3349 23949 3352
rect 23983 3349 23995 3383
rect 23937 3343 23995 3349
rect 24302 3340 24308 3392
rect 24360 3380 24366 3392
rect 24688 3380 24716 3420
rect 25130 3408 25136 3420
rect 25188 3408 25194 3460
rect 27062 3408 27068 3460
rect 27120 3448 27126 3460
rect 27338 3448 27344 3460
rect 27120 3420 27344 3448
rect 27120 3408 27126 3420
rect 27338 3408 27344 3420
rect 27396 3408 27402 3460
rect 28350 3448 28356 3460
rect 28290 3420 28356 3448
rect 28350 3408 28356 3420
rect 28408 3408 28414 3460
rect 28810 3408 28816 3460
rect 28868 3448 28874 3460
rect 30469 3451 30527 3457
rect 30469 3448 30481 3451
rect 28868 3420 30481 3448
rect 28868 3408 28874 3420
rect 30469 3417 30481 3420
rect 30515 3417 30527 3451
rect 30469 3411 30527 3417
rect 24360 3352 24716 3380
rect 24360 3340 24366 3352
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 26234 3380 26240 3392
rect 24820 3352 26240 3380
rect 24820 3340 24826 3352
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 26329 3383 26387 3389
rect 26329 3349 26341 3383
rect 26375 3380 26387 3383
rect 26878 3380 26884 3392
rect 26375 3352 26884 3380
rect 26375 3349 26387 3352
rect 26329 3343 26387 3349
rect 26878 3340 26884 3352
rect 26936 3340 26942 3392
rect 28994 3380 29000 3392
rect 28955 3352 29000 3380
rect 28994 3340 29000 3352
rect 29052 3340 29058 3392
rect 29730 3340 29736 3392
rect 29788 3380 29794 3392
rect 31018 3380 31024 3392
rect 29788 3352 31024 3380
rect 29788 3340 29794 3352
rect 31018 3340 31024 3352
rect 31076 3340 31082 3392
rect 31128 3380 31156 3556
rect 32140 3556 32496 3584
rect 31481 3519 31539 3525
rect 31481 3485 31493 3519
rect 31527 3516 31539 3519
rect 31754 3516 31760 3528
rect 31527 3488 31760 3516
rect 31527 3485 31539 3488
rect 31481 3479 31539 3485
rect 31754 3476 31760 3488
rect 31812 3516 31818 3528
rect 32030 3516 32036 3528
rect 31812 3488 32036 3516
rect 31812 3476 31818 3488
rect 32030 3476 32036 3488
rect 32088 3476 32094 3528
rect 32140 3525 32168 3556
rect 32490 3544 32496 3556
rect 32548 3584 32554 3596
rect 32548 3556 35112 3584
rect 32548 3544 32554 3556
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 32214 3476 32220 3528
rect 32272 3516 32278 3528
rect 32769 3519 32827 3525
rect 32769 3516 32781 3519
rect 32272 3488 32781 3516
rect 32272 3476 32278 3488
rect 32769 3485 32781 3488
rect 32815 3516 32827 3519
rect 32950 3516 32956 3528
rect 32815 3488 32956 3516
rect 32815 3485 32827 3488
rect 32769 3479 32827 3485
rect 32950 3476 32956 3488
rect 33008 3476 33014 3528
rect 35084 3525 35112 3556
rect 35069 3519 35127 3525
rect 35069 3485 35081 3519
rect 35115 3485 35127 3519
rect 35069 3479 35127 3485
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 35952 3488 36093 3516
rect 35952 3476 35958 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 31570 3408 31576 3460
rect 31628 3448 31634 3460
rect 35161 3451 35219 3457
rect 35161 3448 35173 3451
rect 31628 3420 35173 3448
rect 31628 3408 31634 3420
rect 35161 3417 35173 3420
rect 35207 3417 35219 3451
rect 35161 3411 35219 3417
rect 32677 3383 32735 3389
rect 32677 3380 32689 3383
rect 31128 3352 32689 3380
rect 32677 3349 32689 3352
rect 32723 3349 32735 3383
rect 36262 3380 36268 3392
rect 36223 3352 36268 3380
rect 32677 3343 32735 3349
rect 36262 3340 36268 3352
rect 36320 3340 36326 3392
rect 1104 3290 36892 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 36892 3290
rect 1104 3216 36892 3238
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 9674 3176 9680 3188
rect 8895 3148 9680 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 15838 3176 15844 3188
rect 11532 3148 15844 3176
rect 11532 3120 11560 3148
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 9401 3111 9459 3117
rect 9401 3108 9413 3111
rect 8628 3080 9413 3108
rect 8628 3068 8634 3080
rect 9401 3077 9413 3080
rect 9447 3108 9459 3111
rect 11054 3108 11060 3120
rect 9447 3080 11060 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 11149 3111 11207 3117
rect 11149 3077 11161 3111
rect 11195 3108 11207 3111
rect 11514 3108 11520 3120
rect 11195 3080 11520 3108
rect 11195 3077 11207 3080
rect 11149 3071 11207 3077
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 12986 3068 12992 3120
rect 13044 3068 13050 3120
rect 13446 3108 13452 3120
rect 13407 3080 13452 3108
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2406 3040 2412 3052
rect 1903 3012 2412 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 2556 3012 8769 3040
rect 2556 3000 2562 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 13740 3049 13768 3148
rect 15838 3136 15844 3148
rect 15896 3176 15902 3188
rect 16298 3176 16304 3188
rect 15896 3148 16304 3176
rect 15896 3136 15902 3148
rect 16298 3136 16304 3148
rect 16356 3176 16362 3188
rect 16356 3148 16528 3176
rect 16356 3136 16362 3148
rect 15010 3068 15016 3120
rect 15068 3068 15074 3120
rect 16025 3111 16083 3117
rect 16025 3077 16037 3111
rect 16071 3108 16083 3111
rect 16390 3108 16396 3120
rect 16071 3080 16396 3108
rect 16071 3077 16083 3080
rect 16025 3071 16083 3077
rect 16390 3068 16396 3080
rect 16448 3068 16454 3120
rect 13725 3043 13783 3049
rect 9640 3012 12296 3040
rect 9640 3000 9646 3012
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 9490 2972 9496 2984
rect 7791 2944 9496 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11940 2944 11989 2972
rect 11940 2932 11946 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 12268 2972 12296 3012
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16500 3040 16528 3148
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 21358 3176 21364 3188
rect 17184 3148 21364 3176
rect 17184 3136 17190 3148
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 21450 3136 21456 3188
rect 21508 3176 21514 3188
rect 21508 3148 22140 3176
rect 21508 3136 21514 3148
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 19058 3108 19064 3120
rect 17920 3080 19064 3108
rect 17920 3068 17926 3080
rect 16850 3040 16856 3052
rect 16347 3012 16528 3040
rect 16811 3012 16856 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 18800 3049 18828 3080
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 20806 3068 20812 3120
rect 20864 3108 20870 3120
rect 22005 3111 22063 3117
rect 22005 3108 22017 3111
rect 20864 3080 22017 3108
rect 20864 3068 20870 3080
rect 22005 3077 22017 3080
rect 22051 3077 22063 3111
rect 22112 3108 22140 3148
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 26602 3176 26608 3188
rect 22244 3148 26608 3176
rect 22244 3136 22250 3148
rect 26602 3136 26608 3148
rect 26660 3136 26666 3188
rect 26786 3136 26792 3188
rect 26844 3176 26850 3188
rect 27433 3179 27491 3185
rect 27433 3176 27445 3179
rect 26844 3148 27445 3176
rect 26844 3136 26850 3148
rect 27433 3145 27445 3148
rect 27479 3145 27491 3179
rect 27433 3139 27491 3145
rect 28350 3136 28356 3188
rect 28408 3176 28414 3188
rect 32398 3176 32404 3188
rect 28408 3148 31754 3176
rect 32359 3148 32404 3176
rect 28408 3136 28414 3148
rect 22462 3108 22468 3120
rect 22112 3080 22468 3108
rect 22005 3071 22063 3077
rect 22462 3068 22468 3080
rect 22520 3068 22526 3120
rect 24854 3108 24860 3120
rect 23322 3080 24860 3108
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 26142 3068 26148 3120
rect 26200 3108 26206 3120
rect 26513 3111 26571 3117
rect 26513 3108 26525 3111
rect 26200 3080 26525 3108
rect 26200 3068 26206 3080
rect 26513 3077 26525 3080
rect 26559 3108 26571 3111
rect 27614 3108 27620 3120
rect 26559 3080 27620 3108
rect 26559 3077 26571 3080
rect 26513 3071 26571 3077
rect 27614 3068 27620 3080
rect 27672 3068 27678 3120
rect 28810 3068 28816 3120
rect 28868 3108 28874 3120
rect 28905 3111 28963 3117
rect 28905 3108 28917 3111
rect 28868 3080 28917 3108
rect 28868 3068 28874 3080
rect 28905 3077 28917 3080
rect 28951 3077 28963 3111
rect 28905 3071 28963 3077
rect 28994 3068 29000 3120
rect 29052 3108 29058 3120
rect 30834 3108 30840 3120
rect 29052 3080 30840 3108
rect 29052 3068 29058 3080
rect 30834 3068 30840 3080
rect 30892 3068 30898 3120
rect 31726 3108 31754 3148
rect 32398 3136 32404 3148
rect 32456 3136 32462 3188
rect 34425 3179 34483 3185
rect 34425 3145 34437 3179
rect 34471 3176 34483 3179
rect 34471 3148 36308 3176
rect 34471 3145 34483 3148
rect 34425 3139 34483 3145
rect 33045 3111 33103 3117
rect 33045 3108 33057 3111
rect 31726 3080 33057 3108
rect 33045 3077 33057 3080
rect 33091 3077 33103 3111
rect 33045 3071 33103 3077
rect 36280 3052 36308 3148
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 16960 3012 18061 3040
rect 16960 2972 16988 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3009 18843 3043
rect 24029 3043 24087 3049
rect 20194 3012 22094 3040
rect 18785 3003 18843 3009
rect 12268 2944 16988 2972
rect 11977 2935 12035 2941
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18748 2944 19073 2972
rect 18748 2932 18754 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20809 2975 20867 2981
rect 20809 2972 20821 2975
rect 19484 2944 20821 2972
rect 19484 2932 19490 2944
rect 20809 2941 20821 2944
rect 20855 2972 20867 2975
rect 21269 2975 21327 2981
rect 21269 2972 21281 2975
rect 20855 2944 21281 2972
rect 20855 2941 20867 2944
rect 20809 2935 20867 2941
rect 21269 2941 21281 2944
rect 21315 2941 21327 2975
rect 22066 2972 22094 3012
rect 24029 3009 24041 3043
rect 24075 3040 24087 3043
rect 24486 3040 24492 3052
rect 24075 3012 24492 3040
rect 24075 3009 24087 3012
rect 24029 3003 24087 3009
rect 24486 3000 24492 3012
rect 24544 3000 24550 3052
rect 29546 3040 29552 3052
rect 25898 3012 29552 3040
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 29638 3000 29644 3052
rect 29696 3040 29702 3052
rect 29733 3043 29791 3049
rect 29733 3040 29745 3043
rect 29696 3012 29745 3040
rect 29696 3000 29702 3012
rect 29733 3009 29745 3012
rect 29779 3040 29791 3043
rect 31205 3043 31263 3049
rect 29779 3012 30420 3040
rect 29779 3009 29791 3012
rect 29733 3003 29791 3009
rect 23753 2975 23811 2981
rect 22066 2944 22784 2972
rect 21269 2935 21327 2941
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2904 8355 2907
rect 22646 2904 22652 2916
rect 8343 2876 12434 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 12406 2848 12434 2876
rect 20088 2876 22652 2904
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 72 2808 1685 2836
rect 72 2796 78 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 1854 2796 1860 2848
rect 1912 2836 1918 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 1912 2808 2329 2836
rect 1912 2796 1918 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2317 2799 2375 2805
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 2961 2839 3019 2845
rect 2961 2836 2973 2839
rect 2832 2808 2973 2836
rect 2832 2796 2838 2808
rect 2961 2805 2973 2808
rect 3007 2805 3019 2839
rect 12406 2808 12440 2848
rect 2961 2799 3019 2805
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 12768 2808 14565 2836
rect 12768 2796 12774 2808
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 14553 2799 14611 2805
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 16356 2808 17049 2836
rect 16356 2796 16362 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 18104 2808 18245 2836
rect 18104 2796 18110 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 20088 2836 20116 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 18656 2808 20116 2836
rect 18656 2796 18662 2808
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 21450 2836 21456 2848
rect 20220 2808 21456 2836
rect 20220 2796 20226 2808
rect 21450 2796 21456 2808
rect 21508 2796 21514 2848
rect 22756 2836 22784 2944
rect 23753 2941 23765 2975
rect 23799 2972 23811 2975
rect 24302 2972 24308 2984
rect 23799 2944 24308 2972
rect 23799 2941 23811 2944
rect 23753 2935 23811 2941
rect 24302 2932 24308 2944
rect 24360 2932 24366 2984
rect 24394 2932 24400 2984
rect 24452 2972 24458 2984
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 24452 2944 24777 2972
rect 24452 2932 24458 2944
rect 24765 2941 24777 2944
rect 24811 2941 24823 2975
rect 24765 2935 24823 2941
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 24912 2944 26464 2972
rect 24912 2932 24918 2944
rect 26436 2904 26464 2944
rect 26602 2932 26608 2984
rect 26660 2972 26666 2984
rect 30009 2975 30067 2981
rect 30009 2972 30021 2975
rect 26660 2944 30021 2972
rect 26660 2932 26666 2944
rect 30009 2941 30021 2944
rect 30055 2941 30067 2975
rect 30392 2972 30420 3012
rect 31205 3009 31217 3043
rect 31251 3040 31263 3043
rect 32493 3043 32551 3049
rect 32493 3040 32505 3043
rect 31251 3012 32505 3040
rect 31251 3009 31263 3012
rect 31205 3003 31263 3009
rect 32493 3009 32505 3012
rect 32539 3009 32551 3043
rect 32950 3040 32956 3052
rect 32911 3012 32956 3040
rect 32493 3003 32551 3009
rect 31757 2975 31815 2981
rect 31757 2972 31769 2975
rect 30392 2944 31769 2972
rect 30009 2935 30067 2941
rect 31757 2941 31769 2944
rect 31803 2941 31815 2975
rect 32508 2972 32536 3003
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 34977 3043 35035 3049
rect 34977 3009 34989 3043
rect 35023 3040 35035 3043
rect 35621 3043 35679 3049
rect 35621 3040 35633 3043
rect 35023 3012 35633 3040
rect 35023 3009 35035 3012
rect 34977 3003 35035 3009
rect 35621 3009 35633 3012
rect 35667 3040 35679 3043
rect 35986 3040 35992 3052
rect 35667 3012 35992 3040
rect 35667 3009 35679 3012
rect 35621 3003 35679 3009
rect 35986 3000 35992 3012
rect 36044 3000 36050 3052
rect 36262 3040 36268 3052
rect 36223 3012 36268 3040
rect 36262 3000 36268 3012
rect 36320 3000 36326 3052
rect 32508 2944 35480 2972
rect 31757 2935 31815 2941
rect 31570 2904 31576 2916
rect 26436 2876 31576 2904
rect 31570 2864 31576 2876
rect 31628 2864 31634 2916
rect 32858 2864 32864 2916
rect 32916 2904 32922 2916
rect 35452 2913 35480 2944
rect 33597 2907 33655 2913
rect 33597 2904 33609 2907
rect 32916 2876 33609 2904
rect 32916 2864 32922 2876
rect 33597 2873 33609 2876
rect 33643 2873 33655 2907
rect 33597 2867 33655 2873
rect 35437 2907 35495 2913
rect 35437 2873 35449 2907
rect 35483 2873 35495 2907
rect 35437 2867 35495 2873
rect 24026 2836 24032 2848
rect 22756 2808 24032 2836
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 30558 2836 30564 2848
rect 27764 2808 30564 2836
rect 27764 2796 27770 2808
rect 30558 2796 30564 2808
rect 30616 2796 30622 2848
rect 31018 2836 31024 2848
rect 30979 2808 31024 2836
rect 31018 2796 31024 2808
rect 31076 2796 31082 2848
rect 31110 2796 31116 2848
rect 31168 2836 31174 2848
rect 36173 2839 36231 2845
rect 36173 2836 36185 2839
rect 31168 2808 36185 2836
rect 31168 2796 31174 2808
rect 36173 2805 36185 2808
rect 36219 2805 36231 2839
rect 36173 2799 36231 2805
rect 1104 2746 36892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36892 2746
rect 1104 2672 36892 2694
rect 2498 2632 2504 2644
rect 2459 2604 2504 2632
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 15896 2604 27292 2632
rect 15896 2592 15902 2604
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 5534 2564 5540 2576
rect 4203 2536 5540 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 24581 2567 24639 2573
rect 24581 2564 24593 2567
rect 16632 2536 19564 2564
rect 16632 2524 16638 2536
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11572 2468 11989 2496
rect 11572 2456 11578 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2496 14611 2499
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 14599 2468 17141 2496
rect 14599 2465 14611 2468
rect 14553 2459 14611 2465
rect 17129 2465 17141 2468
rect 17175 2496 17187 2499
rect 17862 2496 17868 2508
rect 17175 2468 17868 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17862 2456 17868 2468
rect 17920 2496 17926 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 17920 2468 19441 2496
rect 17920 2456 17926 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19536 2496 19564 2536
rect 20732 2536 24593 2564
rect 20732 2496 20760 2536
rect 24581 2533 24593 2536
rect 24627 2533 24639 2567
rect 24581 2527 24639 2533
rect 19536 2468 20760 2496
rect 21453 2499 21511 2505
rect 19429 2459 19487 2465
rect 21453 2465 21465 2499
rect 21499 2496 21511 2499
rect 21910 2496 21916 2508
rect 21499 2468 21916 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 21910 2456 21916 2468
rect 21968 2456 21974 2508
rect 22094 2496 22100 2508
rect 22055 2468 22100 2496
rect 22094 2456 22100 2468
rect 22152 2456 22158 2508
rect 25958 2456 25964 2508
rect 26016 2496 26022 2508
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 26016 2468 26065 2496
rect 26016 2456 26022 2468
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26326 2496 26332 2508
rect 26287 2468 26332 2496
rect 26053 2459 26111 2465
rect 26326 2456 26332 2468
rect 26384 2496 26390 2508
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 26384 2468 27169 2496
rect 26384 2456 26390 2468
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 27264 2496 27292 2604
rect 28626 2592 28632 2644
rect 28684 2632 28690 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 28684 2604 28917 2632
rect 28684 2592 28690 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 34238 2632 34244 2644
rect 34199 2604 34244 2632
rect 28905 2595 28963 2601
rect 34238 2592 34244 2604
rect 34296 2592 34302 2644
rect 29178 2564 29184 2576
rect 28460 2536 29184 2564
rect 28460 2496 28488 2536
rect 29178 2524 29184 2536
rect 29236 2524 29242 2576
rect 27264 2468 28488 2496
rect 27157 2459 27215 2465
rect 28626 2456 28632 2508
rect 28684 2456 28690 2508
rect 28902 2456 28908 2508
rect 28960 2496 28966 2508
rect 30285 2499 30343 2505
rect 30285 2496 30297 2499
rect 28960 2468 30297 2496
rect 28960 2456 28966 2468
rect 30285 2465 30297 2468
rect 30331 2465 30343 2499
rect 30558 2496 30564 2508
rect 30519 2468 30564 2496
rect 30285 2459 30343 2465
rect 30558 2456 30564 2468
rect 30616 2496 30622 2508
rect 32309 2499 32367 2505
rect 32309 2496 32321 2499
rect 30616 2468 32321 2496
rect 30616 2456 30622 2468
rect 32309 2465 32321 2468
rect 32355 2465 32367 2499
rect 32309 2459 32367 2465
rect 1854 2428 1860 2440
rect 1815 2400 1860 2428
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2774 2428 2780 2440
rect 2363 2400 2780 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3344 2400 3985 2428
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3344 2301 3372 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5350 2428 5356 2440
rect 4939 2400 5356 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 9122 2428 9128 2440
rect 8159 2400 9128 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9490 2428 9496 2440
rect 9451 2400 9496 2428
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10502 2428 10508 2440
rect 10459 2400 10508 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 10870 2428 10876 2440
rect 10831 2400 10876 2428
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 16224 2400 19196 2428
rect 9677 2363 9735 2369
rect 9677 2329 9689 2363
rect 9723 2360 9735 2363
rect 10778 2360 10784 2372
rect 9723 2332 10784 2360
rect 9723 2329 9735 2332
rect 9677 2323 9735 2329
rect 10778 2320 10784 2332
rect 10836 2320 10842 2372
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 12253 2363 12311 2369
rect 12253 2360 12265 2363
rect 11664 2332 12265 2360
rect 11664 2320 11670 2332
rect 12253 2329 12265 2332
rect 12299 2329 12311 2363
rect 13630 2360 13636 2372
rect 13478 2332 13636 2360
rect 12253 2323 12311 2329
rect 13630 2320 13636 2332
rect 13688 2320 13694 2372
rect 14458 2320 14464 2372
rect 14516 2360 14522 2372
rect 14829 2363 14887 2369
rect 14829 2360 14841 2363
rect 14516 2332 14841 2360
rect 14516 2320 14522 2332
rect 14829 2329 14841 2332
rect 14875 2329 14887 2363
rect 14829 2323 14887 2329
rect 15838 2320 15844 2372
rect 15896 2320 15902 2372
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4580 2264 4721 2292
rect 4580 2252 4586 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 7374 2292 7380 2304
rect 7335 2264 7380 2292
rect 6733 2255 6791 2261
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2292 10287 2295
rect 10962 2292 10968 2304
rect 10275 2264 10968 2292
rect 10275 2261 10287 2264
rect 10229 2255 10287 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11057 2295 11115 2301
rect 11057 2261 11069 2295
rect 11103 2292 11115 2295
rect 12894 2292 12900 2304
rect 11103 2264 12900 2292
rect 11103 2261 11115 2264
rect 11057 2255 11115 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 13725 2295 13783 2301
rect 13725 2261 13737 2295
rect 13771 2292 13783 2295
rect 16224 2292 16252 2400
rect 19168 2372 19196 2400
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 28644 2428 28672 2456
rect 31294 2428 31300 2440
rect 21232 2400 24978 2428
rect 28644 2400 29224 2428
rect 31255 2400 31300 2428
rect 21232 2388 21238 2400
rect 17402 2360 17408 2372
rect 16316 2332 17408 2360
rect 16316 2301 16344 2332
rect 17402 2320 17408 2332
rect 17460 2320 17466 2372
rect 18877 2363 18935 2369
rect 18877 2329 18889 2363
rect 18923 2329 18935 2363
rect 18877 2323 18935 2329
rect 13771 2264 16252 2292
rect 16301 2295 16359 2301
rect 13771 2261 13783 2264
rect 13725 2255 13783 2261
rect 16301 2261 16313 2295
rect 16347 2261 16359 2295
rect 18892 2292 18920 2323
rect 19150 2320 19156 2372
rect 19208 2360 19214 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19208 2332 19717 2360
rect 19208 2320 19214 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 21082 2360 21088 2372
rect 20930 2332 21088 2360
rect 19705 2323 19763 2329
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 23753 2363 23811 2369
rect 23753 2329 23765 2363
rect 23799 2329 23811 2363
rect 23753 2323 23811 2329
rect 19242 2292 19248 2304
rect 18892 2264 19248 2292
rect 16301 2255 16359 2261
rect 19242 2252 19248 2264
rect 19300 2292 19306 2304
rect 23768 2292 23796 2323
rect 26050 2320 26056 2372
rect 26108 2360 26114 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 26108 2332 27445 2360
rect 26108 2320 26114 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 29086 2360 29092 2372
rect 28658 2332 29092 2360
rect 27433 2323 27491 2329
rect 29086 2320 29092 2332
rect 29144 2320 29150 2372
rect 29196 2360 29224 2400
rect 31294 2388 31300 2400
rect 31352 2388 31358 2440
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32916 2400 32965 2428
rect 32916 2388 32922 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33244 2360 33272 2391
rect 34238 2388 34244 2440
rect 34296 2428 34302 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34296 2400 34897 2428
rect 34296 2388 34302 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35342 2388 35348 2440
rect 35400 2428 35406 2440
rect 36081 2431 36139 2437
rect 36081 2428 36093 2431
rect 35400 2400 36093 2428
rect 35400 2388 35406 2400
rect 36081 2397 36093 2400
rect 36127 2397 36139 2431
rect 36081 2391 36139 2397
rect 29196 2332 33272 2360
rect 28810 2292 28816 2304
rect 19300 2264 28816 2292
rect 19300 2252 19306 2264
rect 28810 2252 28816 2264
rect 28868 2252 28874 2304
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31113 2295 31171 2301
rect 31113 2292 31125 2295
rect 30984 2264 31125 2292
rect 30984 2252 30990 2264
rect 31113 2261 31125 2264
rect 31159 2261 31171 2295
rect 31113 2255 31171 2261
rect 34422 2252 34428 2304
rect 34480 2292 34486 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34480 2264 35081 2292
rect 34480 2252 34486 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36265 2295 36323 2301
rect 36265 2292 36277 2295
rect 36136 2264 36277 2292
rect 36136 2252 36142 2264
rect 36265 2261 36277 2264
rect 36311 2261 36323 2295
rect 36265 2255 36323 2261
rect 1104 2202 36892 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 36892 2202
rect 1104 2128 36892 2150
rect 7374 2048 7380 2100
rect 7432 2088 7438 2100
rect 10870 2088 10876 2100
rect 7432 2060 10876 2088
rect 7432 2048 7438 2060
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 17402 2048 17408 2100
rect 17460 2088 17466 2100
rect 24670 2088 24676 2100
rect 17460 2060 24676 2088
rect 17460 2048 17466 2060
rect 24670 2048 24676 2060
rect 24728 2048 24734 2100
rect 21082 1980 21088 2032
rect 21140 2020 21146 2032
rect 25590 2020 25596 2032
rect 21140 1992 25596 2020
rect 21140 1980 21146 1992
rect 25590 1980 25596 1992
rect 25648 1980 25654 2032
rect 15930 1912 15936 1964
rect 15988 1952 15994 1964
rect 21910 1952 21916 1964
rect 15988 1924 21916 1952
rect 15988 1912 15994 1924
rect 21910 1912 21916 1924
rect 21968 1912 21974 1964
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16120 37408 16172 37460
rect 2412 37315 2464 37324
rect 2412 37281 2421 37315
rect 2421 37281 2455 37315
rect 2455 37281 2464 37315
rect 2412 37272 2464 37281
rect 12440 37272 12492 37324
rect 3516 37204 3568 37256
rect 4620 37204 4672 37256
rect 6460 37204 6512 37256
rect 7656 37204 7708 37256
rect 9680 37204 9732 37256
rect 12072 37204 12124 37256
rect 12900 37204 12952 37256
rect 26424 37408 26476 37460
rect 16672 37272 16724 37324
rect 19340 37272 19392 37324
rect 18512 37204 18564 37256
rect 19984 37204 20036 37256
rect 22008 37247 22060 37256
rect 22008 37213 22017 37247
rect 22017 37213 22051 37247
rect 22051 37213 22060 37247
rect 22008 37204 22060 37213
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 27436 37247 27488 37256
rect 27436 37213 27445 37247
rect 27445 37213 27479 37247
rect 27479 37213 27488 37247
rect 27436 37204 27488 37213
rect 28448 37247 28500 37256
rect 28448 37213 28457 37247
rect 28457 37213 28491 37247
rect 28491 37213 28500 37247
rect 28448 37204 28500 37213
rect 29920 37204 29972 37256
rect 31024 37247 31076 37256
rect 31024 37213 31033 37247
rect 31033 37213 31067 37247
rect 31067 37213 31076 37247
rect 31024 37204 31076 37213
rect 27344 37136 27396 37188
rect 34796 37204 34848 37256
rect 36084 37247 36136 37256
rect 36084 37213 36093 37247
rect 36093 37213 36127 37247
rect 36127 37213 36136 37247
rect 36084 37204 36136 37213
rect 3240 37111 3292 37120
rect 3240 37077 3249 37111
rect 3249 37077 3283 37111
rect 3283 37077 3292 37111
rect 3240 37068 3292 37077
rect 4804 37111 4856 37120
rect 4804 37077 4813 37111
rect 4813 37077 4847 37111
rect 4847 37077 4856 37111
rect 4804 37068 4856 37077
rect 6736 37111 6788 37120
rect 6736 37077 6745 37111
rect 6745 37077 6779 37111
rect 6779 37077 6788 37111
rect 6736 37068 6788 37077
rect 7748 37068 7800 37120
rect 9956 37111 10008 37120
rect 9956 37077 9965 37111
rect 9965 37077 9999 37111
rect 9999 37077 10008 37111
rect 9956 37068 10008 37077
rect 11060 37068 11112 37120
rect 12532 37068 12584 37120
rect 14832 37068 14884 37120
rect 15660 37111 15712 37120
rect 15660 37077 15669 37111
rect 15669 37077 15703 37111
rect 15703 37077 15712 37111
rect 15660 37068 15712 37077
rect 18052 37068 18104 37120
rect 21272 37068 21324 37120
rect 22560 37068 22612 37120
rect 24492 37068 24544 37120
rect 27712 37068 27764 37120
rect 29644 37068 29696 37120
rect 30932 37068 30984 37120
rect 33140 37111 33192 37120
rect 33140 37077 33149 37111
rect 33149 37077 33183 37111
rect 33183 37077 33192 37111
rect 33140 37068 33192 37077
rect 34520 37068 34572 37120
rect 36176 37068 36228 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2780 36864 2832 36916
rect 7656 36907 7708 36916
rect 7656 36873 7665 36907
rect 7665 36873 7699 36907
rect 7699 36873 7708 36907
rect 7656 36864 7708 36873
rect 12072 36907 12124 36916
rect 12072 36873 12081 36907
rect 12081 36873 12115 36907
rect 12115 36873 12124 36907
rect 12072 36864 12124 36873
rect 19340 36907 19392 36916
rect 19340 36873 19349 36907
rect 19349 36873 19383 36907
rect 19383 36873 19392 36907
rect 19340 36864 19392 36873
rect 27344 36907 27396 36916
rect 27344 36873 27353 36907
rect 27353 36873 27387 36907
rect 27387 36873 27396 36907
rect 27344 36864 27396 36873
rect 31024 36864 31076 36916
rect 35532 36907 35584 36916
rect 35532 36873 35541 36907
rect 35541 36873 35575 36907
rect 35575 36873 35584 36907
rect 35532 36864 35584 36873
rect 37372 36864 37424 36916
rect 1308 36796 1360 36848
rect 1952 36728 2004 36780
rect 8300 36728 8352 36780
rect 12532 36728 12584 36780
rect 13176 36728 13228 36780
rect 19984 36728 20036 36780
rect 20260 36728 20312 36780
rect 28356 36728 28408 36780
rect 35992 36728 36044 36780
rect 35900 36660 35952 36712
rect 2596 36592 2648 36644
rect 3516 36567 3568 36576
rect 3516 36533 3525 36567
rect 3525 36533 3559 36567
rect 3559 36533 3568 36567
rect 3516 36524 3568 36533
rect 8300 36567 8352 36576
rect 8300 36533 8309 36567
rect 8309 36533 8343 36567
rect 8343 36533 8352 36567
rect 8300 36524 8352 36533
rect 18512 36567 18564 36576
rect 18512 36533 18521 36567
rect 18521 36533 18555 36567
rect 18555 36533 18564 36567
rect 18512 36524 18564 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1308 36320 1360 36372
rect 35532 36159 35584 36168
rect 35532 36125 35541 36159
rect 35541 36125 35575 36159
rect 35575 36125 35584 36159
rect 35532 36116 35584 36125
rect 35808 36159 35860 36168
rect 35808 36125 35817 36159
rect 35817 36125 35851 36159
rect 35851 36125 35860 36159
rect 35808 36116 35860 36125
rect 1676 36091 1728 36100
rect 1676 36057 1685 36091
rect 1685 36057 1719 36091
rect 1719 36057 1728 36091
rect 1676 36048 1728 36057
rect 17592 35980 17644 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1676 35819 1728 35828
rect 1676 35785 1685 35819
rect 1685 35785 1719 35819
rect 1719 35785 1728 35819
rect 1676 35776 1728 35785
rect 2412 35776 2464 35828
rect 28448 35776 28500 35828
rect 36084 35819 36136 35828
rect 36084 35785 36093 35819
rect 36093 35785 36127 35819
rect 36127 35785 36136 35819
rect 36084 35776 36136 35785
rect 27160 35683 27212 35692
rect 27160 35649 27169 35683
rect 27169 35649 27203 35683
rect 27203 35649 27212 35683
rect 27160 35640 27212 35649
rect 34520 35640 34572 35692
rect 35808 35640 35860 35692
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 22008 35232 22060 35284
rect 7564 35028 7616 35080
rect 1676 34935 1728 34944
rect 1676 34901 1685 34935
rect 1685 34901 1719 34935
rect 1719 34901 1728 34935
rect 1676 34892 1728 34901
rect 26608 35028 26660 35080
rect 36360 35071 36412 35080
rect 36360 35037 36369 35071
rect 36369 35037 36403 35071
rect 36403 35037 36412 35071
rect 36360 35028 36412 35037
rect 24400 34892 24452 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 36360 34731 36412 34740
rect 36360 34697 36369 34731
rect 36369 34697 36403 34731
rect 36403 34697 36412 34731
rect 36360 34688 36412 34697
rect 24400 34484 24452 34536
rect 36084 34484 36136 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 27160 32852 27212 32904
rect 36360 32895 36412 32904
rect 36360 32861 36369 32895
rect 36369 32861 36403 32895
rect 36403 32861 36412 32895
rect 36360 32852 36412 32861
rect 1676 32827 1728 32836
rect 1676 32793 1685 32827
rect 1685 32793 1719 32827
rect 1719 32793 1728 32827
rect 1676 32784 1728 32793
rect 2228 32784 2280 32836
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1676 32555 1728 32564
rect 1676 32521 1685 32555
rect 1685 32521 1719 32555
rect 1719 32521 1728 32555
rect 1676 32512 1728 32521
rect 22744 32512 22796 32564
rect 36360 32555 36412 32564
rect 36360 32521 36369 32555
rect 36369 32521 36403 32555
rect 36403 32521 36412 32555
rect 36360 32512 36412 32521
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 36084 31943 36136 31952
rect 36084 31909 36093 31943
rect 36093 31909 36127 31943
rect 36127 31909 36136 31943
rect 36084 31900 36136 31909
rect 22008 31764 22060 31816
rect 35808 31764 35860 31816
rect 1584 31696 1636 31748
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 35900 31424 35952 31476
rect 1584 31399 1636 31408
rect 1584 31365 1593 31399
rect 1593 31365 1627 31399
rect 1627 31365 1636 31399
rect 1584 31356 1636 31365
rect 29828 31288 29880 31340
rect 29828 31084 29880 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 29920 30311 29972 30320
rect 29920 30277 29929 30311
rect 29929 30277 29963 30311
rect 29963 30277 29972 30311
rect 29920 30268 29972 30277
rect 24124 30200 24176 30252
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 24584 29792 24636 29844
rect 34796 29792 34848 29844
rect 1584 29520 1636 29572
rect 2044 29520 2096 29572
rect 24492 29452 24544 29504
rect 25596 29452 25648 29504
rect 29736 29520 29788 29572
rect 36360 29520 36412 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 36360 29291 36412 29300
rect 36360 29257 36369 29291
rect 36369 29257 36403 29291
rect 36403 29257 36412 29291
rect 36360 29248 36412 29257
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2320 28024 2372 28076
rect 13176 28067 13228 28076
rect 13176 28033 13185 28067
rect 13185 28033 13219 28067
rect 13219 28033 13228 28067
rect 13176 28024 13228 28033
rect 20260 28067 20312 28076
rect 20260 28033 20269 28067
rect 20269 28033 20303 28067
rect 20303 28033 20312 28067
rect 20260 28024 20312 28033
rect 36268 28067 36320 28076
rect 36268 28033 36277 28067
rect 36277 28033 36311 28067
rect 36311 28033 36320 28067
rect 36268 28024 36320 28033
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 14096 27888 14148 27940
rect 35348 27888 35400 27940
rect 2320 27863 2372 27872
rect 2320 27829 2329 27863
rect 2329 27829 2363 27863
rect 2363 27829 2372 27863
rect 2320 27820 2372 27829
rect 21456 27820 21508 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 7564 27591 7616 27600
rect 7564 27557 7573 27591
rect 7573 27557 7607 27591
rect 7607 27557 7616 27591
rect 7564 27548 7616 27557
rect 3516 27480 3568 27532
rect 14464 27412 14516 27464
rect 34520 27412 34572 27464
rect 8116 27319 8168 27328
rect 8116 27285 8125 27319
rect 8125 27285 8159 27319
rect 8159 27285 8168 27319
rect 8116 27276 8168 27285
rect 25504 27276 25556 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 27160 26528 27212 26580
rect 35808 26460 35860 26512
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 2412 26299 2464 26308
rect 2412 26265 2421 26299
rect 2421 26265 2455 26299
rect 2455 26265 2464 26299
rect 2412 26256 2464 26265
rect 21916 26256 21968 26308
rect 1676 26231 1728 26240
rect 1676 26197 1685 26231
rect 1685 26197 1719 26231
rect 1719 26197 1728 26231
rect 1676 26188 1728 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 26608 24760 26660 24812
rect 2412 24556 2464 24608
rect 26608 24599 26660 24608
rect 26608 24565 26617 24599
rect 26617 24565 26651 24599
rect 26651 24565 26660 24599
rect 26608 24556 26660 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 1584 24080 1636 24132
rect 7564 24080 7616 24132
rect 36176 24055 36228 24064
rect 36176 24021 36185 24055
rect 36185 24021 36219 24055
rect 36219 24021 36228 24055
rect 36176 24012 36228 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 24400 23851 24452 23860
rect 24400 23817 24409 23851
rect 24409 23817 24443 23851
rect 24443 23817 24452 23851
rect 24400 23808 24452 23817
rect 24860 23468 24912 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 22008 23196 22060 23248
rect 21456 23171 21508 23180
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 17868 22992 17920 23044
rect 20996 22992 21048 23044
rect 20076 22967 20128 22976
rect 20076 22933 20085 22967
rect 20085 22933 20119 22967
rect 20119 22933 20128 22967
rect 20076 22924 20128 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 2136 22584 2188 22636
rect 1676 22491 1728 22500
rect 1676 22457 1685 22491
rect 1685 22457 1719 22491
rect 1719 22457 1728 22491
rect 1676 22448 1728 22457
rect 19984 22380 20036 22432
rect 26608 22584 26660 22636
rect 32496 22584 32548 22636
rect 36268 22491 36320 22500
rect 36268 22457 36277 22491
rect 36277 22457 36311 22491
rect 36311 22457 36320 22491
rect 36268 22448 36320 22457
rect 23848 22380 23900 22432
rect 26608 22380 26660 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 21456 22040 21508 22092
rect 22836 21904 22888 21956
rect 23572 21904 23624 21956
rect 15292 21836 15344 21888
rect 17592 21836 17644 21888
rect 20720 21836 20772 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 22836 21675 22888 21684
rect 22836 21641 22845 21675
rect 22845 21641 22879 21675
rect 22879 21641 22888 21675
rect 22836 21632 22888 21641
rect 15292 21607 15344 21616
rect 15292 21573 15301 21607
rect 15301 21573 15335 21607
rect 15335 21573 15344 21607
rect 15292 21564 15344 21573
rect 15384 21607 15436 21616
rect 15384 21573 15393 21607
rect 15393 21573 15427 21607
rect 15427 21573 15436 21607
rect 15384 21564 15436 21573
rect 16672 21564 16724 21616
rect 17868 21564 17920 21616
rect 19984 21607 20036 21616
rect 19984 21573 19993 21607
rect 19993 21573 20027 21607
rect 20027 21573 20036 21607
rect 19984 21564 20036 21573
rect 20720 21607 20772 21616
rect 20720 21573 20729 21607
rect 20729 21573 20763 21607
rect 20763 21573 20772 21607
rect 20720 21564 20772 21573
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 21916 21428 21968 21480
rect 23756 21360 23808 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 20812 21335 20864 21344
rect 20812 21301 20821 21335
rect 20821 21301 20855 21335
rect 20855 21301 20864 21335
rect 20812 21292 20864 21301
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 25320 21292 25372 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 20812 21088 20864 21140
rect 34244 21088 34296 21140
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 22284 20884 22336 20936
rect 24952 20927 25004 20936
rect 24952 20893 24961 20927
rect 24961 20893 24995 20927
rect 24995 20893 25004 20927
rect 24952 20884 25004 20893
rect 29828 20884 29880 20936
rect 35900 20884 35952 20936
rect 20904 20859 20956 20868
rect 20904 20825 20913 20859
rect 20913 20825 20947 20859
rect 20947 20825 20956 20859
rect 20904 20816 20956 20825
rect 20996 20859 21048 20868
rect 20996 20825 21005 20859
rect 21005 20825 21039 20859
rect 21039 20825 21048 20859
rect 21548 20859 21600 20868
rect 20996 20816 21048 20825
rect 21548 20825 21557 20859
rect 21557 20825 21591 20859
rect 21591 20825 21600 20859
rect 21548 20816 21600 20825
rect 17224 20748 17276 20800
rect 22744 20748 22796 20800
rect 25228 20748 25280 20800
rect 25872 20748 25924 20800
rect 36268 20791 36320 20800
rect 36268 20757 36277 20791
rect 36277 20757 36311 20791
rect 36311 20757 36320 20791
rect 36268 20748 36320 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 15384 20544 15436 20596
rect 20904 20544 20956 20596
rect 21916 20544 21968 20596
rect 16948 20476 17000 20528
rect 19616 20476 19668 20528
rect 22376 20476 22428 20528
rect 22744 20519 22796 20528
rect 22744 20485 22753 20519
rect 22753 20485 22787 20519
rect 22787 20485 22796 20519
rect 22744 20476 22796 20485
rect 36084 20544 36136 20596
rect 23388 20476 23440 20528
rect 27436 20476 27488 20528
rect 15200 20408 15252 20460
rect 25320 20408 25372 20460
rect 25872 20451 25924 20460
rect 25872 20417 25881 20451
rect 25881 20417 25915 20451
rect 25915 20417 25924 20451
rect 25872 20408 25924 20417
rect 29092 20408 29144 20460
rect 19340 20340 19392 20392
rect 20076 20340 20128 20392
rect 23296 20340 23348 20392
rect 22192 20272 22244 20324
rect 27160 20272 27212 20324
rect 2688 20204 2740 20256
rect 18512 20204 18564 20256
rect 25964 20247 26016 20256
rect 25964 20213 25973 20247
rect 25973 20213 26007 20247
rect 26007 20213 26016 20247
rect 25964 20204 26016 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 14648 19796 14700 19848
rect 25872 20000 25924 20052
rect 22284 19932 22336 19984
rect 25228 19907 25280 19916
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 22100 19839 22152 19848
rect 22100 19805 22109 19839
rect 22109 19805 22143 19839
rect 22143 19805 22152 19839
rect 22100 19796 22152 19805
rect 17960 19728 18012 19780
rect 18696 19728 18748 19780
rect 22284 19728 22336 19780
rect 22928 19728 22980 19780
rect 2136 19660 2188 19712
rect 2320 19660 2372 19712
rect 15292 19660 15344 19712
rect 17684 19703 17736 19712
rect 17684 19669 17693 19703
rect 17693 19669 17727 19703
rect 17727 19669 17736 19703
rect 17684 19660 17736 19669
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 23388 19771 23440 19780
rect 23388 19737 23397 19771
rect 23397 19737 23431 19771
rect 23431 19737 23440 19771
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 23388 19728 23440 19737
rect 23480 19660 23532 19712
rect 24584 19771 24636 19780
rect 24584 19737 24593 19771
rect 24593 19737 24627 19771
rect 24627 19737 24636 19771
rect 24584 19728 24636 19737
rect 25964 19771 26016 19780
rect 25964 19737 25973 19771
rect 25973 19737 26007 19771
rect 26007 19737 26016 19771
rect 25964 19728 26016 19737
rect 27068 19771 27120 19780
rect 27068 19737 27077 19771
rect 27077 19737 27111 19771
rect 27111 19737 27120 19771
rect 27068 19728 27120 19737
rect 27160 19771 27212 19780
rect 27160 19737 27169 19771
rect 27169 19737 27203 19771
rect 27203 19737 27212 19771
rect 27160 19728 27212 19737
rect 27620 19660 27672 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 15476 19456 15528 19508
rect 17316 19431 17368 19440
rect 17316 19397 17325 19431
rect 17325 19397 17359 19431
rect 17359 19397 17368 19431
rect 17316 19388 17368 19397
rect 20996 19456 21048 19508
rect 20904 19388 20956 19440
rect 21456 19388 21508 19440
rect 25504 19388 25556 19440
rect 27068 19456 27120 19508
rect 32496 19499 32548 19508
rect 32496 19465 32505 19499
rect 32505 19465 32539 19499
rect 32539 19465 32548 19499
rect 32496 19456 32548 19465
rect 35900 19388 35952 19440
rect 1584 19320 1636 19372
rect 16028 19320 16080 19372
rect 17040 19320 17092 19372
rect 20628 19320 20680 19372
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 6828 19184 6880 19236
rect 15384 19184 15436 19236
rect 19432 19252 19484 19304
rect 21088 19252 21140 19304
rect 32312 19363 32364 19372
rect 21640 19252 21692 19304
rect 22100 19252 22152 19304
rect 23296 19295 23348 19304
rect 23296 19261 23305 19295
rect 23305 19261 23339 19295
rect 23339 19261 23348 19295
rect 23296 19252 23348 19261
rect 23572 19295 23624 19304
rect 23572 19261 23581 19295
rect 23581 19261 23615 19295
rect 23615 19261 23624 19295
rect 23572 19252 23624 19261
rect 18788 19184 18840 19236
rect 21548 19184 21600 19236
rect 24584 19252 24636 19304
rect 27068 19252 27120 19304
rect 25596 19184 25648 19236
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 36084 19363 36136 19372
rect 36084 19329 36093 19363
rect 36093 19329 36127 19363
rect 36127 19329 36136 19363
rect 36084 19320 36136 19329
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 16120 19116 16172 19168
rect 17960 19116 18012 19168
rect 19156 19116 19208 19168
rect 20076 19116 20128 19168
rect 21272 19116 21324 19168
rect 21364 19116 21416 19168
rect 22560 19116 22612 19168
rect 25872 19116 25924 19168
rect 36268 19159 36320 19168
rect 36268 19125 36277 19159
rect 36277 19125 36311 19159
rect 36311 19125 36320 19159
rect 36268 19116 36320 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 14280 18912 14332 18964
rect 15476 18912 15528 18964
rect 15844 18912 15896 18964
rect 17316 18912 17368 18964
rect 20812 18912 20864 18964
rect 25596 18912 25648 18964
rect 25964 18912 26016 18964
rect 27068 18912 27120 18964
rect 14556 18708 14608 18760
rect 15200 18708 15252 18760
rect 15936 18708 15988 18760
rect 16120 18708 16172 18760
rect 18788 18819 18840 18828
rect 18788 18785 18797 18819
rect 18797 18785 18831 18819
rect 18831 18785 18840 18819
rect 18788 18776 18840 18785
rect 20536 18844 20588 18896
rect 21364 18776 21416 18828
rect 22560 18776 22612 18828
rect 20996 18708 21048 18760
rect 21824 18751 21876 18760
rect 14740 18615 14792 18624
rect 14740 18581 14749 18615
rect 14749 18581 14783 18615
rect 14783 18581 14792 18615
rect 14740 18572 14792 18581
rect 15476 18572 15528 18624
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 17960 18640 18012 18692
rect 19984 18640 20036 18692
rect 21824 18717 21833 18751
rect 21833 18717 21867 18751
rect 21867 18717 21876 18751
rect 21824 18708 21876 18717
rect 22284 18708 22336 18760
rect 26608 18776 26660 18828
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 27160 18751 27212 18760
rect 27160 18717 27169 18751
rect 27169 18717 27203 18751
rect 27203 18717 27212 18751
rect 27160 18708 27212 18717
rect 18328 18572 18380 18624
rect 18604 18572 18656 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 21456 18572 21508 18624
rect 22744 18572 22796 18624
rect 24032 18640 24084 18692
rect 24860 18640 24912 18692
rect 25872 18683 25924 18692
rect 25872 18649 25881 18683
rect 25881 18649 25915 18683
rect 25915 18649 25924 18683
rect 25872 18640 25924 18649
rect 24952 18572 25004 18624
rect 25596 18572 25648 18624
rect 27712 18572 27764 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 14464 18368 14516 18420
rect 15016 18368 15068 18420
rect 14096 18343 14148 18352
rect 14096 18309 14105 18343
rect 14105 18309 14139 18343
rect 14139 18309 14148 18343
rect 14096 18300 14148 18309
rect 15292 18300 15344 18352
rect 15660 18300 15712 18352
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 13268 18071 13320 18080
rect 13268 18037 13277 18071
rect 13277 18037 13311 18071
rect 13311 18037 13320 18071
rect 13268 18028 13320 18037
rect 15108 18164 15160 18216
rect 15384 18164 15436 18216
rect 18788 18368 18840 18420
rect 21640 18368 21692 18420
rect 24032 18411 24084 18420
rect 24032 18377 24041 18411
rect 24041 18377 24075 18411
rect 24075 18377 24084 18411
rect 24032 18368 24084 18377
rect 26700 18368 26752 18420
rect 28816 18368 28868 18420
rect 32312 18368 32364 18420
rect 16764 18300 16816 18352
rect 19432 18300 19484 18352
rect 20260 18343 20312 18352
rect 20260 18309 20269 18343
rect 20269 18309 20303 18343
rect 20303 18309 20312 18343
rect 20260 18300 20312 18309
rect 22192 18300 22244 18352
rect 16396 18232 16448 18284
rect 18604 18232 18656 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 23664 18300 23716 18352
rect 24124 18300 24176 18352
rect 25596 18343 25648 18352
rect 25596 18309 25605 18343
rect 25605 18309 25639 18343
rect 25639 18309 25648 18343
rect 25596 18300 25648 18309
rect 21272 18232 21324 18241
rect 17224 18164 17276 18216
rect 20168 18207 20220 18216
rect 20168 18173 20177 18207
rect 20177 18173 20211 18207
rect 20211 18173 20220 18207
rect 20168 18164 20220 18173
rect 24768 18232 24820 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 23756 18164 23808 18216
rect 24124 18164 24176 18216
rect 24216 18164 24268 18216
rect 25504 18207 25556 18216
rect 25504 18173 25513 18207
rect 25513 18173 25547 18207
rect 25547 18173 25556 18207
rect 25504 18164 25556 18173
rect 27620 18164 27672 18216
rect 18144 18096 18196 18148
rect 18328 18096 18380 18148
rect 25320 18096 25372 18148
rect 15844 18028 15896 18080
rect 16488 18028 16540 18080
rect 18052 18028 18104 18080
rect 20812 18028 20864 18080
rect 22468 18028 22520 18080
rect 22652 18028 22704 18080
rect 27068 18028 27120 18080
rect 27252 18071 27304 18080
rect 27252 18037 27261 18071
rect 27261 18037 27295 18071
rect 27295 18037 27304 18071
rect 27252 18028 27304 18037
rect 28816 18028 28868 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 6368 17824 6420 17876
rect 6828 17824 6880 17876
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 12440 17824 12492 17833
rect 13176 17824 13228 17876
rect 13452 17620 13504 17672
rect 20168 17824 20220 17876
rect 15384 17756 15436 17808
rect 16120 17756 16172 17808
rect 21088 17756 21140 17808
rect 22836 17756 22888 17808
rect 27344 17756 27396 17808
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 15292 17688 15344 17740
rect 17224 17688 17276 17740
rect 19340 17688 19392 17740
rect 20168 17688 20220 17740
rect 22376 17688 22428 17740
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 25780 17688 25832 17740
rect 19156 17620 19208 17672
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 20812 17620 20864 17629
rect 15476 17595 15528 17604
rect 15476 17561 15485 17595
rect 15485 17561 15519 17595
rect 15519 17561 15528 17595
rect 15476 17552 15528 17561
rect 15568 17595 15620 17604
rect 15568 17561 15577 17595
rect 15577 17561 15611 17595
rect 15611 17561 15620 17595
rect 15568 17552 15620 17561
rect 16304 17595 16356 17604
rect 16304 17561 16313 17595
rect 16313 17561 16347 17595
rect 16347 17561 16356 17595
rect 16304 17552 16356 17561
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 16488 17484 16540 17536
rect 17040 17552 17092 17604
rect 18144 17552 18196 17604
rect 18236 17484 18288 17536
rect 19248 17484 19300 17536
rect 20352 17552 20404 17604
rect 21456 17595 21508 17604
rect 21456 17561 21465 17595
rect 21465 17561 21499 17595
rect 21499 17561 21508 17595
rect 21456 17552 21508 17561
rect 23020 17595 23072 17604
rect 23020 17561 23029 17595
rect 23029 17561 23063 17595
rect 23063 17561 23072 17595
rect 23020 17552 23072 17561
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 22100 17484 22152 17536
rect 22376 17484 22428 17536
rect 25596 17552 25648 17604
rect 28356 17824 28408 17876
rect 27896 17756 27948 17808
rect 27712 17688 27764 17740
rect 24308 17484 24360 17536
rect 27528 17552 27580 17604
rect 27712 17595 27764 17604
rect 27712 17561 27721 17595
rect 27721 17561 27755 17595
rect 27755 17561 27764 17595
rect 27712 17552 27764 17561
rect 26608 17484 26660 17536
rect 29000 17484 29052 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 9956 17323 10008 17332
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 11336 17144 11388 17196
rect 16120 17280 16172 17332
rect 16304 17280 16356 17332
rect 16948 17323 17000 17332
rect 16948 17289 16957 17323
rect 16957 17289 16991 17323
rect 16991 17289 17000 17323
rect 16948 17280 17000 17289
rect 20168 17280 20220 17332
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 14096 17144 14148 17196
rect 14188 17144 14240 17196
rect 14740 17144 14792 17196
rect 13084 17076 13136 17128
rect 15108 17076 15160 17128
rect 18052 17255 18104 17264
rect 15844 17144 15896 17196
rect 16764 17144 16816 17196
rect 2596 17008 2648 17060
rect 13360 17008 13412 17060
rect 14188 17008 14240 17060
rect 16764 17008 16816 17060
rect 18052 17221 18061 17255
rect 18061 17221 18095 17255
rect 18095 17221 18104 17255
rect 18052 17212 18104 17221
rect 19248 17255 19300 17264
rect 19248 17221 19257 17255
rect 19257 17221 19291 17255
rect 19291 17221 19300 17255
rect 19248 17212 19300 17221
rect 20720 17212 20772 17264
rect 20904 17255 20956 17264
rect 20904 17221 20913 17255
rect 20913 17221 20947 17255
rect 20947 17221 20956 17255
rect 20904 17212 20956 17221
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 18144 17119 18196 17128
rect 18144 17085 18153 17119
rect 18153 17085 18187 17119
rect 18187 17085 18196 17119
rect 18144 17076 18196 17085
rect 24860 17280 24912 17332
rect 27620 17280 27672 17332
rect 29736 17280 29788 17332
rect 22100 17119 22152 17128
rect 22100 17085 22109 17119
rect 22109 17085 22143 17119
rect 22143 17085 22152 17119
rect 22100 17076 22152 17085
rect 5356 16940 5408 16992
rect 11336 16940 11388 16992
rect 13452 16940 13504 16992
rect 16212 16940 16264 16992
rect 16672 16940 16724 16992
rect 18880 17008 18932 17060
rect 22836 17076 22888 17128
rect 24952 17255 25004 17264
rect 23480 17076 23532 17128
rect 24308 17119 24360 17128
rect 24308 17085 24317 17119
rect 24317 17085 24351 17119
rect 24351 17085 24360 17119
rect 24308 17076 24360 17085
rect 23572 17008 23624 17060
rect 24584 17008 24636 17060
rect 24952 17221 24961 17255
rect 24961 17221 24995 17255
rect 24995 17221 25004 17255
rect 24952 17212 25004 17221
rect 25596 17212 25648 17264
rect 29184 17212 29236 17264
rect 25044 17076 25096 17128
rect 25688 17076 25740 17128
rect 26608 17144 26660 17196
rect 28816 17144 28868 17196
rect 29000 17144 29052 17196
rect 28632 17119 28684 17128
rect 25228 17008 25280 17060
rect 25596 17008 25648 17060
rect 20352 16940 20404 16992
rect 21088 16940 21140 16992
rect 23296 16940 23348 16992
rect 28632 17085 28641 17119
rect 28641 17085 28675 17119
rect 28675 17085 28684 17119
rect 28632 17076 28684 17085
rect 36268 17051 36320 17060
rect 36268 17017 36277 17051
rect 36277 17017 36311 17051
rect 36311 17017 36320 17051
rect 36268 17008 36320 17017
rect 26976 16940 27028 16992
rect 28724 16940 28776 16992
rect 30288 16983 30340 16992
rect 30288 16949 30297 16983
rect 30297 16949 30331 16983
rect 30331 16949 30340 16983
rect 30288 16940 30340 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 15200 16736 15252 16788
rect 15568 16736 15620 16788
rect 17776 16779 17828 16788
rect 17776 16745 17785 16779
rect 17785 16745 17819 16779
rect 17819 16745 17828 16779
rect 17776 16736 17828 16745
rect 15016 16711 15068 16720
rect 6736 16532 6788 16584
rect 15016 16677 15025 16711
rect 15025 16677 15059 16711
rect 15059 16677 15068 16711
rect 15016 16668 15068 16677
rect 12992 16600 13044 16652
rect 17684 16668 17736 16720
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 2136 16396 2188 16448
rect 2688 16396 2740 16448
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 12992 16396 13044 16448
rect 16672 16600 16724 16652
rect 16948 16600 17000 16652
rect 20628 16736 20680 16788
rect 20904 16736 20956 16788
rect 29828 16779 29880 16788
rect 29828 16745 29837 16779
rect 29837 16745 29871 16779
rect 29871 16745 29880 16779
rect 29828 16736 29880 16745
rect 18236 16668 18288 16720
rect 22928 16668 22980 16720
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 21548 16600 21600 16652
rect 24216 16668 24268 16720
rect 24584 16668 24636 16720
rect 26608 16668 26660 16720
rect 25780 16643 25832 16652
rect 25780 16609 25789 16643
rect 25789 16609 25823 16643
rect 25823 16609 25832 16643
rect 25780 16600 25832 16609
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 28264 16643 28316 16652
rect 28264 16609 28273 16643
rect 28273 16609 28307 16643
rect 28307 16609 28316 16643
rect 28264 16600 28316 16609
rect 30288 16643 30340 16652
rect 30288 16609 30297 16643
rect 30297 16609 30331 16643
rect 30331 16609 30340 16643
rect 30288 16600 30340 16609
rect 13912 16464 13964 16516
rect 15844 16464 15896 16516
rect 15016 16396 15068 16448
rect 18880 16464 18932 16516
rect 20168 16464 20220 16516
rect 20444 16507 20496 16516
rect 20444 16473 20453 16507
rect 20453 16473 20487 16507
rect 20487 16473 20496 16507
rect 20444 16464 20496 16473
rect 20536 16464 20588 16516
rect 22744 16507 22796 16516
rect 16948 16396 17000 16448
rect 20076 16396 20128 16448
rect 22744 16473 22753 16507
rect 22753 16473 22787 16507
rect 22787 16473 22796 16507
rect 22744 16464 22796 16473
rect 22836 16464 22888 16516
rect 23480 16507 23532 16516
rect 23480 16473 23489 16507
rect 23489 16473 23523 16507
rect 23523 16473 23532 16507
rect 23480 16464 23532 16473
rect 25044 16507 25096 16516
rect 25044 16473 25053 16507
rect 25053 16473 25087 16507
rect 25087 16473 25096 16507
rect 25044 16464 25096 16473
rect 25412 16464 25464 16516
rect 26976 16507 27028 16516
rect 25596 16396 25648 16448
rect 26976 16473 26985 16507
rect 26985 16473 27019 16507
rect 27019 16473 27028 16507
rect 26976 16464 27028 16473
rect 27068 16507 27120 16516
rect 27068 16473 27077 16507
rect 27077 16473 27111 16507
rect 27111 16473 27120 16507
rect 28172 16507 28224 16516
rect 27068 16464 27120 16473
rect 28172 16473 28181 16507
rect 28181 16473 28215 16507
rect 28215 16473 28224 16507
rect 28172 16464 28224 16473
rect 30288 16464 30340 16516
rect 28356 16396 28408 16448
rect 31116 16396 31168 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2320 16235 2372 16244
rect 2320 16201 2329 16235
rect 2329 16201 2363 16235
rect 2363 16201 2372 16235
rect 2320 16192 2372 16201
rect 9956 16192 10008 16244
rect 12348 16192 12400 16244
rect 12532 16192 12584 16244
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 2688 16056 2740 16108
rect 18144 16192 18196 16244
rect 19248 16192 19300 16244
rect 22376 16192 22428 16244
rect 18052 16124 18104 16176
rect 23572 16124 23624 16176
rect 27252 16192 27304 16244
rect 27896 16235 27948 16244
rect 27896 16201 27905 16235
rect 27905 16201 27939 16235
rect 27939 16201 27948 16235
rect 27896 16192 27948 16201
rect 28172 16192 28224 16244
rect 30288 16235 30340 16244
rect 30288 16201 30297 16235
rect 30297 16201 30331 16235
rect 30331 16201 30340 16235
rect 30288 16192 30340 16201
rect 24308 16124 24360 16176
rect 25412 16124 25464 16176
rect 26608 16124 26660 16176
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 2228 15988 2280 16040
rect 12992 15988 13044 16040
rect 2044 15920 2096 15972
rect 11612 15920 11664 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2688 15852 2740 15904
rect 13360 16056 13412 16108
rect 14372 16099 14424 16108
rect 14372 16065 14381 16099
rect 14381 16065 14415 16099
rect 14415 16065 14424 16099
rect 14372 16056 14424 16065
rect 18880 16056 18932 16108
rect 20352 16056 20404 16108
rect 21824 16056 21876 16108
rect 13452 15988 13504 16040
rect 15292 15988 15344 16040
rect 15108 15920 15160 15972
rect 15752 15963 15804 15972
rect 15752 15929 15761 15963
rect 15761 15929 15795 15963
rect 15795 15929 15804 15963
rect 15752 15920 15804 15929
rect 15844 15920 15896 15972
rect 18512 15963 18564 15972
rect 14648 15852 14700 15904
rect 15936 15852 15988 15904
rect 16212 15852 16264 15904
rect 18144 15852 18196 15904
rect 18512 15929 18521 15963
rect 18521 15929 18555 15963
rect 18555 15929 18564 15963
rect 18512 15920 18564 15929
rect 19340 16031 19392 16040
rect 19340 15997 19349 16031
rect 19349 15997 19383 16031
rect 19383 15997 19392 16031
rect 19340 15988 19392 15997
rect 19524 15988 19576 16040
rect 22652 15988 22704 16040
rect 23296 15988 23348 16040
rect 23480 15988 23532 16040
rect 24308 16031 24360 16040
rect 20352 15920 20404 15972
rect 22468 15920 22520 15972
rect 20812 15852 20864 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 24308 15997 24317 16031
rect 24317 15997 24351 16031
rect 24351 15997 24360 16031
rect 24308 15988 24360 15997
rect 25780 16031 25832 16040
rect 25780 15997 25789 16031
rect 25789 15997 25823 16031
rect 25823 15997 25832 16031
rect 25780 15988 25832 15997
rect 25872 15988 25924 16040
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 28632 16056 28684 16108
rect 31116 16099 31168 16108
rect 31116 16065 31125 16099
rect 31125 16065 31159 16099
rect 31159 16065 31168 16099
rect 31116 16056 31168 16065
rect 29920 15988 29972 16040
rect 27528 15920 27580 15972
rect 23112 15852 23164 15904
rect 24308 15852 24360 15904
rect 27068 15852 27120 15904
rect 27344 15852 27396 15904
rect 29828 15852 29880 15904
rect 36268 15895 36320 15904
rect 36268 15861 36277 15895
rect 36277 15861 36311 15895
rect 36311 15861 36320 15895
rect 36268 15852 36320 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1860 15648 1912 15700
rect 6736 15648 6788 15700
rect 15752 15648 15804 15700
rect 11152 15623 11204 15632
rect 11152 15589 11161 15623
rect 11161 15589 11195 15623
rect 11195 15589 11204 15623
rect 11152 15580 11204 15589
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 12348 15512 12400 15564
rect 13636 15555 13688 15564
rect 12716 15444 12768 15496
rect 13636 15521 13645 15555
rect 13645 15521 13679 15555
rect 13679 15521 13688 15555
rect 13636 15512 13688 15521
rect 13728 15444 13780 15496
rect 14832 15580 14884 15632
rect 16580 15580 16632 15632
rect 17316 15648 17368 15700
rect 23296 15648 23348 15700
rect 23572 15691 23624 15700
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 36084 15648 36136 15700
rect 19432 15580 19484 15632
rect 20812 15580 20864 15632
rect 18236 15512 18288 15564
rect 20536 15512 20588 15564
rect 20904 15512 20956 15564
rect 23756 15580 23808 15632
rect 25504 15580 25556 15632
rect 25872 15580 25924 15632
rect 25964 15580 26016 15632
rect 28080 15580 28132 15632
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 15844 15444 15896 15496
rect 19340 15444 19392 15496
rect 19524 15487 19576 15496
rect 19524 15453 19533 15487
rect 19533 15453 19567 15487
rect 19567 15453 19576 15487
rect 19524 15444 19576 15453
rect 20168 15444 20220 15496
rect 24400 15444 24452 15496
rect 27896 15512 27948 15564
rect 28632 15512 28684 15564
rect 29092 15555 29144 15564
rect 29092 15521 29101 15555
rect 29101 15521 29135 15555
rect 29135 15521 29144 15555
rect 29092 15512 29144 15521
rect 28264 15444 28316 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 14832 15376 14884 15428
rect 15108 15419 15160 15428
rect 15108 15385 15117 15419
rect 15117 15385 15151 15419
rect 15151 15385 15160 15419
rect 15108 15376 15160 15385
rect 15476 15376 15528 15428
rect 17224 15419 17276 15428
rect 17224 15385 17233 15419
rect 17233 15385 17267 15419
rect 17267 15385 17276 15419
rect 17224 15376 17276 15385
rect 17316 15419 17368 15428
rect 17316 15385 17325 15419
rect 17325 15385 17359 15419
rect 17359 15385 17368 15419
rect 17316 15376 17368 15385
rect 18144 15376 18196 15428
rect 19248 15376 19300 15428
rect 21272 15419 21324 15428
rect 21272 15385 21281 15419
rect 21281 15385 21315 15419
rect 21315 15385 21324 15419
rect 21272 15376 21324 15385
rect 11980 15308 12032 15360
rect 12624 15308 12676 15360
rect 13452 15308 13504 15360
rect 14096 15308 14148 15360
rect 16028 15308 16080 15360
rect 16120 15351 16172 15360
rect 16120 15317 16129 15351
rect 16129 15317 16163 15351
rect 16163 15317 16172 15351
rect 16120 15308 16172 15317
rect 17868 15308 17920 15360
rect 20168 15308 20220 15360
rect 20352 15308 20404 15360
rect 22376 15376 22428 15428
rect 22836 15376 22888 15428
rect 23480 15376 23532 15428
rect 25136 15419 25188 15428
rect 25136 15385 25145 15419
rect 25145 15385 25179 15419
rect 25179 15385 25188 15419
rect 25136 15376 25188 15385
rect 25412 15376 25464 15428
rect 27528 15419 27580 15428
rect 24676 15308 24728 15360
rect 24860 15308 24912 15360
rect 27528 15385 27537 15419
rect 27537 15385 27571 15419
rect 27571 15385 27580 15419
rect 27528 15376 27580 15385
rect 27804 15376 27856 15428
rect 28540 15419 28592 15428
rect 28540 15385 28549 15419
rect 28549 15385 28583 15419
rect 28583 15385 28592 15419
rect 28540 15376 28592 15385
rect 29276 15308 29328 15360
rect 29828 15351 29880 15360
rect 29828 15317 29837 15351
rect 29837 15317 29871 15351
rect 29871 15317 29880 15351
rect 29828 15308 29880 15317
rect 30472 15351 30524 15360
rect 30472 15317 30481 15351
rect 30481 15317 30515 15351
rect 30515 15317 30524 15351
rect 30472 15308 30524 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2596 15104 2648 15156
rect 17132 15104 17184 15156
rect 18052 15104 18104 15156
rect 20904 15147 20956 15156
rect 7564 15036 7616 15088
rect 9956 15079 10008 15088
rect 9956 15045 9965 15079
rect 9965 15045 9999 15079
rect 9999 15045 10008 15079
rect 9956 15036 10008 15045
rect 11152 15079 11204 15088
rect 11152 15045 11161 15079
rect 11161 15045 11195 15079
rect 11195 15045 11204 15079
rect 11152 15036 11204 15045
rect 13820 15036 13872 15088
rect 14372 15079 14424 15088
rect 14372 15045 14381 15079
rect 14381 15045 14415 15079
rect 14415 15045 14424 15079
rect 14372 15036 14424 15045
rect 18236 15036 18288 15088
rect 20076 15036 20128 15088
rect 20904 15113 20913 15147
rect 20913 15113 20947 15147
rect 20947 15113 20956 15147
rect 20904 15104 20956 15113
rect 22468 15104 22520 15156
rect 20536 15036 20588 15088
rect 22560 15079 22612 15088
rect 11796 14968 11848 15020
rect 15384 14968 15436 15020
rect 16396 14968 16448 15020
rect 17224 14968 17276 15020
rect 18696 14968 18748 15020
rect 8116 14900 8168 14952
rect 13544 14900 13596 14952
rect 14004 14900 14056 14952
rect 14096 14900 14148 14952
rect 14464 14900 14516 14952
rect 17868 14943 17920 14952
rect 8300 14832 8352 14884
rect 16764 14832 16816 14884
rect 13636 14764 13688 14816
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 22560 15045 22569 15079
rect 22569 15045 22603 15079
rect 22603 15045 22612 15079
rect 22560 15036 22612 15045
rect 22652 15036 22704 15088
rect 24308 15036 24360 15088
rect 24676 15104 24728 15156
rect 26884 15104 26936 15156
rect 28632 15147 28684 15156
rect 28632 15113 28641 15147
rect 28641 15113 28675 15147
rect 28675 15113 28684 15147
rect 28632 15104 28684 15113
rect 29092 15104 29144 15156
rect 35992 15147 36044 15156
rect 35992 15113 36001 15147
rect 36001 15113 36035 15147
rect 36035 15113 36044 15147
rect 35992 15104 36044 15113
rect 36176 15104 36228 15156
rect 25780 15079 25832 15088
rect 25780 15045 25789 15079
rect 25789 15045 25823 15079
rect 25823 15045 25832 15079
rect 25780 15036 25832 15045
rect 27620 15079 27672 15088
rect 27620 15045 27629 15079
rect 27629 15045 27663 15079
rect 27663 15045 27672 15079
rect 27620 15036 27672 15045
rect 29828 14968 29880 15020
rect 17132 14832 17184 14884
rect 17960 14764 18012 14816
rect 18328 14764 18380 14816
rect 19708 14875 19760 14884
rect 19708 14841 19717 14875
rect 19717 14841 19751 14875
rect 19751 14841 19760 14875
rect 19708 14832 19760 14841
rect 20536 14832 20588 14884
rect 20720 14764 20772 14816
rect 22376 14900 22428 14952
rect 23296 14943 23348 14952
rect 22192 14832 22244 14884
rect 23296 14909 23305 14943
rect 23305 14909 23339 14943
rect 23339 14909 23348 14943
rect 23296 14900 23348 14909
rect 23940 14943 23992 14952
rect 23940 14909 23949 14943
rect 23949 14909 23983 14943
rect 23983 14909 23992 14943
rect 23940 14900 23992 14909
rect 24584 14900 24636 14952
rect 25688 14943 25740 14952
rect 25688 14909 25697 14943
rect 25697 14909 25731 14943
rect 25731 14909 25740 14943
rect 25688 14900 25740 14909
rect 26332 14943 26384 14952
rect 26332 14909 26341 14943
rect 26341 14909 26375 14943
rect 26375 14909 26384 14943
rect 26332 14900 26384 14909
rect 27344 14900 27396 14952
rect 22928 14764 22980 14816
rect 23204 14832 23256 14884
rect 26424 14832 26476 14884
rect 27712 14900 27764 14952
rect 29000 14900 29052 14952
rect 29276 14943 29328 14952
rect 29276 14909 29285 14943
rect 29285 14909 29319 14943
rect 29319 14909 29328 14943
rect 29276 14900 29328 14909
rect 26792 14764 26844 14816
rect 28172 14764 28224 14816
rect 31116 14832 31168 14884
rect 30012 14764 30064 14816
rect 36176 14968 36228 15020
rect 31760 14764 31812 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 11244 14560 11296 14612
rect 14372 14560 14424 14612
rect 14740 14560 14792 14612
rect 20812 14560 20864 14612
rect 21272 14603 21324 14612
rect 21272 14569 21281 14603
rect 21281 14569 21315 14603
rect 21315 14569 21324 14603
rect 21272 14560 21324 14569
rect 21364 14560 21416 14612
rect 21548 14560 21600 14612
rect 23848 14560 23900 14612
rect 25780 14560 25832 14612
rect 26792 14560 26844 14612
rect 28264 14560 28316 14612
rect 11336 14424 11388 14476
rect 12900 14424 12952 14476
rect 14004 14492 14056 14544
rect 15476 14492 15528 14544
rect 26240 14535 26292 14544
rect 26240 14501 26249 14535
rect 26249 14501 26283 14535
rect 26283 14501 26292 14535
rect 26240 14492 26292 14501
rect 16764 14424 16816 14476
rect 17684 14424 17736 14476
rect 17776 14424 17828 14476
rect 18420 14424 18472 14476
rect 23204 14424 23256 14476
rect 23664 14424 23716 14476
rect 27068 14424 27120 14476
rect 30472 14424 30524 14476
rect 9956 14356 10008 14408
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 21180 14356 21232 14408
rect 12532 14288 12584 14340
rect 12716 14288 12768 14340
rect 15476 14331 15528 14340
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 11060 14220 11112 14272
rect 11336 14220 11388 14272
rect 12348 14220 12400 14272
rect 15476 14297 15485 14331
rect 15485 14297 15519 14331
rect 15519 14297 15528 14331
rect 15476 14288 15528 14297
rect 16672 14331 16724 14340
rect 16672 14297 16681 14331
rect 16681 14297 16715 14331
rect 16715 14297 16724 14331
rect 16672 14288 16724 14297
rect 16028 14220 16080 14272
rect 18328 14331 18380 14340
rect 18328 14297 18337 14331
rect 18337 14297 18371 14331
rect 18371 14297 18380 14331
rect 18328 14288 18380 14297
rect 20168 14288 20220 14340
rect 21088 14288 21140 14340
rect 22376 14331 22428 14340
rect 22376 14297 22385 14331
rect 22385 14297 22419 14331
rect 22419 14297 22428 14331
rect 22376 14288 22428 14297
rect 23848 14399 23900 14408
rect 23848 14365 23857 14399
rect 23857 14365 23891 14399
rect 23891 14365 23900 14399
rect 23848 14356 23900 14365
rect 28080 14399 28132 14408
rect 28080 14365 28089 14399
rect 28089 14365 28123 14399
rect 28123 14365 28132 14399
rect 28080 14356 28132 14365
rect 28356 14356 28408 14408
rect 29000 14356 29052 14408
rect 19340 14220 19392 14272
rect 20076 14220 20128 14272
rect 20720 14220 20772 14272
rect 21916 14220 21968 14272
rect 22008 14220 22060 14272
rect 22100 14220 22152 14272
rect 25320 14220 25372 14272
rect 25596 14331 25648 14340
rect 25596 14297 25605 14331
rect 25605 14297 25639 14331
rect 25639 14297 25648 14331
rect 25596 14288 25648 14297
rect 26976 14288 27028 14340
rect 27252 14288 27304 14340
rect 30104 14288 30156 14340
rect 30564 14356 30616 14408
rect 31760 14356 31812 14408
rect 30472 14263 30524 14272
rect 30472 14229 30481 14263
rect 30481 14229 30515 14263
rect 30515 14229 30524 14263
rect 30472 14220 30524 14229
rect 31116 14220 31168 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 13452 14016 13504 14068
rect 12624 13991 12676 14000
rect 12624 13957 12633 13991
rect 12633 13957 12667 13991
rect 12667 13957 12676 13991
rect 12624 13948 12676 13957
rect 14004 13948 14056 14000
rect 16396 14016 16448 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 9128 13923 9180 13932
rect 9128 13889 9137 13923
rect 9137 13889 9171 13923
rect 9171 13889 9180 13923
rect 9128 13880 9180 13889
rect 11612 13880 11664 13932
rect 11704 13880 11756 13932
rect 11520 13812 11572 13864
rect 12348 13812 12400 13864
rect 10968 13744 11020 13796
rect 11060 13744 11112 13796
rect 12624 13812 12676 13864
rect 14096 13880 14148 13932
rect 13636 13812 13688 13864
rect 15752 13991 15804 14000
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 20076 14016 20128 14068
rect 22008 14016 22060 14068
rect 22560 14016 22612 14068
rect 22652 14016 22704 14068
rect 23388 14016 23440 14068
rect 25228 14016 25280 14068
rect 15752 13948 15804 13957
rect 17408 13991 17460 14000
rect 17408 13957 17417 13991
rect 17417 13957 17451 13991
rect 17451 13957 17460 13991
rect 17408 13948 17460 13957
rect 17684 13948 17736 14000
rect 18236 13948 18288 14000
rect 18972 13991 19024 14000
rect 18972 13957 18981 13991
rect 18981 13957 19015 13991
rect 19015 13957 19024 13991
rect 18972 13948 19024 13957
rect 19064 13948 19116 14000
rect 20536 13991 20588 14000
rect 20536 13957 20545 13991
rect 20545 13957 20579 13991
rect 20579 13957 20588 13991
rect 20536 13948 20588 13957
rect 23572 13991 23624 14000
rect 23572 13957 23581 13991
rect 23581 13957 23615 13991
rect 23615 13957 23624 13991
rect 23572 13948 23624 13957
rect 26424 13948 26476 14000
rect 26884 13948 26936 14000
rect 30472 14016 30524 14068
rect 35992 14016 36044 14068
rect 27896 13948 27948 14000
rect 29092 13991 29144 14000
rect 29092 13957 29101 13991
rect 29101 13957 29135 13991
rect 29135 13957 29144 13991
rect 29092 13948 29144 13957
rect 21180 13880 21232 13932
rect 22100 13880 22152 13932
rect 22652 13923 22704 13932
rect 22652 13889 22661 13923
rect 22661 13889 22695 13923
rect 22695 13889 22704 13923
rect 22652 13880 22704 13889
rect 16764 13812 16816 13864
rect 18420 13812 18472 13864
rect 19524 13855 19576 13864
rect 19524 13821 19533 13855
rect 19533 13821 19567 13855
rect 19567 13821 19576 13855
rect 19524 13812 19576 13821
rect 14372 13744 14424 13796
rect 15016 13787 15068 13796
rect 15016 13753 15025 13787
rect 15025 13753 15059 13787
rect 15059 13753 15068 13787
rect 15016 13744 15068 13753
rect 17960 13744 18012 13796
rect 18236 13744 18288 13796
rect 19800 13744 19852 13796
rect 20076 13744 20128 13796
rect 20260 13812 20312 13864
rect 21732 13812 21784 13864
rect 23664 13812 23716 13864
rect 26976 13880 27028 13932
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 10692 13676 10744 13728
rect 12348 13676 12400 13728
rect 12992 13676 13044 13728
rect 17040 13676 17092 13728
rect 18420 13676 18472 13728
rect 25412 13812 25464 13864
rect 25964 13812 26016 13864
rect 24952 13744 25004 13796
rect 28080 13812 28132 13864
rect 28448 13855 28500 13864
rect 28448 13821 28457 13855
rect 28457 13821 28491 13855
rect 28491 13821 28500 13855
rect 28448 13812 28500 13821
rect 30104 13948 30156 14000
rect 29460 13812 29512 13864
rect 30380 13880 30432 13932
rect 36360 13923 36412 13932
rect 36360 13889 36369 13923
rect 36369 13889 36403 13923
rect 36403 13889 36412 13923
rect 36360 13880 36412 13889
rect 26240 13676 26292 13728
rect 26516 13676 26568 13728
rect 31576 13744 31628 13796
rect 29644 13719 29696 13728
rect 29644 13685 29653 13719
rect 29653 13685 29687 13719
rect 29687 13685 29696 13719
rect 29644 13676 29696 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10968 13472 11020 13524
rect 11704 13472 11756 13524
rect 12072 13472 12124 13524
rect 17408 13472 17460 13524
rect 18880 13515 18932 13524
rect 18880 13481 18889 13515
rect 18889 13481 18923 13515
rect 18923 13481 18932 13515
rect 18880 13472 18932 13481
rect 12716 13404 12768 13456
rect 13728 13404 13780 13456
rect 15844 13404 15896 13456
rect 20720 13404 20772 13456
rect 22008 13472 22060 13524
rect 22928 13472 22980 13524
rect 24860 13472 24912 13524
rect 25320 13515 25372 13524
rect 25320 13481 25329 13515
rect 25329 13481 25363 13515
rect 25363 13481 25372 13515
rect 25320 13472 25372 13481
rect 31576 13515 31628 13524
rect 1952 13268 2004 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9496 13268 9548 13320
rect 10784 13200 10836 13252
rect 11060 13243 11112 13252
rect 11060 13209 11069 13243
rect 11069 13209 11103 13243
rect 11103 13209 11112 13243
rect 11060 13200 11112 13209
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 11980 13200 12032 13252
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 13544 13336 13596 13388
rect 14004 13336 14056 13388
rect 15568 13336 15620 13388
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 16396 13336 16448 13345
rect 19524 13379 19576 13388
rect 19524 13345 19533 13379
rect 19533 13345 19567 13379
rect 19567 13345 19576 13379
rect 19524 13336 19576 13345
rect 19800 13379 19852 13388
rect 19800 13345 19809 13379
rect 19809 13345 19843 13379
rect 19843 13345 19852 13379
rect 19800 13336 19852 13345
rect 21088 13379 21140 13388
rect 21088 13345 21097 13379
rect 21097 13345 21131 13379
rect 21131 13345 21140 13379
rect 21088 13336 21140 13345
rect 21456 13336 21508 13388
rect 21732 13379 21784 13388
rect 21732 13345 21741 13379
rect 21741 13345 21775 13379
rect 21775 13345 21784 13379
rect 21732 13336 21784 13345
rect 22836 13404 22888 13456
rect 23572 13404 23624 13456
rect 25964 13404 26016 13456
rect 31576 13481 31585 13515
rect 31585 13481 31619 13515
rect 31619 13481 31628 13515
rect 31576 13472 31628 13481
rect 24860 13336 24912 13388
rect 27436 13336 27488 13388
rect 27528 13336 27580 13388
rect 28080 13336 28132 13388
rect 29184 13336 29236 13388
rect 12900 13268 12952 13320
rect 17592 13268 17644 13320
rect 19340 13268 19392 13320
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 24492 13268 24544 13320
rect 25688 13268 25740 13320
rect 15016 13243 15068 13252
rect 12624 13132 12676 13184
rect 15016 13209 15025 13243
rect 15025 13209 15059 13243
rect 15059 13209 15068 13243
rect 15016 13200 15068 13209
rect 15844 13243 15896 13252
rect 15844 13209 15853 13243
rect 15853 13209 15887 13243
rect 15887 13209 15896 13243
rect 15844 13200 15896 13209
rect 16672 13200 16724 13252
rect 16304 13132 16356 13184
rect 16488 13132 16540 13184
rect 17132 13200 17184 13252
rect 18144 13175 18196 13184
rect 18144 13141 18153 13175
rect 18153 13141 18187 13175
rect 18187 13141 18196 13175
rect 18144 13132 18196 13141
rect 19340 13132 19392 13184
rect 22284 13243 22336 13252
rect 22284 13209 22293 13243
rect 22293 13209 22327 13243
rect 22327 13209 22336 13243
rect 22284 13200 22336 13209
rect 22928 13243 22980 13252
rect 20996 13132 21048 13184
rect 21364 13132 21416 13184
rect 22928 13209 22937 13243
rect 22937 13209 22971 13243
rect 22971 13209 22980 13243
rect 26332 13268 26384 13320
rect 29000 13311 29052 13320
rect 29000 13277 29009 13311
rect 29009 13277 29043 13311
rect 29043 13277 29052 13311
rect 29000 13268 29052 13277
rect 30380 13404 30432 13456
rect 26240 13243 26292 13252
rect 22928 13200 22980 13209
rect 26240 13209 26249 13243
rect 26249 13209 26283 13243
rect 26283 13209 26292 13243
rect 26240 13200 26292 13209
rect 22468 13132 22520 13184
rect 27068 13132 27120 13184
rect 27712 13200 27764 13252
rect 27988 13243 28040 13252
rect 27988 13209 27997 13243
rect 27997 13209 28031 13243
rect 28031 13209 28040 13243
rect 27988 13200 28040 13209
rect 29644 13200 29696 13252
rect 36176 13336 36228 13388
rect 30288 13243 30340 13252
rect 30288 13209 30297 13243
rect 30297 13209 30331 13243
rect 30331 13209 30340 13243
rect 30288 13200 30340 13209
rect 31576 13132 31628 13184
rect 35900 13132 35952 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1860 12928 1912 12980
rect 4804 12928 4856 12980
rect 8392 12928 8444 12980
rect 11888 12928 11940 12980
rect 12072 12971 12124 12980
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 12348 12928 12400 12980
rect 8300 12792 8352 12844
rect 9496 12792 9548 12844
rect 9864 12792 9916 12844
rect 11428 12860 11480 12912
rect 11612 12792 11664 12844
rect 12072 12792 12124 12844
rect 12900 12860 12952 12912
rect 14832 12860 14884 12912
rect 15476 12860 15528 12912
rect 16856 12860 16908 12912
rect 17224 12860 17276 12912
rect 17500 12903 17552 12912
rect 17500 12869 17509 12903
rect 17509 12869 17543 12903
rect 17543 12869 17552 12903
rect 17500 12860 17552 12869
rect 18420 12903 18472 12912
rect 18420 12869 18429 12903
rect 18429 12869 18463 12903
rect 18463 12869 18472 12903
rect 18420 12860 18472 12869
rect 18972 12928 19024 12980
rect 21364 12971 21416 12980
rect 19524 12860 19576 12912
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 21732 12860 21784 12912
rect 27436 12928 27488 12980
rect 29736 12928 29788 12980
rect 30288 12928 30340 12980
rect 31576 12928 31628 12980
rect 35348 12928 35400 12980
rect 26056 12860 26108 12912
rect 18880 12792 18932 12844
rect 19432 12792 19484 12844
rect 21180 12792 21232 12844
rect 12348 12724 12400 12776
rect 12072 12588 12124 12640
rect 12440 12656 12492 12708
rect 12532 12656 12584 12708
rect 13360 12724 13412 12776
rect 13728 12656 13780 12708
rect 14280 12724 14332 12776
rect 15200 12724 15252 12776
rect 15844 12724 15896 12776
rect 17960 12724 18012 12776
rect 20720 12767 20772 12776
rect 19064 12656 19116 12708
rect 19800 12656 19852 12708
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 23480 12792 23532 12844
rect 23756 12792 23808 12844
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 24216 12792 24268 12844
rect 25412 12792 25464 12844
rect 21456 12724 21508 12776
rect 22376 12724 22428 12776
rect 23664 12724 23716 12776
rect 25964 12724 26016 12776
rect 13636 12588 13688 12640
rect 16120 12588 16172 12640
rect 18880 12588 18932 12640
rect 18972 12588 19024 12640
rect 19892 12588 19944 12640
rect 20444 12588 20496 12640
rect 23388 12656 23440 12708
rect 24584 12656 24636 12708
rect 26148 12656 26200 12708
rect 27068 12792 27120 12844
rect 27436 12792 27488 12844
rect 28724 12792 28776 12844
rect 29276 12792 29328 12844
rect 30472 12792 30524 12844
rect 26332 12724 26384 12776
rect 30748 12792 30800 12844
rect 31576 12724 31628 12776
rect 27068 12656 27120 12708
rect 30932 12656 30984 12708
rect 22836 12588 22888 12640
rect 25136 12588 25188 12640
rect 25320 12588 25372 12640
rect 27436 12588 27488 12640
rect 30656 12588 30708 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 8300 12248 8352 12300
rect 13084 12384 13136 12436
rect 13728 12384 13780 12436
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8668 12180 8720 12232
rect 9864 12180 9916 12232
rect 10692 12180 10744 12232
rect 11152 12180 11204 12232
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12256 12316 12308 12368
rect 15200 12316 15252 12368
rect 16304 12384 16356 12436
rect 16672 12316 16724 12368
rect 13176 12248 13228 12300
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 11336 12180 11388 12232
rect 11612 12180 11664 12232
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 12348 12180 12400 12232
rect 19800 12316 19852 12368
rect 19248 12248 19300 12300
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 20536 12384 20588 12436
rect 21824 12427 21876 12436
rect 21824 12393 21833 12427
rect 21833 12393 21867 12427
rect 21867 12393 21876 12427
rect 21824 12384 21876 12393
rect 23020 12384 23072 12436
rect 24768 12384 24820 12436
rect 29092 12384 29144 12436
rect 30932 12427 30984 12436
rect 30932 12393 30941 12427
rect 30941 12393 30975 12427
rect 30975 12393 30984 12427
rect 30932 12384 30984 12393
rect 31576 12427 31628 12436
rect 31576 12393 31585 12427
rect 31585 12393 31619 12427
rect 31619 12393 31628 12427
rect 31576 12384 31628 12393
rect 22836 12248 22888 12300
rect 26148 12248 26200 12300
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 16028 12180 16080 12232
rect 19156 12180 19208 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 20260 12180 20312 12232
rect 21272 12180 21324 12232
rect 23388 12180 23440 12232
rect 25412 12180 25464 12232
rect 25688 12180 25740 12232
rect 13544 12112 13596 12164
rect 14740 12155 14792 12164
rect 14740 12121 14749 12155
rect 14749 12121 14783 12155
rect 14783 12121 14792 12155
rect 14740 12112 14792 12121
rect 16580 12155 16632 12164
rect 16580 12121 16589 12155
rect 16589 12121 16623 12155
rect 16623 12121 16632 12155
rect 16580 12112 16632 12121
rect 16672 12155 16724 12164
rect 16672 12121 16681 12155
rect 16681 12121 16715 12155
rect 16715 12121 16724 12155
rect 16672 12112 16724 12121
rect 16856 12112 16908 12164
rect 22928 12155 22980 12164
rect 1860 12044 1912 12096
rect 8024 12044 8076 12096
rect 9588 12044 9640 12096
rect 11060 12044 11112 12096
rect 12440 12044 12492 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 15476 12044 15528 12096
rect 15936 12044 15988 12096
rect 16028 12044 16080 12096
rect 18788 12044 18840 12096
rect 19248 12044 19300 12096
rect 21272 12044 21324 12096
rect 22928 12121 22937 12155
rect 22937 12121 22971 12155
rect 22971 12121 22980 12155
rect 22928 12112 22980 12121
rect 24768 12112 24820 12164
rect 25596 12112 25648 12164
rect 25780 12155 25832 12164
rect 25780 12121 25789 12155
rect 25789 12121 25823 12155
rect 25823 12121 25832 12155
rect 25780 12112 25832 12121
rect 23664 12087 23716 12096
rect 23664 12053 23673 12087
rect 23673 12053 23707 12087
rect 23707 12053 23716 12087
rect 23664 12044 23716 12053
rect 23756 12044 23808 12096
rect 24032 12044 24084 12096
rect 26148 12112 26200 12164
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 26608 12180 26660 12189
rect 27068 12248 27120 12300
rect 30472 12316 30524 12368
rect 27344 12044 27396 12096
rect 29644 12112 29696 12164
rect 29828 12112 29880 12164
rect 30472 12155 30524 12164
rect 30472 12121 30481 12155
rect 30481 12121 30515 12155
rect 30515 12121 30524 12155
rect 30472 12112 30524 12121
rect 30656 12112 30708 12164
rect 31760 12112 31812 12164
rect 28448 12044 28500 12096
rect 32404 12044 32456 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 11152 11840 11204 11892
rect 12348 11840 12400 11892
rect 8760 11704 8812 11756
rect 11336 11772 11388 11824
rect 11520 11772 11572 11824
rect 12440 11772 12492 11824
rect 13636 11772 13688 11824
rect 14648 11815 14700 11824
rect 14648 11781 14657 11815
rect 14657 11781 14691 11815
rect 14691 11781 14700 11815
rect 15752 11840 15804 11892
rect 16764 11840 16816 11892
rect 20996 11840 21048 11892
rect 22284 11840 22336 11892
rect 22744 11840 22796 11892
rect 23388 11840 23440 11892
rect 25044 11840 25096 11892
rect 26424 11840 26476 11892
rect 27252 11883 27304 11892
rect 27252 11849 27261 11883
rect 27261 11849 27295 11883
rect 27295 11849 27304 11883
rect 27252 11840 27304 11849
rect 27804 11840 27856 11892
rect 28448 11840 28500 11892
rect 14648 11772 14700 11781
rect 10692 11704 10744 11756
rect 11060 11704 11112 11756
rect 14372 11704 14424 11756
rect 11796 11679 11848 11688
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 10876 11568 10928 11620
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12716 11636 12768 11688
rect 13268 11636 13320 11688
rect 15844 11704 15896 11756
rect 16212 11704 16264 11756
rect 17868 11747 17920 11756
rect 15292 11636 15344 11688
rect 16856 11636 16908 11688
rect 17868 11713 17877 11747
rect 17877 11713 17911 11747
rect 17911 11713 17920 11747
rect 17868 11704 17920 11713
rect 17960 11636 18012 11688
rect 13636 11568 13688 11620
rect 20444 11815 20496 11824
rect 20444 11781 20453 11815
rect 20453 11781 20487 11815
rect 20487 11781 20496 11815
rect 20444 11772 20496 11781
rect 20720 11772 20772 11824
rect 22560 11772 22612 11824
rect 23112 11772 23164 11824
rect 28816 11772 28868 11824
rect 21916 11704 21968 11756
rect 25228 11704 25280 11756
rect 25688 11704 25740 11756
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 18788 11679 18840 11688
rect 18788 11645 18797 11679
rect 18797 11645 18831 11679
rect 18831 11645 18840 11679
rect 22928 11679 22980 11688
rect 18788 11636 18840 11645
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 26240 11704 26292 11756
rect 27344 11747 27396 11756
rect 27344 11713 27353 11747
rect 27353 11713 27387 11747
rect 27387 11713 27396 11747
rect 27344 11704 27396 11713
rect 27528 11704 27580 11756
rect 28172 11704 28224 11756
rect 28448 11704 28500 11756
rect 29552 11704 29604 11756
rect 29736 11747 29788 11756
rect 29736 11713 29745 11747
rect 29745 11713 29779 11747
rect 29779 11713 29788 11747
rect 29736 11704 29788 11713
rect 36268 11747 36320 11756
rect 36268 11713 36277 11747
rect 36277 11713 36311 11747
rect 36311 11713 36320 11747
rect 36268 11704 36320 11713
rect 8208 11500 8260 11552
rect 10048 11500 10100 11552
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 15752 11500 15804 11552
rect 17868 11500 17920 11552
rect 20076 11500 20128 11552
rect 20812 11500 20864 11552
rect 28632 11568 28684 11620
rect 29000 11568 29052 11620
rect 29368 11568 29420 11620
rect 36084 11611 36136 11620
rect 36084 11577 36093 11611
rect 36093 11577 36127 11611
rect 36127 11577 36136 11611
rect 36084 11568 36136 11577
rect 25044 11500 25096 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 25596 11500 25648 11552
rect 30104 11500 30156 11552
rect 31668 11500 31720 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2504 11296 2556 11348
rect 9864 11296 9916 11348
rect 10416 11296 10468 11348
rect 13912 11296 13964 11348
rect 16580 11296 16632 11348
rect 10692 11228 10744 11280
rect 11060 11228 11112 11280
rect 11336 11271 11388 11280
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 12072 11228 12124 11280
rect 11888 11160 11940 11212
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 14188 11160 14240 11212
rect 15200 11160 15252 11212
rect 16580 11160 16632 11212
rect 17132 11160 17184 11212
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 12624 11092 12676 11144
rect 13636 11092 13688 11144
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 8024 11067 8076 11076
rect 8024 11033 8033 11067
rect 8033 11033 8067 11067
rect 8067 11033 8076 11067
rect 8024 11024 8076 11033
rect 9680 11024 9732 11076
rect 10876 11067 10928 11076
rect 10876 11033 10885 11067
rect 10885 11033 10919 11067
rect 10919 11033 10928 11067
rect 10876 11024 10928 11033
rect 12256 11024 12308 11076
rect 12992 11067 13044 11076
rect 12992 11033 13001 11067
rect 13001 11033 13035 11067
rect 13035 11033 13044 11067
rect 12992 11024 13044 11033
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 18052 11296 18104 11348
rect 20444 11296 20496 11348
rect 23204 11296 23256 11348
rect 25596 11296 25648 11348
rect 27896 11339 27948 11348
rect 27896 11305 27905 11339
rect 27905 11305 27939 11339
rect 27939 11305 27948 11339
rect 27896 11296 27948 11305
rect 29828 11339 29880 11348
rect 17500 11228 17552 11280
rect 17776 11228 17828 11280
rect 18236 11228 18288 11280
rect 21640 11228 21692 11280
rect 23296 11228 23348 11280
rect 27344 11228 27396 11280
rect 28724 11228 28776 11280
rect 29000 11228 29052 11280
rect 29828 11305 29837 11339
rect 29837 11305 29871 11339
rect 29871 11305 29880 11339
rect 29828 11296 29880 11305
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 19432 11160 19484 11212
rect 19984 11160 20036 11212
rect 20628 11160 20680 11212
rect 23664 11160 23716 11212
rect 11704 10956 11756 11008
rect 13360 10956 13412 11008
rect 14188 10956 14240 11008
rect 14464 10956 14516 11008
rect 15200 10999 15252 11008
rect 15200 10965 15209 10999
rect 15209 10965 15243 10999
rect 15243 10965 15252 10999
rect 15200 10956 15252 10965
rect 17316 11024 17368 11076
rect 17960 11024 18012 11076
rect 18788 11024 18840 11076
rect 22468 11092 22520 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 20720 11024 20772 11076
rect 18328 10956 18380 11008
rect 19524 10956 19576 11008
rect 20352 10956 20404 11008
rect 20996 10956 21048 11008
rect 21548 10956 21600 11008
rect 25780 11092 25832 11144
rect 26700 11135 26752 11144
rect 23572 11024 23624 11076
rect 24676 11067 24728 11076
rect 24676 11033 24685 11067
rect 24685 11033 24719 11067
rect 24719 11033 24728 11067
rect 24676 11024 24728 11033
rect 26700 11101 26709 11135
rect 26709 11101 26743 11135
rect 26743 11101 26752 11135
rect 26700 11092 26752 11101
rect 27344 11135 27396 11144
rect 27344 11101 27353 11135
rect 27353 11101 27387 11135
rect 27387 11101 27396 11135
rect 27344 11092 27396 11101
rect 28264 11092 28316 11144
rect 28540 11135 28592 11144
rect 28540 11101 28549 11135
rect 28549 11101 28583 11135
rect 28583 11101 28592 11135
rect 28540 11092 28592 11101
rect 28632 11135 28684 11144
rect 28632 11101 28641 11135
rect 28641 11101 28675 11135
rect 28675 11101 28684 11135
rect 29184 11135 29236 11144
rect 28632 11092 28684 11101
rect 29184 11101 29193 11135
rect 29193 11101 29227 11135
rect 29227 11101 29236 11135
rect 29184 11092 29236 11101
rect 29552 11092 29604 11144
rect 30104 11092 30156 11144
rect 24216 10956 24268 11008
rect 28448 11024 28500 11076
rect 24952 10956 25004 11008
rect 26148 10956 26200 11008
rect 27252 10999 27304 11008
rect 27252 10965 27261 10999
rect 27261 10965 27295 10999
rect 27295 10965 27304 10999
rect 27252 10956 27304 10965
rect 28632 10956 28684 11008
rect 31668 11092 31720 11144
rect 35532 11024 35584 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 7932 10752 7984 10804
rect 8760 10795 8812 10804
rect 8760 10761 8769 10795
rect 8769 10761 8803 10795
rect 8803 10761 8812 10795
rect 8760 10752 8812 10761
rect 10508 10727 10560 10736
rect 10508 10693 10517 10727
rect 10517 10693 10551 10727
rect 10551 10693 10560 10727
rect 10508 10684 10560 10693
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 10140 10616 10192 10668
rect 13084 10752 13136 10804
rect 16304 10752 16356 10804
rect 19340 10752 19392 10804
rect 20168 10752 20220 10804
rect 21272 10752 21324 10804
rect 21364 10752 21416 10804
rect 24952 10752 25004 10804
rect 25504 10752 25556 10804
rect 26056 10752 26108 10804
rect 27988 10752 28040 10804
rect 35532 10795 35584 10804
rect 35532 10761 35541 10795
rect 35541 10761 35575 10795
rect 35575 10761 35584 10795
rect 35532 10752 35584 10761
rect 11888 10684 11940 10736
rect 14832 10684 14884 10736
rect 17224 10684 17276 10736
rect 19248 10684 19300 10736
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 12900 10616 12952 10668
rect 11244 10548 11296 10600
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 9864 10480 9916 10532
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14464 10591 14516 10600
rect 14004 10548 14056 10557
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 12532 10412 12584 10464
rect 13636 10412 13688 10464
rect 16948 10616 17000 10668
rect 20260 10684 20312 10736
rect 22008 10684 22060 10736
rect 22744 10684 22796 10736
rect 16580 10548 16632 10600
rect 21272 10616 21324 10668
rect 23112 10684 23164 10736
rect 23664 10727 23716 10736
rect 23664 10693 23673 10727
rect 23673 10693 23707 10727
rect 23707 10693 23716 10727
rect 23664 10684 23716 10693
rect 25412 10684 25464 10736
rect 22928 10616 22980 10668
rect 26700 10684 26752 10736
rect 28080 10727 28132 10736
rect 28080 10693 28089 10727
rect 28089 10693 28123 10727
rect 28123 10693 28132 10727
rect 28080 10684 28132 10693
rect 26424 10616 26476 10668
rect 26884 10616 26936 10668
rect 29184 10616 29236 10668
rect 30012 10616 30064 10668
rect 30196 10616 30248 10668
rect 17132 10480 17184 10532
rect 19616 10480 19668 10532
rect 16028 10412 16080 10464
rect 16304 10412 16356 10464
rect 17960 10412 18012 10464
rect 20444 10548 20496 10600
rect 21088 10480 21140 10532
rect 27252 10548 27304 10600
rect 28724 10591 28776 10600
rect 28724 10557 28733 10591
rect 28733 10557 28767 10591
rect 28767 10557 28776 10591
rect 28724 10548 28776 10557
rect 35992 10616 36044 10668
rect 19984 10412 20036 10464
rect 20536 10412 20588 10464
rect 21364 10412 21416 10464
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 23388 10412 23440 10464
rect 26700 10480 26752 10532
rect 27160 10480 27212 10532
rect 24768 10412 24820 10464
rect 30380 10412 30432 10464
rect 36268 10455 36320 10464
rect 36268 10421 36277 10455
rect 36277 10421 36311 10455
rect 36311 10421 36320 10455
rect 36268 10412 36320 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 9404 10208 9456 10260
rect 11980 10208 12032 10260
rect 12992 10208 13044 10260
rect 15568 10208 15620 10260
rect 16028 10208 16080 10260
rect 18328 10208 18380 10260
rect 12900 10140 12952 10192
rect 13544 10140 13596 10192
rect 16764 10140 16816 10192
rect 17684 10140 17736 10192
rect 18052 10140 18104 10192
rect 18880 10208 18932 10260
rect 21456 10208 21508 10260
rect 21824 10208 21876 10260
rect 19340 10140 19392 10192
rect 20260 10140 20312 10192
rect 21916 10140 21968 10192
rect 9772 10072 9824 10124
rect 1768 9936 1820 9988
rect 2688 9936 2740 9988
rect 11888 10004 11940 10056
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 9772 9868 9824 9920
rect 12164 9868 12216 9920
rect 13452 10004 13504 10056
rect 14372 10004 14424 10056
rect 14648 10072 14700 10124
rect 16580 10072 16632 10124
rect 17592 10072 17644 10124
rect 21548 10072 21600 10124
rect 22744 10140 22796 10192
rect 25688 10208 25740 10260
rect 27620 10208 27672 10260
rect 23940 10140 23992 10192
rect 24860 10140 24912 10192
rect 28724 10140 28776 10192
rect 30380 10140 30432 10192
rect 30196 10072 30248 10124
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 18788 10004 18840 10056
rect 20168 10004 20220 10056
rect 20536 10047 20588 10056
rect 20536 10013 20545 10047
rect 20545 10013 20579 10047
rect 20579 10013 20588 10047
rect 20536 10004 20588 10013
rect 21916 10004 21968 10056
rect 24216 10004 24268 10056
rect 15384 9979 15436 9988
rect 15384 9945 15393 9979
rect 15393 9945 15427 9979
rect 15427 9945 15436 9979
rect 15384 9936 15436 9945
rect 16856 9936 16908 9988
rect 17316 9936 17368 9988
rect 18328 9936 18380 9988
rect 20720 9936 20772 9988
rect 20812 9979 20864 9988
rect 20812 9945 20821 9979
rect 20821 9945 20855 9979
rect 20855 9945 20864 9979
rect 20812 9936 20864 9945
rect 24676 10004 24728 10056
rect 26608 10047 26660 10056
rect 26608 10013 26617 10047
rect 26617 10013 26651 10047
rect 26651 10013 26660 10047
rect 27068 10047 27120 10056
rect 26608 10004 26660 10013
rect 27068 10013 27077 10047
rect 27077 10013 27111 10047
rect 27111 10013 27120 10047
rect 27068 10004 27120 10013
rect 27896 10047 27948 10056
rect 27896 10013 27905 10047
rect 27905 10013 27939 10047
rect 27939 10013 27948 10047
rect 27896 10004 27948 10013
rect 29184 10047 29236 10056
rect 29184 10013 29193 10047
rect 29193 10013 29227 10047
rect 29227 10013 29236 10047
rect 29184 10004 29236 10013
rect 30932 10004 30984 10056
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 17592 9868 17644 9920
rect 18052 9868 18104 9920
rect 18972 9868 19024 9920
rect 21088 9868 21140 9920
rect 21456 9868 21508 9920
rect 24860 9936 24912 9988
rect 23756 9911 23808 9920
rect 23756 9877 23765 9911
rect 23765 9877 23799 9911
rect 23799 9877 23808 9911
rect 23756 9868 23808 9877
rect 24032 9868 24084 9920
rect 24768 9868 24820 9920
rect 27620 9936 27672 9988
rect 28356 9936 28408 9988
rect 28724 9936 28776 9988
rect 29092 9936 29144 9988
rect 30196 9936 30248 9988
rect 27712 9868 27764 9920
rect 27988 9868 28040 9920
rect 30380 9979 30432 9988
rect 30380 9945 30389 9979
rect 30389 9945 30423 9979
rect 30423 9945 30432 9979
rect 30380 9936 30432 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 13084 9664 13136 9716
rect 15660 9664 15712 9716
rect 15844 9664 15896 9716
rect 32036 9664 32088 9716
rect 11428 9596 11480 9648
rect 11980 9596 12032 9648
rect 12532 9596 12584 9648
rect 14740 9596 14792 9648
rect 11704 9528 11756 9580
rect 10508 9503 10560 9512
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 12164 9460 12216 9512
rect 12256 9460 12308 9512
rect 14004 9528 14056 9580
rect 17040 9596 17092 9648
rect 18144 9596 18196 9648
rect 20352 9596 20404 9648
rect 25228 9596 25280 9648
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 25688 9596 25740 9648
rect 17316 9528 17368 9580
rect 20168 9528 20220 9580
rect 12716 9392 12768 9444
rect 15292 9460 15344 9512
rect 15660 9460 15712 9512
rect 16580 9460 16632 9512
rect 17776 9460 17828 9512
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 10968 9324 11020 9376
rect 14648 9324 14700 9376
rect 17040 9392 17092 9444
rect 19248 9392 19300 9444
rect 21456 9528 21508 9580
rect 15568 9324 15620 9376
rect 15844 9324 15896 9376
rect 17408 9324 17460 9376
rect 18052 9324 18104 9376
rect 18696 9324 18748 9376
rect 18880 9324 18932 9376
rect 19984 9324 20036 9376
rect 20352 9324 20404 9376
rect 20720 9324 20772 9376
rect 24492 9571 24544 9580
rect 24492 9537 24501 9571
rect 24501 9537 24535 9571
rect 24535 9537 24544 9571
rect 24492 9528 24544 9537
rect 25780 9528 25832 9580
rect 27344 9571 27396 9580
rect 27344 9537 27353 9571
rect 27353 9537 27387 9571
rect 27387 9537 27396 9571
rect 27344 9528 27396 9537
rect 27804 9528 27856 9580
rect 29552 9596 29604 9648
rect 29644 9596 29696 9648
rect 30564 9639 30616 9648
rect 30564 9605 30573 9639
rect 30573 9605 30607 9639
rect 30607 9605 30616 9639
rect 30564 9596 30616 9605
rect 30656 9639 30708 9648
rect 30656 9605 30665 9639
rect 30665 9605 30699 9639
rect 30699 9605 30708 9639
rect 30656 9596 30708 9605
rect 23848 9460 23900 9512
rect 26608 9460 26660 9512
rect 27896 9460 27948 9512
rect 29000 9528 29052 9580
rect 35992 9528 36044 9580
rect 26516 9392 26568 9444
rect 27160 9392 27212 9444
rect 24032 9324 24084 9376
rect 24216 9324 24268 9376
rect 26240 9324 26292 9376
rect 27804 9324 27856 9376
rect 28540 9367 28592 9376
rect 28540 9333 28549 9367
rect 28549 9333 28583 9367
rect 28583 9333 28592 9367
rect 28540 9324 28592 9333
rect 36084 9367 36136 9376
rect 36084 9333 36093 9367
rect 36093 9333 36127 9367
rect 36127 9333 36136 9367
rect 36084 9324 36136 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9772 9120 9824 9172
rect 10508 9163 10560 9172
rect 10508 9129 10517 9163
rect 10517 9129 10551 9163
rect 10551 9129 10560 9163
rect 10508 9120 10560 9129
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 12164 9120 12216 9172
rect 14280 9120 14332 9172
rect 15936 9120 15988 9172
rect 11060 9052 11112 9104
rect 13268 9095 13320 9104
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9680 8916 9732 8968
rect 13268 9061 13277 9095
rect 13277 9061 13311 9095
rect 13311 9061 13320 9095
rect 13268 9052 13320 9061
rect 18144 9120 18196 9172
rect 20076 9120 20128 9172
rect 22376 9120 22428 9172
rect 25228 9120 25280 9172
rect 17316 9052 17368 9104
rect 26056 9052 26108 9104
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 15476 8984 15528 9036
rect 18328 8984 18380 9036
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 11704 8916 11756 8968
rect 11796 8916 11848 8968
rect 13544 8916 13596 8968
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 15016 8916 15068 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 20444 8984 20496 9036
rect 20904 8984 20956 9036
rect 22928 8984 22980 9036
rect 24492 8984 24544 9036
rect 25504 8984 25556 9036
rect 26148 8984 26200 9036
rect 19984 8916 20036 8968
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 23112 8916 23164 8968
rect 26240 8916 26292 8968
rect 9956 8848 10008 8900
rect 12716 8848 12768 8900
rect 14924 8848 14976 8900
rect 18052 8891 18104 8900
rect 13360 8780 13412 8832
rect 15660 8780 15712 8832
rect 16028 8780 16080 8832
rect 16580 8780 16632 8832
rect 18052 8857 18061 8891
rect 18061 8857 18095 8891
rect 18095 8857 18104 8891
rect 18052 8848 18104 8857
rect 18144 8848 18196 8900
rect 20444 8848 20496 8900
rect 22100 8848 22152 8900
rect 24032 8891 24084 8900
rect 22376 8780 22428 8832
rect 24032 8857 24041 8891
rect 24041 8857 24075 8891
rect 24075 8857 24084 8891
rect 24032 8848 24084 8857
rect 26608 8984 26660 9036
rect 29552 9052 29604 9104
rect 27804 8984 27856 9036
rect 29184 8984 29236 9036
rect 30196 8984 30248 9036
rect 29828 8916 29880 8968
rect 30288 8916 30340 8968
rect 26608 8891 26660 8900
rect 26608 8857 26617 8891
rect 26617 8857 26651 8891
rect 26651 8857 26660 8891
rect 26608 8848 26660 8857
rect 26976 8848 27028 8900
rect 29184 8848 29236 8900
rect 31760 8848 31812 8900
rect 29276 8780 29328 8832
rect 29644 8780 29696 8832
rect 29920 8780 29972 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 13820 8576 13872 8628
rect 15384 8576 15436 8628
rect 15936 8576 15988 8628
rect 17776 8576 17828 8628
rect 20628 8576 20680 8628
rect 21548 8576 21600 8628
rect 21824 8576 21876 8628
rect 10140 8551 10192 8560
rect 10140 8517 10149 8551
rect 10149 8517 10183 8551
rect 10183 8517 10192 8551
rect 10140 8508 10192 8517
rect 10692 8551 10744 8560
rect 10692 8517 10701 8551
rect 10701 8517 10735 8551
rect 10735 8517 10744 8551
rect 10692 8508 10744 8517
rect 10784 8551 10836 8560
rect 10784 8517 10793 8551
rect 10793 8517 10827 8551
rect 10827 8517 10836 8551
rect 10784 8508 10836 8517
rect 13544 8508 13596 8560
rect 16028 8551 16080 8560
rect 16028 8517 16037 8551
rect 16037 8517 16071 8551
rect 16071 8517 16080 8551
rect 16856 8551 16908 8560
rect 16028 8508 16080 8517
rect 16856 8517 16865 8551
rect 16865 8517 16899 8551
rect 16899 8517 16908 8551
rect 16856 8508 16908 8517
rect 1584 8440 1636 8492
rect 13820 8440 13872 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 17592 8508 17644 8560
rect 17960 8508 18012 8560
rect 21180 8508 21232 8560
rect 22744 8508 22796 8560
rect 24216 8508 24268 8560
rect 24676 8576 24728 8628
rect 26608 8576 26660 8628
rect 27712 8576 27764 8628
rect 26516 8508 26568 8560
rect 30012 8508 30064 8560
rect 20260 8440 20312 8492
rect 21824 8440 21876 8492
rect 22928 8483 22980 8492
rect 22928 8449 22937 8483
rect 22937 8449 22971 8483
rect 22971 8449 22980 8483
rect 22928 8440 22980 8449
rect 27344 8440 27396 8492
rect 12716 8372 12768 8424
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 9680 8347 9732 8356
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 9680 8304 9732 8313
rect 11612 8304 11664 8356
rect 16580 8372 16632 8424
rect 17960 8372 18012 8424
rect 18144 8372 18196 8424
rect 19432 8372 19484 8424
rect 20536 8372 20588 8424
rect 22376 8372 22428 8424
rect 20260 8304 20312 8356
rect 15476 8236 15528 8288
rect 16028 8236 16080 8288
rect 21272 8304 21324 8356
rect 22284 8347 22336 8356
rect 22284 8313 22293 8347
rect 22293 8313 22327 8347
rect 22327 8313 22336 8347
rect 22284 8304 22336 8313
rect 22836 8304 22888 8356
rect 23664 8372 23716 8424
rect 26240 8415 26292 8424
rect 26240 8381 26249 8415
rect 26249 8381 26283 8415
rect 26283 8381 26292 8415
rect 26240 8372 26292 8381
rect 26424 8372 26476 8424
rect 27712 8440 27764 8492
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 28724 8440 28776 8492
rect 29828 8483 29880 8492
rect 29828 8449 29837 8483
rect 29837 8449 29871 8483
rect 29871 8449 29880 8483
rect 29828 8440 29880 8449
rect 28816 8372 28868 8424
rect 36084 8483 36136 8492
rect 36084 8449 36093 8483
rect 36093 8449 36127 8483
rect 36127 8449 36136 8483
rect 36084 8440 36136 8449
rect 24400 8304 24452 8356
rect 25688 8304 25740 8356
rect 24676 8236 24728 8288
rect 24860 8236 24912 8288
rect 26700 8236 26752 8288
rect 28448 8304 28500 8356
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 31300 8279 31352 8288
rect 31300 8245 31309 8279
rect 31309 8245 31343 8279
rect 31343 8245 31352 8279
rect 31300 8236 31352 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 10692 8032 10744 8084
rect 12624 8032 12676 8084
rect 13544 8032 13596 8084
rect 10784 7964 10836 8016
rect 10508 7896 10560 7948
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 11888 7828 11940 7880
rect 21180 8032 21232 8084
rect 23388 8032 23440 8084
rect 31300 8032 31352 8084
rect 19064 7964 19116 8016
rect 19432 7964 19484 8016
rect 14096 7828 14148 7880
rect 16580 7896 16632 7948
rect 17224 7896 17276 7948
rect 20628 7896 20680 7948
rect 22192 7939 22244 7948
rect 22192 7905 22201 7939
rect 22201 7905 22235 7939
rect 22235 7905 22244 7939
rect 24308 7964 24360 8016
rect 28080 7964 28132 8016
rect 22192 7896 22244 7905
rect 23664 7896 23716 7948
rect 24492 7896 24544 7948
rect 24860 7939 24912 7948
rect 24860 7905 24869 7939
rect 24869 7905 24903 7939
rect 24903 7905 24912 7939
rect 24860 7896 24912 7905
rect 25872 7896 25924 7948
rect 13728 7803 13780 7812
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 11060 7692 11112 7744
rect 13728 7769 13737 7803
rect 13737 7769 13771 7803
rect 13771 7769 13780 7803
rect 17592 7828 17644 7880
rect 18512 7828 18564 7880
rect 19248 7828 19300 7880
rect 26148 7828 26200 7880
rect 29000 7896 29052 7948
rect 30288 7896 30340 7948
rect 13728 7760 13780 7769
rect 17684 7760 17736 7812
rect 20904 7760 20956 7812
rect 21824 7760 21876 7812
rect 23756 7760 23808 7812
rect 27160 7760 27212 7812
rect 28356 7828 28408 7880
rect 28540 7828 28592 7880
rect 29828 7871 29880 7880
rect 29828 7837 29837 7871
rect 29837 7837 29871 7871
rect 29871 7837 29880 7871
rect 29828 7828 29880 7837
rect 32496 7828 32548 7880
rect 29368 7760 29420 7812
rect 16120 7692 16172 7744
rect 20168 7692 20220 7744
rect 22192 7692 22244 7744
rect 24952 7692 25004 7744
rect 26148 7692 26200 7744
rect 26516 7692 26568 7744
rect 26700 7692 26752 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 12072 7488 12124 7540
rect 12532 7488 12584 7540
rect 13636 7488 13688 7540
rect 2136 7420 2188 7472
rect 10140 7420 10192 7472
rect 10968 7463 11020 7472
rect 10968 7429 10977 7463
rect 10977 7429 11011 7463
rect 11011 7429 11020 7463
rect 10968 7420 11020 7429
rect 11336 7420 11388 7472
rect 13544 7420 13596 7472
rect 1584 7352 1636 7404
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 13728 7352 13780 7404
rect 20168 7488 20220 7540
rect 17224 7420 17276 7472
rect 17868 7420 17920 7472
rect 23388 7488 23440 7540
rect 29184 7531 29236 7540
rect 14188 7284 14240 7336
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 19064 7352 19116 7404
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 21824 7420 21876 7472
rect 22744 7420 22796 7472
rect 21272 7352 21324 7404
rect 20628 7284 20680 7293
rect 22744 7284 22796 7336
rect 24216 7420 24268 7472
rect 25596 7420 25648 7472
rect 29184 7497 29193 7531
rect 29193 7497 29227 7531
rect 29227 7497 29236 7531
rect 29184 7488 29236 7497
rect 25504 7352 25556 7404
rect 26700 7420 26752 7472
rect 35900 7420 35952 7472
rect 27896 7352 27948 7404
rect 28080 7352 28132 7404
rect 28540 7352 28592 7404
rect 29000 7352 29052 7404
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23940 7327 23992 7336
rect 23664 7284 23716 7293
rect 23940 7293 23949 7327
rect 23949 7293 23983 7327
rect 23983 7293 23992 7327
rect 23940 7284 23992 7293
rect 24032 7284 24084 7336
rect 29552 7352 29604 7404
rect 35808 7352 35860 7404
rect 2136 7148 2188 7200
rect 9680 7148 9732 7200
rect 12072 7148 12124 7200
rect 14280 7148 14332 7200
rect 18420 7148 18472 7200
rect 18880 7191 18932 7200
rect 18880 7157 18889 7191
rect 18889 7157 18923 7191
rect 18923 7157 18932 7191
rect 18880 7148 18932 7157
rect 20996 7216 21048 7268
rect 21456 7148 21508 7200
rect 22192 7216 22244 7268
rect 23572 7148 23624 7200
rect 27252 7191 27304 7200
rect 27252 7157 27261 7191
rect 27261 7157 27295 7191
rect 27295 7157 27304 7191
rect 27252 7148 27304 7157
rect 27528 7148 27580 7200
rect 28540 7191 28592 7200
rect 28540 7157 28549 7191
rect 28549 7157 28583 7191
rect 28583 7157 28592 7191
rect 28540 7148 28592 7157
rect 30380 7148 30432 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 10968 6944 11020 6996
rect 11520 6944 11572 6996
rect 12072 6944 12124 6996
rect 14280 6944 14332 6996
rect 14924 6944 14976 6996
rect 15200 6987 15252 6996
rect 15200 6953 15230 6987
rect 15230 6953 15252 6987
rect 15200 6944 15252 6953
rect 15568 6944 15620 6996
rect 20904 6944 20956 6996
rect 21824 6944 21876 6996
rect 27252 6944 27304 6996
rect 14188 6876 14240 6928
rect 9772 6808 9824 6860
rect 10140 6808 10192 6860
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 13544 6808 13596 6860
rect 14464 6808 14516 6860
rect 17868 6876 17920 6928
rect 19432 6876 19484 6928
rect 21916 6876 21968 6928
rect 28540 6876 28592 6928
rect 17500 6808 17552 6860
rect 18052 6808 18104 6860
rect 22100 6808 22152 6860
rect 24400 6808 24452 6860
rect 24492 6808 24544 6860
rect 24768 6808 24820 6860
rect 9404 6715 9456 6724
rect 9404 6681 9413 6715
rect 9413 6681 9447 6715
rect 9447 6681 9456 6715
rect 9404 6672 9456 6681
rect 19340 6740 19392 6792
rect 23204 6740 23256 6792
rect 16948 6715 17000 6724
rect 11244 6604 11296 6656
rect 12440 6604 12492 6656
rect 13912 6604 13964 6656
rect 14556 6604 14608 6656
rect 16948 6681 16957 6715
rect 16957 6681 16991 6715
rect 16991 6681 17000 6715
rect 16948 6672 17000 6681
rect 18236 6672 18288 6724
rect 18512 6672 18564 6724
rect 19064 6672 19116 6724
rect 21916 6672 21968 6724
rect 23940 6672 23992 6724
rect 17132 6604 17184 6656
rect 20812 6604 20864 6656
rect 21456 6604 21508 6656
rect 23020 6604 23072 6656
rect 23204 6647 23256 6656
rect 23204 6613 23213 6647
rect 23213 6613 23247 6647
rect 23247 6613 23256 6647
rect 23204 6604 23256 6613
rect 23664 6647 23716 6656
rect 23664 6613 23673 6647
rect 23673 6613 23707 6647
rect 23707 6613 23716 6647
rect 23664 6604 23716 6613
rect 26608 6740 26660 6792
rect 28080 6740 28132 6792
rect 28816 6783 28868 6792
rect 28816 6749 28825 6783
rect 28825 6749 28859 6783
rect 28859 6749 28868 6783
rect 28816 6740 28868 6749
rect 29000 6740 29052 6792
rect 30288 6740 30340 6792
rect 32496 6783 32548 6792
rect 32496 6749 32505 6783
rect 32505 6749 32539 6783
rect 32539 6749 32548 6783
rect 32496 6740 32548 6749
rect 26700 6672 26752 6724
rect 31852 6672 31904 6724
rect 27252 6604 27304 6656
rect 28080 6647 28132 6656
rect 28080 6613 28089 6647
rect 28089 6613 28123 6647
rect 28123 6613 28132 6647
rect 28080 6604 28132 6613
rect 28724 6647 28776 6656
rect 28724 6613 28733 6647
rect 28733 6613 28767 6647
rect 28767 6613 28776 6647
rect 28724 6604 28776 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 8208 6400 8260 6452
rect 9772 6400 9824 6452
rect 11980 6400 12032 6452
rect 11428 6332 11480 6384
rect 14464 6400 14516 6452
rect 13912 6332 13964 6384
rect 17132 6400 17184 6452
rect 20260 6400 20312 6452
rect 22100 6400 22152 6452
rect 20628 6332 20680 6384
rect 23664 6400 23716 6452
rect 23848 6400 23900 6452
rect 26240 6400 26292 6452
rect 22284 6375 22336 6384
rect 13728 6264 13780 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 21272 6264 21324 6316
rect 22284 6341 22293 6375
rect 22293 6341 22327 6375
rect 22327 6341 22336 6375
rect 22284 6332 22336 6341
rect 23296 6332 23348 6384
rect 24952 6332 25004 6384
rect 27804 6375 27856 6384
rect 27804 6341 27813 6375
rect 27813 6341 27847 6375
rect 27847 6341 27856 6375
rect 27804 6332 27856 6341
rect 27896 6307 27948 6316
rect 9680 6196 9732 6248
rect 13820 6196 13872 6248
rect 14372 6196 14424 6248
rect 14648 6196 14700 6248
rect 16856 6196 16908 6248
rect 17592 6196 17644 6248
rect 19248 6196 19300 6248
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 11520 6060 11572 6112
rect 11704 6060 11756 6112
rect 12348 6060 12400 6112
rect 13912 6128 13964 6180
rect 15016 6128 15068 6180
rect 14004 6060 14056 6112
rect 18512 6128 18564 6180
rect 18880 6128 18932 6180
rect 22284 6196 22336 6248
rect 23020 6196 23072 6248
rect 24584 6239 24636 6248
rect 24584 6205 24593 6239
rect 24593 6205 24627 6239
rect 24627 6205 24636 6239
rect 24584 6196 24636 6205
rect 27896 6273 27905 6307
rect 27905 6273 27939 6307
rect 27939 6273 27948 6307
rect 27896 6264 27948 6273
rect 29552 6264 29604 6316
rect 30288 6264 30340 6316
rect 27528 6196 27580 6248
rect 16948 6060 17000 6112
rect 22928 6060 22980 6112
rect 23480 6060 23532 6112
rect 26976 6060 27028 6112
rect 27252 6103 27304 6112
rect 27252 6069 27261 6103
rect 27261 6069 27295 6103
rect 27295 6069 27304 6103
rect 27252 6060 27304 6069
rect 29092 6060 29144 6112
rect 29644 6103 29696 6112
rect 29644 6069 29653 6103
rect 29653 6069 29687 6103
rect 29687 6069 29696 6103
rect 29644 6060 29696 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 9404 5856 9456 5908
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 12256 5856 12308 5908
rect 13912 5856 13964 5908
rect 14004 5856 14056 5908
rect 22192 5856 22244 5908
rect 24860 5856 24912 5908
rect 25964 5856 26016 5908
rect 26240 5856 26292 5908
rect 31760 5899 31812 5908
rect 31760 5865 31769 5899
rect 31769 5865 31803 5899
rect 31803 5865 31812 5899
rect 31760 5856 31812 5865
rect 9128 5788 9180 5840
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 14096 5788 14148 5840
rect 14924 5831 14976 5840
rect 14924 5797 14933 5831
rect 14933 5797 14967 5831
rect 14967 5797 14976 5831
rect 14924 5788 14976 5797
rect 18328 5788 18380 5840
rect 18512 5788 18564 5840
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 17592 5763 17644 5772
rect 17592 5729 17601 5763
rect 17601 5729 17635 5763
rect 17635 5729 17644 5763
rect 17592 5720 17644 5729
rect 17868 5720 17920 5772
rect 21548 5788 21600 5840
rect 20352 5720 20404 5772
rect 23848 5720 23900 5772
rect 24584 5720 24636 5772
rect 11152 5652 11204 5704
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 13544 5652 13596 5704
rect 15844 5652 15896 5704
rect 11796 5584 11848 5636
rect 11980 5584 12032 5636
rect 13636 5584 13688 5636
rect 16304 5584 16356 5636
rect 18052 5584 18104 5636
rect 13728 5559 13780 5568
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 14556 5516 14608 5568
rect 21456 5652 21508 5704
rect 23388 5652 23440 5704
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 30288 5652 30340 5704
rect 31208 5652 31260 5704
rect 21088 5584 21140 5636
rect 19248 5516 19300 5568
rect 21272 5516 21324 5568
rect 21732 5516 21784 5568
rect 24768 5584 24820 5636
rect 25504 5584 25556 5636
rect 25964 5584 26016 5636
rect 23572 5559 23624 5568
rect 23572 5525 23581 5559
rect 23581 5525 23615 5559
rect 23615 5525 23624 5559
rect 23572 5516 23624 5525
rect 27344 5559 27396 5568
rect 27344 5525 27353 5559
rect 27353 5525 27387 5559
rect 27387 5525 27396 5559
rect 27344 5516 27396 5525
rect 29184 5516 29236 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 11060 5312 11112 5364
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 12072 5312 12124 5364
rect 9772 5287 9824 5296
rect 9772 5253 9781 5287
rect 9781 5253 9815 5287
rect 9815 5253 9824 5287
rect 9772 5244 9824 5253
rect 15752 5312 15804 5364
rect 16212 5355 16264 5364
rect 16212 5321 16221 5355
rect 16221 5321 16255 5355
rect 16255 5321 16264 5355
rect 16212 5312 16264 5321
rect 17960 5312 18012 5364
rect 14372 5244 14424 5296
rect 14464 5244 14516 5296
rect 14832 5244 14884 5296
rect 16488 5244 16540 5296
rect 18512 5244 18564 5296
rect 21732 5244 21784 5296
rect 1584 5176 1636 5228
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 16120 5176 16172 5228
rect 17592 5176 17644 5228
rect 21916 5176 21968 5228
rect 23204 5244 23256 5296
rect 25872 5244 25924 5296
rect 26424 5312 26476 5364
rect 27068 5312 27120 5364
rect 26884 5244 26936 5296
rect 24584 5219 24636 5228
rect 24584 5185 24593 5219
rect 24593 5185 24627 5219
rect 24627 5185 24636 5219
rect 24584 5176 24636 5185
rect 26240 5176 26292 5228
rect 30104 5244 30156 5296
rect 27896 5176 27948 5228
rect 30012 5176 30064 5228
rect 36176 5176 36228 5228
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 9864 5108 9916 5160
rect 13544 4972 13596 5024
rect 15844 5040 15896 5092
rect 16396 5040 16448 5092
rect 16672 5040 16724 5092
rect 21640 5108 21692 5160
rect 15752 4972 15804 5024
rect 21456 4972 21508 5024
rect 23112 4972 23164 5024
rect 23388 4972 23440 5024
rect 26792 5108 26844 5160
rect 27252 5108 27304 5160
rect 28816 5108 28868 5160
rect 36360 5151 36412 5160
rect 36360 5117 36369 5151
rect 36369 5117 36403 5151
rect 36403 5117 36412 5151
rect 36360 5108 36412 5117
rect 24308 4972 24360 5024
rect 28724 5040 28776 5092
rect 25964 4972 26016 5024
rect 29460 5040 29512 5092
rect 29000 5015 29052 5024
rect 29000 4981 29009 5015
rect 29009 4981 29043 5015
rect 29043 4981 29052 5015
rect 29000 4972 29052 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 9128 4811 9180 4820
rect 9128 4777 9137 4811
rect 9137 4777 9171 4811
rect 9171 4777 9180 4811
rect 9128 4768 9180 4777
rect 9772 4811 9824 4820
rect 9772 4777 9781 4811
rect 9781 4777 9815 4811
rect 9815 4777 9824 4811
rect 9772 4768 9824 4777
rect 11336 4768 11388 4820
rect 12164 4768 12216 4820
rect 14004 4768 14056 4820
rect 11704 4632 11756 4684
rect 17408 4768 17460 4820
rect 18788 4811 18840 4820
rect 18788 4777 18797 4811
rect 18797 4777 18831 4811
rect 18831 4777 18840 4811
rect 18788 4768 18840 4777
rect 15476 4700 15528 4752
rect 18052 4700 18104 4752
rect 9128 4564 9180 4616
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 16396 4632 16448 4684
rect 17868 4632 17920 4684
rect 15568 4496 15620 4548
rect 17040 4564 17092 4616
rect 15936 4539 15988 4548
rect 15936 4505 15945 4539
rect 15945 4505 15979 4539
rect 15979 4505 15988 4539
rect 15936 4496 15988 4505
rect 18236 4700 18288 4752
rect 20720 4768 20772 4820
rect 18788 4632 18840 4684
rect 19616 4632 19668 4684
rect 20076 4632 20128 4684
rect 20720 4632 20772 4684
rect 19064 4564 19116 4616
rect 24308 4768 24360 4820
rect 14924 4428 14976 4480
rect 15844 4428 15896 4480
rect 18696 4428 18748 4480
rect 24308 4632 24360 4684
rect 22100 4564 22152 4616
rect 29000 4768 29052 4820
rect 30564 4768 30616 4820
rect 36360 4811 36412 4820
rect 36360 4777 36369 4811
rect 36369 4777 36403 4811
rect 36403 4777 36412 4811
rect 36360 4768 36412 4777
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 24860 4675 24912 4684
rect 24860 4641 24869 4675
rect 24869 4641 24903 4675
rect 24903 4641 24912 4675
rect 24860 4632 24912 4641
rect 26608 4632 26660 4684
rect 26700 4632 26752 4684
rect 26976 4632 27028 4684
rect 26516 4564 26568 4616
rect 27620 4564 27672 4616
rect 27804 4564 27856 4616
rect 28632 4564 28684 4616
rect 21548 4428 21600 4480
rect 22836 4496 22888 4548
rect 26240 4496 26292 4548
rect 27344 4496 27396 4548
rect 24124 4428 24176 4480
rect 27620 4428 27672 4480
rect 28724 4428 28776 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 13268 4224 13320 4276
rect 10784 4088 10836 4140
rect 11336 4088 11388 4140
rect 12237 4199 12289 4208
rect 12237 4165 12252 4199
rect 12252 4165 12286 4199
rect 12286 4165 12289 4199
rect 12237 4156 12289 4165
rect 13544 4156 13596 4208
rect 15844 4224 15896 4276
rect 15568 4156 15620 4208
rect 16212 4224 16264 4276
rect 16856 4224 16908 4276
rect 18512 4156 18564 4208
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16856 4131 16908 4140
rect 16304 4088 16356 4097
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 18696 4224 18748 4276
rect 21916 4224 21968 4276
rect 22468 4224 22520 4276
rect 23388 4224 23440 4276
rect 26516 4267 26568 4276
rect 19432 4156 19484 4208
rect 21824 4156 21876 4208
rect 23480 4156 23532 4208
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 20996 4088 21048 4140
rect 21548 4088 21600 4140
rect 26516 4233 26525 4267
rect 26525 4233 26559 4267
rect 26559 4233 26568 4267
rect 26516 4224 26568 4233
rect 26608 4224 26660 4276
rect 31392 4224 31444 4276
rect 26056 4156 26108 4208
rect 29644 4156 29696 4208
rect 26332 4088 26384 4140
rect 29000 4088 29052 4140
rect 30012 4131 30064 4140
rect 30012 4097 30021 4131
rect 30021 4097 30055 4131
rect 30055 4097 30064 4131
rect 31760 4156 31812 4208
rect 30748 4131 30800 4140
rect 30012 4088 30064 4097
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 30748 4088 30800 4097
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 11244 3952 11296 4004
rect 13452 4020 13504 4072
rect 13820 4020 13872 4072
rect 17132 4063 17184 4072
rect 14464 3952 14516 4004
rect 13636 3884 13688 3936
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14556 3884 14608 3936
rect 16764 3884 16816 3936
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 20904 4020 20956 4072
rect 20720 3952 20772 4004
rect 21824 3952 21876 4004
rect 23848 4020 23900 4072
rect 25044 4020 25096 4072
rect 26056 4020 26108 4072
rect 26884 4020 26936 4072
rect 23388 3884 23440 3936
rect 25872 3952 25924 4004
rect 28540 4020 28592 4072
rect 28632 4063 28684 4072
rect 28632 4029 28641 4063
rect 28641 4029 28675 4063
rect 28675 4029 28684 4063
rect 28632 4020 28684 4029
rect 30472 3952 30524 4004
rect 35900 3995 35952 4004
rect 35900 3961 35909 3995
rect 35909 3961 35943 3995
rect 35943 3961 35952 3995
rect 35900 3952 35952 3961
rect 26424 3884 26476 3936
rect 26792 3884 26844 3936
rect 29000 3884 29052 3936
rect 29552 3884 29604 3936
rect 31300 3884 31352 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 11612 3680 11664 3732
rect 12440 3680 12492 3732
rect 13728 3680 13780 3732
rect 13636 3612 13688 3664
rect 11888 3544 11940 3596
rect 14556 3544 14608 3596
rect 7840 3476 7892 3528
rect 5540 3408 5592 3460
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11980 3519 12032 3528
rect 11520 3476 11572 3485
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 14188 3476 14240 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 15108 3544 15160 3596
rect 16856 3544 16908 3596
rect 18328 3544 18380 3596
rect 15844 3476 15896 3528
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 2412 3383 2464 3392
rect 2412 3349 2421 3383
rect 2421 3349 2455 3383
rect 2455 3349 2464 3383
rect 2412 3340 2464 3349
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 10784 3408 10836 3460
rect 11152 3408 11204 3460
rect 11796 3340 11848 3392
rect 15016 3408 15068 3460
rect 15292 3408 15344 3460
rect 19064 3680 19116 3732
rect 22192 3680 22244 3732
rect 22560 3680 22612 3732
rect 23572 3680 23624 3732
rect 24584 3680 24636 3732
rect 26332 3680 26384 3732
rect 26424 3680 26476 3732
rect 27620 3680 27672 3732
rect 27712 3680 27764 3732
rect 28540 3723 28592 3732
rect 18696 3612 18748 3664
rect 19800 3612 19852 3664
rect 19984 3655 20036 3664
rect 19984 3621 19993 3655
rect 19993 3621 20027 3655
rect 20027 3621 20036 3655
rect 19984 3612 20036 3621
rect 28540 3689 28549 3723
rect 28549 3689 28583 3723
rect 28583 3689 28592 3723
rect 28540 3680 28592 3689
rect 31208 3680 31260 3732
rect 31392 3723 31444 3732
rect 31392 3689 31401 3723
rect 31401 3689 31435 3723
rect 31435 3689 31444 3723
rect 31392 3680 31444 3689
rect 32036 3723 32088 3732
rect 32036 3689 32045 3723
rect 32045 3689 32079 3723
rect 32079 3689 32088 3723
rect 32036 3680 32088 3689
rect 29736 3612 29788 3664
rect 35348 3612 35400 3664
rect 21088 3544 21140 3596
rect 22100 3544 22152 3596
rect 22192 3587 22244 3596
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 24584 3587 24636 3596
rect 22192 3544 22244 3553
rect 24584 3553 24593 3587
rect 24593 3553 24627 3587
rect 24627 3553 24636 3587
rect 24584 3544 24636 3553
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 25228 3544 25280 3596
rect 25872 3544 25924 3596
rect 19340 3476 19392 3528
rect 21824 3476 21876 3528
rect 21456 3451 21508 3460
rect 14832 3340 14884 3392
rect 18604 3340 18656 3392
rect 19340 3340 19392 3392
rect 21456 3417 21465 3451
rect 21465 3417 21499 3451
rect 21499 3417 21508 3451
rect 21456 3408 21508 3417
rect 21732 3340 21784 3392
rect 26332 3476 26384 3528
rect 26792 3519 26844 3528
rect 26792 3485 26801 3519
rect 26801 3485 26835 3519
rect 26835 3485 26844 3519
rect 26792 3476 26844 3485
rect 28448 3476 28500 3528
rect 29736 3476 29788 3528
rect 29920 3476 29972 3528
rect 22468 3451 22520 3460
rect 22468 3417 22477 3451
rect 22477 3417 22511 3451
rect 22511 3417 22520 3451
rect 22468 3408 22520 3417
rect 24400 3408 24452 3460
rect 24308 3340 24360 3392
rect 25136 3408 25188 3460
rect 27068 3451 27120 3460
rect 27068 3417 27077 3451
rect 27077 3417 27111 3451
rect 27111 3417 27120 3451
rect 27068 3408 27120 3417
rect 27344 3408 27396 3460
rect 28356 3408 28408 3460
rect 28816 3408 28868 3460
rect 24768 3340 24820 3392
rect 26240 3340 26292 3392
rect 26884 3340 26936 3392
rect 29000 3383 29052 3392
rect 29000 3349 29009 3383
rect 29009 3349 29043 3383
rect 29043 3349 29052 3383
rect 29000 3340 29052 3349
rect 29736 3340 29788 3392
rect 31024 3340 31076 3392
rect 31760 3476 31812 3528
rect 32036 3476 32088 3528
rect 32496 3544 32548 3596
rect 32220 3476 32272 3528
rect 32956 3476 33008 3528
rect 35900 3476 35952 3528
rect 31576 3408 31628 3460
rect 36268 3383 36320 3392
rect 36268 3349 36277 3383
rect 36277 3349 36311 3383
rect 36311 3349 36320 3383
rect 36268 3340 36320 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 9680 3136 9732 3188
rect 8576 3068 8628 3120
rect 11060 3068 11112 3120
rect 11520 3068 11572 3120
rect 12992 3068 13044 3120
rect 13452 3111 13504 3120
rect 13452 3077 13461 3111
rect 13461 3077 13495 3111
rect 13495 3077 13504 3111
rect 13452 3068 13504 3077
rect 2412 3000 2464 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 9588 3000 9640 3052
rect 15844 3136 15896 3188
rect 16304 3136 16356 3188
rect 15016 3068 15068 3120
rect 16396 3068 16448 3120
rect 9496 2932 9548 2984
rect 11888 2932 11940 2984
rect 17132 3136 17184 3188
rect 21364 3136 21416 3188
rect 21456 3136 21508 3188
rect 17868 3068 17920 3120
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 19064 3068 19116 3120
rect 20812 3068 20864 3120
rect 22192 3136 22244 3188
rect 26608 3136 26660 3188
rect 26792 3136 26844 3188
rect 28356 3136 28408 3188
rect 32404 3179 32456 3188
rect 22468 3068 22520 3120
rect 24860 3068 24912 3120
rect 26148 3068 26200 3120
rect 27620 3068 27672 3120
rect 28816 3068 28868 3120
rect 29000 3068 29052 3120
rect 30840 3068 30892 3120
rect 32404 3145 32413 3179
rect 32413 3145 32447 3179
rect 32447 3145 32456 3179
rect 32404 3136 32456 3145
rect 18696 2932 18748 2984
rect 19432 2932 19484 2984
rect 24492 3043 24544 3052
rect 24492 3009 24501 3043
rect 24501 3009 24535 3043
rect 24535 3009 24544 3043
rect 24492 3000 24544 3009
rect 29552 3000 29604 3052
rect 29644 3000 29696 3052
rect 20 2796 72 2848
rect 1860 2796 1912 2848
rect 2780 2796 2832 2848
rect 12440 2796 12492 2848
rect 12716 2796 12768 2848
rect 16304 2796 16356 2848
rect 18052 2796 18104 2848
rect 18604 2796 18656 2848
rect 22652 2864 22704 2916
rect 20168 2796 20220 2848
rect 21456 2796 21508 2848
rect 24308 2932 24360 2984
rect 24400 2932 24452 2984
rect 24860 2932 24912 2984
rect 26608 2932 26660 2984
rect 32956 3043 33008 3052
rect 32956 3009 32965 3043
rect 32965 3009 32999 3043
rect 32999 3009 33008 3043
rect 32956 3000 33008 3009
rect 35992 3000 36044 3052
rect 36268 3043 36320 3052
rect 36268 3009 36277 3043
rect 36277 3009 36311 3043
rect 36311 3009 36320 3043
rect 36268 3000 36320 3009
rect 31576 2864 31628 2916
rect 32864 2864 32916 2916
rect 24032 2796 24084 2848
rect 27712 2796 27764 2848
rect 30564 2796 30616 2848
rect 31024 2839 31076 2848
rect 31024 2805 31033 2839
rect 31033 2805 31067 2839
rect 31067 2805 31076 2839
rect 31024 2796 31076 2805
rect 31116 2796 31168 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 15844 2592 15896 2644
rect 5540 2524 5592 2576
rect 16580 2524 16632 2576
rect 11520 2456 11572 2508
rect 17868 2456 17920 2508
rect 21916 2456 21968 2508
rect 22100 2499 22152 2508
rect 22100 2465 22109 2499
rect 22109 2465 22143 2499
rect 22143 2465 22152 2499
rect 22100 2456 22152 2465
rect 25964 2456 26016 2508
rect 26332 2499 26384 2508
rect 26332 2465 26341 2499
rect 26341 2465 26375 2499
rect 26375 2465 26384 2499
rect 26332 2456 26384 2465
rect 28632 2592 28684 2644
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 29184 2524 29236 2576
rect 28632 2456 28684 2508
rect 28908 2456 28960 2508
rect 30564 2499 30616 2508
rect 30564 2465 30573 2499
rect 30573 2465 30607 2499
rect 30607 2465 30616 2499
rect 30564 2456 30616 2465
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 2780 2388 2832 2440
rect 1308 2252 1360 2304
rect 3240 2252 3292 2304
rect 5356 2388 5408 2440
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 9128 2388 9180 2440
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 10508 2388 10560 2440
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 10784 2320 10836 2372
rect 11612 2320 11664 2372
rect 13636 2320 13688 2372
rect 14464 2320 14516 2372
rect 15844 2320 15896 2372
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 7380 2295 7432 2304
rect 7380 2261 7389 2295
rect 7389 2261 7423 2295
rect 7423 2261 7432 2295
rect 7380 2252 7432 2261
rect 7748 2252 7800 2304
rect 10968 2252 11020 2304
rect 12900 2252 12952 2304
rect 21180 2388 21232 2440
rect 31300 2431 31352 2440
rect 17408 2320 17460 2372
rect 19156 2320 19208 2372
rect 21088 2320 21140 2372
rect 19248 2252 19300 2304
rect 26056 2320 26108 2372
rect 29092 2320 29144 2372
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 32864 2388 32916 2440
rect 34244 2388 34296 2440
rect 35348 2388 35400 2440
rect 28816 2252 28868 2304
rect 30932 2252 30984 2304
rect 34428 2252 34480 2304
rect 36084 2252 36136 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 7380 2048 7432 2100
rect 10876 2048 10928 2100
rect 17408 2048 17460 2100
rect 24676 2048 24728 2100
rect 21088 1980 21140 2032
rect 25596 1980 25648 2032
rect 15936 1912 15988 1964
rect 21916 1912 21968 1964
<< metal2 >>
rect 1306 39200 1362 39800
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 1320 36854 1348 39200
rect 2410 38176 2466 38185
rect 2410 38111 2466 38120
rect 2424 37330 2452 38111
rect 2412 37324 2464 37330
rect 2412 37266 2464 37272
rect 1308 36848 1360 36854
rect 1308 36790 1360 36796
rect 1320 36378 1348 36790
rect 1952 36780 2004 36786
rect 1952 36722 2004 36728
rect 1308 36372 1360 36378
rect 1308 36314 1360 36320
rect 1674 36136 1730 36145
rect 1674 36071 1676 36080
rect 1728 36071 1730 36080
rect 1676 36042 1728 36048
rect 1688 35834 1716 36042
rect 1676 35828 1728 35834
rect 1676 35770 1728 35776
rect 1676 34944 1728 34950
rect 1676 34886 1728 34892
rect 1688 34785 1716 34886
rect 1674 34776 1730 34785
rect 1674 34711 1730 34720
rect 1676 32836 1728 32842
rect 1676 32778 1728 32784
rect 1688 32745 1716 32778
rect 1674 32736 1730 32745
rect 1674 32671 1730 32680
rect 1688 32570 1716 32671
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31414 1624 31690
rect 1584 31408 1636 31414
rect 1582 31376 1584 31385
rect 1636 31376 1638 31385
rect 1582 31311 1638 31320
rect 1584 29572 1636 29578
rect 1584 29514 1636 29520
rect 1596 29345 1624 29514
rect 1582 29336 1638 29345
rect 1582 29271 1584 29280
rect 1636 29271 1638 29280
rect 1584 29242 1636 29248
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1676 26240 1728 26246
rect 1676 26182 1728 26188
rect 1688 25945 1716 26182
rect 1674 25936 1730 25945
rect 1674 25871 1730 25880
rect 1584 24132 1636 24138
rect 1584 24074 1636 24080
rect 1596 23905 1624 24074
rect 1582 23896 1638 23905
rect 1582 23831 1584 23840
rect 1636 23831 1638 23840
rect 1584 23802 1636 23808
rect 1674 22536 1730 22545
rect 1674 22471 1676 22480
rect 1728 22471 1730 22480
rect 1676 22442 1728 22448
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 20942 1624 21286
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1596 20505 1624 20878
rect 1582 20496 1638 20505
rect 1582 20431 1638 20440
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1596 19145 1624 19314
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1596 18970 1624 19071
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1688 17105 1716 17138
rect 1674 17096 1730 17105
rect 1674 17031 1730 17040
rect 1688 16794 1716 17031
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1872 16574 1900 20878
rect 1964 20602 1992 36722
rect 2424 35834 2452 37266
rect 2792 36922 2820 39471
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 3252 37126 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 6472 37262 6500 39200
rect 3516 37256 3568 37262
rect 3516 37198 3568 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 7656 37256 7708 37262
rect 7656 37198 7708 37204
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 2780 36916 2832 36922
rect 2780 36858 2832 36864
rect 2596 36644 2648 36650
rect 2596 36586 2648 36592
rect 2412 35828 2464 35834
rect 2412 35770 2464 35776
rect 2228 32836 2280 32842
rect 2228 32778 2280 32784
rect 2044 29572 2096 29578
rect 2044 29514 2096 29520
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1872 16546 1992 16574
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1872 15706 1900 16050
rect 1674 15671 1730 15680
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1676 13728 1728 13734
rect 1674 13696 1676 13705
rect 1728 13696 1730 13705
rect 1674 13631 1730 13640
rect 1872 12986 1900 13874
rect 1964 13326 1992 16546
rect 2056 15978 2084 29514
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 2148 19718 2176 22578
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1964 12238 1992 13262
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1674 11656 1730 11665
rect 1674 11591 1676 11600
rect 1728 11591 1730 11600
rect 1676 11562 1728 11568
rect 1872 10674 1900 12038
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8265 1624 8434
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1596 8090 1624 8191
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1780 5370 1808 9930
rect 1858 8392 1914 8401
rect 1858 8327 1860 8336
rect 1912 8327 1914 8336
rect 1860 8298 1912 8304
rect 2148 7478 2176 16390
rect 2240 16046 2268 32778
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2332 27878 2360 28018
rect 2320 27872 2372 27878
rect 2320 27814 2372 27820
rect 2332 21434 2360 27814
rect 2412 26308 2464 26314
rect 2412 26250 2464 26256
rect 2424 24614 2452 26250
rect 2608 26234 2636 36586
rect 3528 36582 3556 37198
rect 4804 37120 4856 37126
rect 4804 37062 4856 37068
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 3516 36576 3568 36582
rect 3516 36518 3568 36524
rect 3528 27538 3556 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3516 27532 3568 27538
rect 3516 27474 3568 27480
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2516 26206 2636 26234
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2332 21406 2452 21434
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2332 16250 2360 19654
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2228 16040 2280 16046
rect 2424 16017 2452 21406
rect 2228 15982 2280 15988
rect 2410 16008 2466 16017
rect 2410 15943 2466 15952
rect 2516 11354 2544 26206
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2596 17060 2648 17066
rect 2596 17002 2648 17008
rect 2608 15162 2636 17002
rect 2700 16454 2728 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2700 15910 2728 16050
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2700 9994 2728 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4816 12986 4844 37062
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2148 7206 2176 7414
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4865 1624 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 1582 4856 1638 4865
rect 4214 4859 4522 4868
rect 1582 4791 1584 4800
rect 1636 4791 1638 4800
rect 1584 4762 1636 4768
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2424 3097 2452 3334
rect 2410 3088 2466 3097
rect 2410 3023 2412 3032
rect 2464 3023 2466 3032
rect 2504 3052 2556 3058
rect 2412 2994 2464 3000
rect 2504 2994 2556 3000
rect 2424 2963 2452 2994
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 32 800 60 2790
rect 1872 2446 1900 2790
rect 2516 2650 2544 2994
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2792 2446 2820 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5368 2650 5396 16934
rect 6380 7886 6408 17818
rect 6748 16590 6776 37062
rect 7668 36922 7696 37198
rect 7760 37126 7788 39200
rect 9692 37262 9720 39200
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 9956 37120 10008 37126
rect 10980 37108 11008 39200
rect 12440 37324 12492 37330
rect 12440 37266 12492 37272
rect 12072 37256 12124 37262
rect 12072 37198 12124 37204
rect 11060 37120 11112 37126
rect 10980 37080 11060 37108
rect 9956 37062 10008 37068
rect 11060 37062 11112 37068
rect 7656 36916 7708 36922
rect 7656 36858 7708 36864
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 8312 36582 8340 36722
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 7564 35080 7616 35086
rect 7564 35022 7616 35028
rect 7576 27606 7604 35022
rect 7564 27600 7616 27606
rect 7564 27542 7616 27548
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 17882 6868 19178
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6748 15706 6776 16526
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 7576 15094 7604 24074
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 8128 14958 8156 27270
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8312 14890 8340 36518
rect 9968 17338 9996 37062
rect 12084 36922 12112 37198
rect 12072 36916 12124 36922
rect 12072 36858 12124 36864
rect 12452 17882 12480 37266
rect 12912 37262 12940 39200
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 14844 37126 14872 39200
rect 16132 37466 16160 39200
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 16672 37324 16724 37330
rect 16672 37266 16724 37272
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 14832 37120 14884 37126
rect 15660 37120 15712 37126
rect 14832 37062 14884 37068
rect 15658 37088 15660 37097
rect 15712 37088 15714 37097
rect 12544 36786 12572 37062
rect 15658 37023 15714 37032
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 13176 36780 13228 36786
rect 13176 36722 13228 36728
rect 13188 28082 13216 36722
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 14096 27940 14148 27946
rect 14096 27882 14148 27888
rect 14108 18358 14136 27882
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9968 16250 9996 17274
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11348 16998 11376 17138
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11164 15094 11192 15574
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 9968 14414 9996 15030
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9140 13326 9168 13874
rect 9508 13326 9536 14214
rect 11072 13802 11100 14214
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12306 8340 12786
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8404 12238 8432 12922
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11082 8064 12038
rect 8680 11898 8708 12174
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7944 10810 7972 11018
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5368 2446 5396 2586
rect 5552 2582 5580 3402
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 6564 2446 6592 7686
rect 8220 6458 8248 11494
rect 8772 10810 8800 11698
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 3534 7880 6054
rect 9140 5846 9168 13262
rect 9508 12850 9536 13262
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9876 12434 9904 12786
rect 10704 12442 10732 13670
rect 10980 13530 11008 13738
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10796 12753 10824 13194
rect 10782 12744 10838 12753
rect 10782 12679 10838 12688
rect 10692 12436 10744 12442
rect 9876 12406 9996 12434
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10266 9444 10406
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 9042 9444 9318
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9416 5914 9444 6666
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9140 4826 9168 5782
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9140 4622 9168 4762
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8588 3126 8616 3334
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 9140 2446 9168 3334
rect 9600 3058 9628 12038
rect 9876 11354 9904 12174
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 9058 9720 11018
rect 9876 10538 9904 11290
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 9926 9812 10066
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9178 9812 9862
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9692 9030 9812 9058
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8362 9720 8910
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9692 7206 9720 8298
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9784 6866 9812 9030
rect 9968 8906 9996 12406
rect 10692 12378 10744 12384
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11762 10732 12174
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10060 11257 10088 11494
rect 10428 11354 10456 11494
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10704 11286 10732 11698
rect 10692 11280 10744 11286
rect 10046 11248 10102 11257
rect 10692 11222 10744 11228
rect 10046 11183 10102 11192
rect 10060 11150 10088 11183
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10508 10736 10560 10742
rect 10506 10704 10508 10713
rect 10560 10704 10562 10713
rect 10140 10668 10192 10674
rect 10506 10639 10562 10648
rect 10140 10610 10192 10616
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 10152 8566 10180 10610
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10520 9178 10548 9454
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10796 8566 10824 12679
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10888 11082 10916 11562
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10980 9382 11008 13466
rect 11072 13258 11100 13738
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 11762 11100 12038
rect 11164 11898 11192 12174
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11150 11792 11206 11801
rect 11060 11756 11112 11762
rect 11150 11727 11206 11736
rect 11060 11698 11112 11704
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10968 9376 11020 9382
rect 10966 9344 10968 9353
rect 11020 9344 11022 9353
rect 10966 9279 11022 9288
rect 10980 9253 11008 9279
rect 11072 9110 11100 11222
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10152 7478 10180 8502
rect 10704 8090 10732 8502
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10152 6866 10180 7414
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9784 6458 9812 6802
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9692 5166 9720 6190
rect 9784 5386 9812 6394
rect 9784 5358 9904 5386
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9692 3194 9720 5102
rect 9784 4826 9812 5238
rect 9876 5166 9904 5358
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9508 2774 9536 2926
rect 9508 2746 9720 2774
rect 9508 2446 9536 2746
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 2792 1465 2820 2382
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 7392 2106 7420 2246
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7760 800 7788 2246
rect 9692 800 9720 2746
rect 10520 2446 10548 7890
rect 10796 4146 10824 7958
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 7002 11008 7414
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11072 5370 11100 7686
rect 11164 6746 11192 11727
rect 11256 10606 11284 14554
rect 11348 14482 11376 16934
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16250 12572 16390
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11624 15609 11652 15914
rect 11610 15600 11666 15609
rect 12360 15570 12388 16186
rect 12622 16144 12678 16153
rect 12622 16079 12624 16088
rect 12676 16079 12678 16088
rect 12624 16050 12676 16056
rect 11610 15535 11666 15544
rect 12348 15564 12400 15570
rect 11624 15502 11652 15535
rect 12348 15506 12400 15512
rect 12728 15502 12756 18226
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 16658 13032 17478
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13096 16590 13124 17070
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16046 13032 16390
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11348 14278 11376 14418
rect 11704 14408 11756 14414
rect 11702 14376 11704 14385
rect 11756 14376 11758 14385
rect 11624 14334 11702 14362
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 12238 11376 14214
rect 11624 13938 11652 14334
rect 11702 14311 11758 14320
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11428 12912 11480 12918
rect 11426 12880 11428 12889
rect 11480 12880 11482 12889
rect 11426 12815 11482 12824
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11532 11830 11560 13806
rect 11716 13530 11744 13874
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11624 12345 11652 12786
rect 11808 12764 11836 14962
rect 11992 13682 12020 15302
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12360 14278 12388 14350
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12348 13864 12400 13870
rect 12544 13852 12572 14282
rect 12636 14006 12664 15302
rect 13188 14634 13216 17818
rect 13280 17202 13308 18022
rect 13452 17672 13504 17678
rect 13504 17620 13584 17626
rect 13452 17614 13584 17620
rect 13464 17598 13584 17614
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13372 16114 13400 17002
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16794 13492 16934
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13464 16046 13492 16730
rect 13556 16674 13584 17598
rect 14108 17202 14136 18294
rect 14292 17678 14320 18906
rect 14476 18426 14504 27406
rect 16684 22094 16712 37266
rect 18064 37126 18092 39200
rect 19352 37330 19380 39200
rect 19340 37324 19392 37330
rect 19340 37266 19392 37272
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18524 36582 18552 37198
rect 19352 36922 19380 37266
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19996 36786 20024 37198
rect 21284 37126 21312 39200
rect 22008 37256 22060 37262
rect 22008 37198 22060 37204
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 20260 36780 20312 36786
rect 20260 36722 20312 36728
rect 18512 36576 18564 36582
rect 18512 36518 18564 36524
rect 17592 36032 17644 36038
rect 17592 35974 17644 35980
rect 16684 22066 16896 22094
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15304 21622 15332 21830
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 15396 20602 15424 21558
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18766 14596 19110
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14660 18578 14688 19790
rect 15212 18766 15240 20402
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 14568 18550 14688 18578
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14200 17066 14228 17138
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 13726 16688 13782 16697
rect 13556 16646 13726 16674
rect 13726 16623 13782 16632
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13464 15366 13492 15982
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13648 15473 13676 15506
rect 13740 15502 13768 16623
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13728 15496 13780 15502
rect 13634 15464 13690 15473
rect 13728 15438 13780 15444
rect 13634 15399 13690 15408
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13544 14952 13596 14958
rect 13542 14920 13544 14929
rect 13596 14920 13598 14929
rect 13542 14855 13598 14864
rect 13636 14816 13688 14822
rect 13688 14764 13768 14770
rect 13636 14758 13768 14764
rect 13648 14742 13768 14758
rect 13096 14606 13216 14634
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12624 13864 12676 13870
rect 12400 13824 12480 13852
rect 12544 13824 12624 13852
rect 12348 13806 12400 13812
rect 12348 13728 12400 13734
rect 11992 13654 12296 13682
rect 12348 13670 12400 13676
rect 11992 13258 12020 13654
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 12084 12986 12112 13466
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11900 12866 11928 12922
rect 11900 12850 12112 12866
rect 11900 12844 12124 12850
rect 11900 12838 12072 12844
rect 12072 12786 12124 12792
rect 11808 12736 12020 12764
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11794 12336 11850 12345
rect 11794 12271 11850 12280
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11336 11824 11388 11830
rect 11520 11824 11572 11830
rect 11388 11784 11468 11812
rect 11336 11766 11388 11772
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11348 7478 11376 11222
rect 11440 9738 11468 11784
rect 11520 11766 11572 11772
rect 11440 9710 11560 9738
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11440 9178 11468 9590
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11532 7002 11560 9710
rect 11624 8362 11652 12174
rect 11808 11694 11836 12271
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 9586 11744 10950
rect 11808 10674 11836 11630
rect 11900 11218 11928 12174
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11992 11132 12020 12736
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 12306 12112 12582
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12176 12186 12204 13330
rect 12268 12866 12296 13654
rect 12360 12986 12388 13670
rect 12452 13172 12480 13824
rect 12624 13806 12676 13812
rect 12728 13462 12756 14282
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12912 13326 12940 14418
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12624 13184 12676 13190
rect 12452 13144 12624 13172
rect 12624 13126 12676 13132
rect 13004 13002 13032 13670
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12452 12974 13032 13002
rect 12268 12838 12388 12866
rect 12360 12782 12388 12838
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12452 12714 12480 12974
rect 12900 12912 12952 12918
rect 12898 12880 12900 12889
rect 12952 12880 12954 12889
rect 12898 12815 12954 12824
rect 12530 12744 12586 12753
rect 12440 12708 12492 12714
rect 12530 12679 12532 12688
rect 12440 12650 12492 12656
rect 12584 12679 12586 12688
rect 12532 12650 12584 12656
rect 13096 12442 13124 14606
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 12782 13400 13330
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12256 12368 12308 12374
rect 12254 12336 12256 12345
rect 12308 12336 12310 12345
rect 12254 12271 12310 12280
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12084 12158 12204 12186
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12084 11694 12112 12158
rect 12360 12050 12388 12174
rect 12176 12022 12388 12050
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 11286 12112 11630
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 11992 11104 12112 11132
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11900 10062 11928 10678
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10266 12020 10542
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11900 9674 11928 9998
rect 11808 9646 11928 9674
rect 11980 9648 12032 9654
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11808 9466 11836 9646
rect 11980 9590 12032 9596
rect 11716 9438 11836 9466
rect 11716 8974 11744 9438
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11164 6718 11652 6746
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10796 3466 10824 4082
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 11072 3126 11100 5306
rect 11164 3466 11192 5646
rect 11256 4010 11284 6598
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11440 5914 11468 6326
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11532 5710 11560 6054
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11348 4146 11376 4762
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11624 3738 11652 6718
rect 11716 6118 11744 8910
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11808 5642 11836 8910
rect 11992 8634 12020 9590
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11716 4690 11744 5306
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11532 3126 11560 3470
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 10874 2544 10930 2553
rect 11532 2514 11560 3062
rect 10874 2479 10930 2488
rect 11520 2508 11572 2514
rect 10888 2446 10916 2479
rect 11520 2450 11572 2456
rect 10508 2440 10560 2446
rect 10876 2440 10928 2446
rect 10508 2382 10560 2388
rect 10782 2408 10838 2417
rect 10876 2382 10928 2388
rect 10782 2343 10784 2352
rect 10836 2343 10838 2352
rect 10784 2314 10836 2320
rect 10888 2106 10916 2382
rect 11624 2378 11652 3674
rect 11900 3602 11928 7822
rect 12084 7546 12112 11104
rect 12176 9926 12204 12022
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12360 11098 12388 11834
rect 12452 11830 12480 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12268 11082 12388 11098
rect 12256 11076 12388 11082
rect 12308 11070 12388 11076
rect 12256 11018 12308 11024
rect 12544 10470 12572 12038
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12268 9518 12296 9998
rect 12544 9654 12572 10406
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12176 9178 12204 9454
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 6866 12020 7278
rect 12084 7206 12112 7482
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11992 6458 12020 6802
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11992 5778 12020 6394
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11992 5250 12020 5578
rect 12084 5370 12112 6938
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11992 5222 12112 5250
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 11808 3398 11836 3431
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11900 2990 11928 3538
rect 11992 3534 12020 4014
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11888 2984 11940 2990
rect 12084 2961 12112 5222
rect 12176 4826 12204 9114
rect 12636 8090 12664 11086
rect 12728 9450 12756 11630
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 10198 12940 10610
rect 13004 10266 13032 11018
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 13096 9722 13124 10746
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12728 9042 12756 9386
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12728 8430 12756 8842
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12348 6112 12400 6118
rect 12452 6066 12480 6598
rect 12400 6060 12480 6066
rect 12348 6054 12480 6060
rect 12360 6038 12480 6054
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12268 4214 12296 5850
rect 12544 4298 12572 7482
rect 13188 4865 13216 12242
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 11218 13308 11630
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 9110 13308 11154
rect 13372 11014 13400 12718
rect 13464 12306 13492 14010
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13556 12170 13584 13330
rect 13648 12646 13676 13806
rect 13740 13462 13768 14742
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12238 13676 12582
rect 13740 12442 13768 12650
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13648 11830 13676 12174
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13648 11150 13676 11562
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8634 13400 8774
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13464 6746 13492 9998
rect 13556 8974 13584 10134
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8566 13584 8910
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13556 7478 13584 8026
rect 13648 7546 13676 10406
rect 13832 8634 13860 15030
rect 13924 11354 13952 16458
rect 14200 16153 14228 17002
rect 14370 16960 14426 16969
rect 14370 16895 14426 16904
rect 14186 16144 14242 16153
rect 14384 16114 14412 16895
rect 14186 16079 14242 16088
rect 14372 16108 14424 16114
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 14958 14136 15302
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14016 14550 14044 14894
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14016 14006 14044 14486
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14002 13424 14058 13433
rect 14002 13359 14004 13368
rect 14056 13359 14058 13368
rect 14004 13330 14056 13336
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 9761 14044 10542
rect 14002 9752 14058 9761
rect 14002 9687 14058 9696
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14016 9353 14044 9522
rect 14002 9344 14058 9353
rect 14002 9279 14058 9288
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 14002 8528 14058 8537
rect 13820 8492 13872 8498
rect 14002 8463 14004 8472
rect 13820 8434 13872 8440
rect 14056 8463 14058 8472
rect 14004 8434 14056 8440
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13556 6866 13584 7414
rect 13740 7410 13768 7754
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13464 6718 13584 6746
rect 13556 5710 13584 6718
rect 13726 6352 13782 6361
rect 13726 6287 13728 6296
rect 13780 6287 13782 6296
rect 13728 6258 13780 6264
rect 13832 6254 13860 8434
rect 14108 7886 14136 13874
rect 14200 11218 14228 16079
rect 14372 16050 14424 16056
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14384 14618 14412 15030
rect 14464 14952 14516 14958
rect 14462 14920 14464 14929
rect 14516 14920 14518 14929
rect 14462 14855 14518 14864
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14292 12073 14320 12718
rect 14278 12064 14334 12073
rect 14278 11999 14334 12008
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 6390 13952 6598
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13634 5672 13690 5681
rect 13556 5114 13584 5646
rect 13634 5607 13636 5616
rect 13688 5607 13690 5616
rect 13636 5578 13688 5584
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13280 5086 13584 5114
rect 13174 4856 13230 4865
rect 13174 4791 13230 4800
rect 12990 4720 13046 4729
rect 12990 4655 13046 4664
rect 12237 4208 12296 4214
rect 12289 4168 12296 4208
rect 12452 4270 12572 4298
rect 12237 4150 12289 4156
rect 12452 3738 12480 4270
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 13004 3126 13032 4655
rect 13280 4282 13308 5086
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13556 4214 13584 4966
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13452 4072 13504 4078
rect 13740 4026 13768 5510
rect 13832 4078 13860 6190
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13924 5914 13952 6122
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5914 14044 6054
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14108 5846 14136 7822
rect 14200 7342 14228 10950
rect 14292 9178 14320 11999
rect 14384 11762 14412 13738
rect 14568 12434 14596 18550
rect 14752 17202 14780 18566
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 15028 16726 15056 18362
rect 15304 18358 15332 19654
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15384 19236 15436 19242
rect 15384 19178 15436 19184
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15396 18222 15424 19178
rect 15488 18970 15516 19450
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15120 17134 15148 18158
rect 15396 17814 15424 18158
rect 15384 17808 15436 17814
rect 15384 17750 15436 17756
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14476 12406 14596 12434
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14476 11014 14504 12406
rect 14660 11914 14688 15846
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14844 15434 14872 15574
rect 14832 15428 14884 15434
rect 14832 15370 14884 15376
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14752 14414 14780 14554
rect 14740 14408 14792 14414
rect 15028 14396 15056 16390
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 15120 15434 15148 15914
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15212 15008 15240 16730
rect 15304 16046 15332 17682
rect 15488 17610 15516 18566
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15580 16794 15608 17546
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15384 15020 15436 15026
rect 15212 14980 15384 15008
rect 15384 14962 15436 14968
rect 15028 14368 15148 14396
rect 14740 14350 14792 14356
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 15028 13258 15056 13738
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14832 12912 14884 12918
rect 14884 12860 15056 12866
rect 14832 12854 15056 12860
rect 14844 12838 15056 12854
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14568 11886 14688 11914
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 7002 14320 7142
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14016 4826 14044 5170
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13452 4014 13504 4020
rect 13464 3126 13492 4014
rect 13556 3998 13768 4026
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13556 3641 13584 3998
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13648 3670 13676 3878
rect 13740 3738 13768 3878
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13636 3664 13688 3670
rect 13542 3632 13598 3641
rect 13636 3606 13688 3612
rect 13542 3567 13598 3576
rect 14200 3534 14228 6870
rect 14384 6254 14412 9998
rect 14476 6866 14504 10542
rect 14568 10010 14596 11886
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14660 10130 14688 11766
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14568 9982 14688 10010
rect 14556 9920 14608 9926
rect 14554 9888 14556 9897
rect 14608 9888 14610 9897
rect 14554 9823 14610 9832
rect 14660 9382 14688 9982
rect 14752 9654 14780 12106
rect 14832 10736 14884 10742
rect 14830 10704 14832 10713
rect 14884 10704 14886 10713
rect 14830 10639 14886 10648
rect 15028 10441 15056 12838
rect 14830 10432 14886 10441
rect 14830 10367 14886 10376
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14476 6458 14504 6802
rect 14568 6662 14596 7278
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14384 5302 14412 6190
rect 14476 5302 14504 6394
rect 14568 5574 14596 6598
rect 14660 6254 14688 9318
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14752 8809 14780 8910
rect 14738 8800 14794 8809
rect 14738 8735 14794 8744
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14844 5302 14872 10367
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 7002 14964 8842
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14936 5846 14964 6938
rect 15028 6186 15056 8910
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14188 3528 14240 3534
rect 14280 3528 14332 3534
rect 14188 3470 14240 3476
rect 14278 3496 14280 3505
rect 14332 3496 14334 3505
rect 14278 3431 14334 3440
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13464 2961 13492 3062
rect 11888 2926 11940 2932
rect 12070 2952 12126 2961
rect 12070 2887 12126 2896
rect 12714 2952 12770 2961
rect 12714 2887 12770 2896
rect 13450 2952 13506 2961
rect 13450 2887 13506 2896
rect 12728 2854 12756 2887
rect 12440 2848 12492 2854
rect 12438 2816 12440 2825
rect 12716 2848 12768 2854
rect 12492 2816 12494 2825
rect 14476 2825 14504 3946
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3602 14596 3878
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 12716 2790 12768 2796
rect 14462 2816 14518 2825
rect 12438 2751 12494 2760
rect 14462 2751 14518 2760
rect 13634 2680 13690 2689
rect 13634 2615 13690 2624
rect 13648 2378 13676 2615
rect 14476 2378 14504 2751
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10980 800 11008 2246
rect 12912 800 12940 2246
rect 14844 800 14872 3334
rect 14936 3210 14964 4422
rect 15120 3602 15148 14368
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15212 12374 15240 12718
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15212 11014 15240 11154
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 7002 15240 10950
rect 15304 9518 15332 11630
rect 15396 9994 15424 14962
rect 15488 14550 15516 15370
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15476 14340 15528 14346
rect 15528 14300 15608 14328
rect 15476 14282 15528 14288
rect 15580 13433 15608 14300
rect 15566 13424 15622 13433
rect 15566 13359 15568 13368
rect 15620 13359 15622 13368
rect 15568 13330 15620 13336
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15488 12102 15516 12854
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15568 10260 15620 10266
rect 15672 10248 15700 18294
rect 15856 18086 15884 18906
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 17202 15884 18022
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15856 15978 15884 16458
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 15764 15706 15792 15914
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15856 15502 15884 15914
rect 15948 15910 15976 18702
rect 16040 17105 16068 19314
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16132 18766 16160 19110
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16132 17338 16160 17750
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16316 17338 16344 17546
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16026 17096 16082 17105
rect 16026 17031 16082 17040
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 16040 15722 16068 17031
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 15910 16252 16934
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 15948 15694 16068 15722
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15948 14090 15976 15694
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16040 14278 16068 15302
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15948 14062 16068 14090
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15764 11898 15792 13942
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15856 13258 15884 13398
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15856 11762 15884 12718
rect 16040 12434 16068 14062
rect 16132 12646 16160 15302
rect 16408 15026 16436 18226
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17626 16528 18022
rect 16500 17598 16620 17626
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16210 14376 16266 14385
rect 16210 14311 16266 14320
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16040 12406 16160 12434
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 12102 16068 12174
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15620 10220 15700 10248
rect 15568 10202 15620 10208
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15396 8634 15424 9930
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15672 9625 15700 9658
rect 15658 9616 15714 9625
rect 15658 9551 15714 9560
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15488 8294 15516 8978
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15580 7154 15608 9318
rect 15672 8838 15700 9454
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15488 7126 15608 7154
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15488 4758 15516 7126
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15580 5778 15608 6938
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15764 5370 15792 11494
rect 15842 10704 15898 10713
rect 15842 10639 15898 10648
rect 15856 9722 15884 10639
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 8514 15884 9318
rect 15948 9178 15976 12038
rect 16028 10464 16080 10470
rect 16026 10432 16028 10441
rect 16080 10432 16082 10441
rect 16026 10367 16082 10376
rect 16040 10266 16068 10367
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16040 8838 16068 8910
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15934 8664 15990 8673
rect 15934 8599 15936 8608
rect 15988 8599 15990 8608
rect 15936 8570 15988 8576
rect 16028 8560 16080 8566
rect 15856 8508 16028 8514
rect 15856 8502 16080 8508
rect 15856 8486 16068 8502
rect 16028 8288 16080 8294
rect 16132 8242 16160 12406
rect 16224 11762 16252 14311
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16408 13394 16436 14010
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16500 13190 16528 17478
rect 16592 15722 16620 17598
rect 16684 16998 16712 21558
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18358 16804 18566
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16776 17066 16804 17138
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16658 16712 16934
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16868 16538 16896 22066
rect 17604 21894 17632 35974
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17604 20942 17632 21830
rect 17880 21622 17908 22986
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16960 17338 16988 20470
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17052 17610 17080 19314
rect 17236 19310 17264 20742
rect 18524 20262 18552 36518
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20272 28082 20300 36722
rect 22020 35290 22048 37198
rect 22572 37126 22600 39200
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22560 37120 22612 37126
rect 22560 37062 22612 37068
rect 22008 35284 22060 35290
rect 22008 35226 22060 35232
rect 22756 32570 22784 37198
rect 24504 37126 24532 39200
rect 26436 37466 26464 39200
rect 26424 37460 26476 37466
rect 26424 37402 26476 37408
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 24400 34944 24452 34950
rect 24400 34886 24452 34892
rect 24412 34542 24440 34886
rect 24400 34536 24452 34542
rect 24400 34478 24452 34484
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22020 31822 22048 32370
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 21468 23186 21496 27814
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21622 20024 22374
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18222 17264 19246
rect 17328 18970 17356 19382
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17236 17746 17264 18158
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17696 16726 17724 19654
rect 17972 19174 18000 19722
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17684 16720 17736 16726
rect 16946 16688 17002 16697
rect 17684 16662 17736 16668
rect 16946 16623 16948 16632
rect 17000 16623 17002 16632
rect 16948 16594 17000 16600
rect 17696 16590 17724 16662
rect 17684 16584 17736 16590
rect 16868 16510 17080 16538
rect 17684 16526 17736 16532
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16592 15694 16896 15722
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16592 14328 16620 15574
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16776 14482 16804 14826
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 14340 16724 14346
rect 16592 14300 16672 14328
rect 16672 14282 16724 14288
rect 16684 13258 16712 14282
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16316 12442 16344 13126
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16684 12170 16712 12310
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16080 8236 16160 8242
rect 16028 8230 16160 8236
rect 16040 8214 16160 8230
rect 16132 7750 16160 8214
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15566 5128 15622 5137
rect 15856 5098 15884 5646
rect 16132 5234 16160 7686
rect 16224 5370 16252 11698
rect 16592 11354 16620 12106
rect 16776 11898 16804 13806
rect 16868 12918 16896 15694
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16868 11694 16896 12106
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16960 11234 16988 16390
rect 17052 13734 17080 16510
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17222 15464 17278 15473
rect 17328 15434 17356 15642
rect 17222 15399 17224 15408
rect 17276 15399 17278 15408
rect 17316 15428 17368 15434
rect 17224 15370 17276 15376
rect 17316 15370 17368 15376
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17144 14890 17172 15098
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16592 11218 16988 11234
rect 16580 11212 16988 11218
rect 16632 11206 16988 11212
rect 17052 13240 17080 13670
rect 17236 13274 17264 14962
rect 17788 14482 17816 16730
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 14958 17908 15302
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17696 14006 17724 14418
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17420 13530 17448 13942
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17592 13320 17644 13326
rect 17132 13252 17184 13258
rect 17052 13212 17132 13240
rect 16580 11154 16632 11160
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16316 10470 16344 10746
rect 16960 10674 16988 11086
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16592 10130 16620 10542
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 9518 16620 10066
rect 16670 9616 16726 9625
rect 16670 9551 16726 9560
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16592 8838 16620 9454
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 8430 16620 8774
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16592 7954 16620 8366
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16302 5808 16358 5817
rect 16302 5743 16358 5752
rect 16316 5642 16344 5743
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15566 5063 15622 5072
rect 15844 5092 15896 5098
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15580 4554 15608 5063
rect 15844 5034 15896 5040
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15660 4684 15712 4690
rect 15764 4672 15792 4966
rect 15712 4644 15792 4672
rect 15660 4626 15712 4632
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15580 4214 15608 4490
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15764 3516 15792 4644
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 4282 15884 4422
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15844 3528 15896 3534
rect 15764 3488 15844 3516
rect 15844 3470 15896 3476
rect 15016 3460 15068 3466
rect 15292 3460 15344 3466
rect 15068 3420 15292 3448
rect 15016 3402 15068 3408
rect 15292 3402 15344 3408
rect 15014 3224 15070 3233
rect 14936 3182 15014 3210
rect 15856 3194 15884 3470
rect 15014 3159 15070 3168
rect 15844 3188 15896 3194
rect 15028 3126 15056 3159
rect 15844 3130 15896 3136
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15856 2378 15884 2586
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 15948 1970 15976 4490
rect 16224 4282 16252 5306
rect 16488 5296 16540 5302
rect 16486 5264 16488 5273
rect 16540 5264 16542 5273
rect 16486 5199 16542 5208
rect 16684 5098 16712 9551
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16408 4690 16436 5034
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3194 16344 4082
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16408 3126 16436 4626
rect 16776 3942 16804 10134
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16868 8809 16896 9930
rect 17052 9654 17080 13212
rect 17236 13246 17356 13274
rect 17880 13274 17908 14894
rect 17972 14822 18000 18634
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18340 18154 18368 18566
rect 18616 18290 18644 18566
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17270 18092 18022
rect 18156 17610 18184 18090
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16969 18184 17070
rect 18142 16960 18198 16969
rect 18142 16895 18198 16904
rect 18156 16250 18184 16895
rect 18248 16726 18276 17478
rect 18236 16720 18288 16726
rect 18236 16662 18288 16668
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 18064 15162 18092 16118
rect 18510 16008 18566 16017
rect 18510 15943 18512 15952
rect 18564 15943 18566 15952
rect 18512 15914 18564 15920
rect 18144 15904 18196 15910
rect 18616 15858 18644 18226
rect 18708 16590 18736 19722
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18800 18834 18828 19178
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18144 15846 18196 15852
rect 18156 15434 18184 15846
rect 18524 15830 18644 15858
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18248 15094 18276 15506
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14346 18368 14758
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18248 13802 18276 13942
rect 18432 13870 18460 14418
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 17592 13262 17644 13268
rect 17132 13194 17184 13200
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17130 12608 17186 12617
rect 17130 12543 17186 12552
rect 17144 11218 17172 12543
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17236 10742 17264 12854
rect 17328 12481 17356 13246
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17314 12472 17370 12481
rect 17370 12416 17448 12434
rect 17314 12407 17448 12416
rect 17328 12406 17448 12407
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17038 9480 17094 9489
rect 17038 9415 17040 9424
rect 17092 9415 17094 9424
rect 17040 9386 17092 9392
rect 16854 8800 16910 8809
rect 16854 8735 16910 8744
rect 16868 8566 16896 8735
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 17144 7528 17172 10474
rect 17236 7954 17264 10678
rect 17328 9994 17356 11018
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 9110 17356 9522
rect 17420 9382 17448 12406
rect 17512 11286 17540 12854
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17052 7500 17172 7528
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16868 4282 16896 6190
rect 16960 6118 16988 6666
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 17052 4622 17080 7500
rect 17236 7478 17264 7890
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17512 6866 17540 11086
rect 17604 10130 17632 13262
rect 17696 13246 17908 13274
rect 17696 10198 17724 13246
rect 17972 12782 18000 13738
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12889 18184 13126
rect 18432 12918 18460 13670
rect 18420 12912 18472 12918
rect 18142 12880 18198 12889
rect 18420 12854 18472 12860
rect 18142 12815 18198 12824
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 18524 12434 18552 15830
rect 18800 15722 18828 18362
rect 19168 17678 19196 19110
rect 19352 17746 19380 20334
rect 19444 19310 19472 21422
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19628 20058 19656 20470
rect 20088 20398 20116 22918
rect 21008 22778 21036 22986
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21468 22098 21496 23122
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20732 21622 20760 21830
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 21928 21486 21956 26250
rect 22020 23254 22048 31758
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23860 22094 23888 22374
rect 23860 22066 23980 22094
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 22848 21690 22876 21898
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21146 20852 21286
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20904 20868 20956 20874
rect 20904 20810 20956 20816
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 20916 20602 20944 20810
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20916 19446 20944 19790
rect 21008 19514 21036 20810
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21468 19446 21496 19654
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 18878 17096 18934 17105
rect 18878 17031 18880 17040
rect 18932 17031 18934 17040
rect 18880 17002 18932 17008
rect 19168 16574 19196 17614
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19260 17270 19288 17478
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19168 16546 19380 16574
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18892 16114 18920 16458
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18432 12406 18552 12434
rect 18616 15694 18828 15722
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 11558 17908 11698
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17682 10024 17738 10033
rect 17682 9959 17738 9968
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 8566 17632 9862
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17604 7886 17632 8502
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17696 7818 17724 9959
rect 17788 9518 17816 11222
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17774 8664 17830 8673
rect 17774 8599 17776 8608
rect 17828 8599 17830 8608
rect 17776 8570 17828 8576
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17880 7478 17908 11494
rect 17972 11082 18000 11630
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 8566 18000 10406
rect 18064 10198 18092 11290
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 9926 18092 9998
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 8906 18092 9318
rect 18156 9178 18184 9590
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17880 6934 17908 7414
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17144 6458 17172 6598
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17420 4826 17448 6258
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17604 5778 17632 6190
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17604 5234 17632 5714
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17880 4690 17908 5714
rect 17972 5370 18000 8366
rect 18064 6866 18092 8842
rect 18156 8430 18184 8842
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18248 6730 18276 11222
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10266 18368 10950
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18340 9897 18368 9930
rect 18326 9888 18382 9897
rect 18326 9823 18382 9832
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 18340 5846 18368 8978
rect 18432 7206 18460 12406
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18524 9042 18552 11630
rect 18616 9466 18644 15694
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18708 12220 18736 14962
rect 18892 13530 18920 16050
rect 19260 15994 19288 16186
rect 19352 16153 19380 16546
rect 19338 16144 19394 16153
rect 19338 16079 19394 16088
rect 19340 16040 19392 16046
rect 19260 15988 19340 15994
rect 19260 15982 19392 15988
rect 19260 15966 19380 15982
rect 19260 15434 19288 15966
rect 19444 15638 19472 18294
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19352 14362 19380 15438
rect 19444 14872 19472 15574
rect 19536 15502 19564 15982
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19708 14884 19760 14890
rect 19444 14844 19708 14872
rect 19708 14826 19760 14832
rect 19352 14334 19472 14362
rect 19340 14272 19392 14278
rect 19338 14240 19340 14249
rect 19392 14240 19394 14249
rect 19338 14175 19394 14184
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 18880 13524 18932 13530
rect 18800 13484 18880 13512
rect 18800 12288 18828 13484
rect 18880 13466 18932 13472
rect 18984 12986 19012 13942
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12646 18920 12786
rect 19076 12714 19104 13942
rect 19340 13320 19392 13326
rect 19338 13288 19340 13297
rect 19392 13288 19394 13297
rect 19338 13223 19394 13232
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12434 19012 12582
rect 18984 12406 19104 12434
rect 18800 12260 19012 12288
rect 18708 12192 18920 12220
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18800 11694 18828 12038
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18800 10062 18828 11018
rect 18892 10266 18920 12192
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18984 10146 19012 12260
rect 18892 10118 19012 10146
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18892 9874 18920 10118
rect 18800 9846 18920 9874
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18616 9438 18736 9466
rect 18708 9382 18736 9438
rect 18696 9376 18748 9382
rect 18602 9344 18658 9353
rect 18696 9318 18748 9324
rect 18602 9279 18658 9288
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18524 6730 18552 7822
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18524 6186 18552 6666
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18524 5846 18552 6122
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 18052 5636 18104 5642
rect 18052 5578 18104 5584
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18064 4758 18092 5578
rect 18052 4752 18104 4758
rect 18236 4752 18288 4758
rect 18052 4694 18104 4700
rect 18234 4720 18236 4729
rect 18288 4720 18290 4729
rect 17868 4684 17920 4690
rect 18234 4655 18290 4664
rect 17868 4626 17920 4632
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16868 4146 16896 4218
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16868 3058 16896 3538
rect 17144 3194 17172 4014
rect 18340 3602 18368 5782
rect 18524 5302 18552 5782
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18512 4208 18564 4214
rect 18510 4176 18512 4185
rect 18564 4176 18566 4185
rect 18510 4111 18566 4120
rect 18616 3652 18644 9279
rect 18800 6066 18828 9846
rect 18878 9480 18934 9489
rect 18878 9415 18934 9424
rect 18892 9382 18920 9415
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18892 6186 18920 7142
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18800 6038 18920 6066
rect 18786 4856 18842 4865
rect 18786 4791 18788 4800
rect 18840 4791 18842 4800
rect 18788 4762 18840 4768
rect 18800 4690 18828 4762
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 4282 18736 4422
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18696 3664 18748 3670
rect 18616 3624 18696 3652
rect 18696 3606 18748 3612
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16578 2952 16634 2961
rect 16578 2887 16634 2896
rect 16304 2848 16356 2854
rect 16132 2796 16304 2802
rect 16132 2790 16356 2796
rect 16132 2774 16344 2790
rect 15936 1964 15988 1970
rect 15936 1906 15988 1912
rect 16132 800 16160 2774
rect 16592 2582 16620 2887
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 17880 2514 17908 3062
rect 18616 2854 18644 3334
rect 18708 2990 18736 3606
rect 18892 3097 18920 6038
rect 18984 3505 19012 9862
rect 19076 8022 19104 12406
rect 19246 12336 19302 12345
rect 19246 12271 19248 12280
rect 19300 12271 19302 12280
rect 19248 12242 19300 12248
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 8016 19116 8022
rect 19064 7958 19116 7964
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19076 6730 19104 7346
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19076 4146 19104 4558
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19076 3738 19104 4082
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18970 3496 19026 3505
rect 18970 3431 19026 3440
rect 19076 3126 19104 3674
rect 19064 3120 19116 3126
rect 18878 3088 18934 3097
rect 19064 3062 19116 3068
rect 18878 3023 18934 3032
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17420 2106 17448 2314
rect 17408 2100 17460 2106
rect 17408 2042 17460 2048
rect 18064 800 18092 2790
rect 19168 2378 19196 12174
rect 19248 12096 19300 12102
rect 19246 12064 19248 12073
rect 19300 12064 19302 12073
rect 19246 11999 19302 12008
rect 19352 10810 19380 13126
rect 19444 12850 19472 14334
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13394 19564 13806
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19812 13394 19840 13738
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19890 12880 19946 12889
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19536 12306 19564 12854
rect 19890 12815 19946 12824
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19812 12374 19840 12650
rect 19904 12646 19932 12815
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11336 19472 12174
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11370 20024 18634
rect 20088 16538 20116 19110
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18358 20300 18566
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20180 17882 20208 18158
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20180 17746 20208 17818
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 20180 17338 20208 17682
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20364 17202 20392 17546
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20364 16998 20392 17138
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20548 16658 20576 18838
rect 20640 16794 20668 19314
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20824 18086 20852 18906
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20824 17678 20852 18022
rect 20812 17672 20864 17678
rect 20810 17640 20812 17649
rect 20864 17640 20866 17649
rect 20810 17575 20866 17584
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 17270 20760 17478
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20916 16794 20944 17206
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20088 16522 20208 16538
rect 20088 16516 20220 16522
rect 20088 16510 20168 16516
rect 20168 16458 20220 16464
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 15094 20116 16390
rect 20180 15502 20208 16458
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20180 14346 20208 15302
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 14074 20116 14214
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20272 13954 20300 16594
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20350 16144 20406 16153
rect 20350 16079 20352 16088
rect 20404 16079 20406 16088
rect 20352 16050 20404 16056
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20364 15366 20392 15914
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20088 13926 20300 13954
rect 20088 13802 20116 13926
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 20166 12744 20222 12753
rect 20166 12679 20222 12688
rect 20180 12322 20208 12679
rect 20272 12345 20300 13806
rect 20350 13424 20406 13433
rect 20350 13359 20406 13368
rect 20088 12294 20208 12322
rect 20258 12336 20314 12345
rect 20088 11558 20116 12294
rect 20258 12271 20314 12280
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19996 11342 20116 11370
rect 19444 11308 19564 11336
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19248 10736 19300 10742
rect 19246 10704 19248 10713
rect 19300 10704 19302 10713
rect 19246 10639 19302 10648
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19260 7886 19288 9386
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19352 6798 19380 10134
rect 19444 8430 19472 11154
rect 19536 11014 19564 11308
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19614 10568 19670 10577
rect 19614 10503 19616 10512
rect 19668 10503 19670 10512
rect 19616 10474 19668 10480
rect 19996 10470 20024 11154
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19982 10296 20038 10305
rect 19982 10231 20038 10240
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9382 20024 10231
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 20088 9178 20116 11342
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20180 10062 20208 10746
rect 20272 10742 20300 12174
rect 20364 11014 20392 13359
rect 20456 12646 20484 16458
rect 20548 15570 20576 16458
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20548 14890 20576 15030
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20548 12442 20576 13942
rect 20640 13569 20668 16730
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15638 20852 15846
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20810 15192 20866 15201
rect 20916 15162 20944 15506
rect 20810 15127 20866 15136
rect 20904 15156 20956 15162
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14278 20760 14758
rect 20824 14618 20852 15127
rect 20904 15098 20956 15104
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 21008 14498 21036 18702
rect 21100 17814 21128 19246
rect 21560 19242 21588 20810
rect 21928 20602 21956 21422
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22112 19310 22140 19790
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21284 18290 21312 19110
rect 21376 18834 21404 19110
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 21468 17610 21496 18566
rect 21652 18426 21680 19246
rect 21824 18760 21876 18766
rect 21822 18728 21824 18737
rect 21876 18728 21878 18737
rect 21822 18663 21878 18672
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 22204 18358 22232 20266
rect 22296 19990 22324 20878
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20534 22784 20742
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22296 19786 22324 19926
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22296 18766 22324 19722
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17134 22140 17478
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21100 14929 21128 16934
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15745 21312 15846
rect 21270 15736 21326 15745
rect 21270 15671 21326 15680
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21086 14920 21142 14929
rect 21086 14855 21142 14864
rect 21284 14618 21312 15370
rect 21560 14618 21588 16594
rect 21822 16144 21878 16153
rect 21822 16079 21824 16088
rect 21876 16079 21878 16088
rect 21824 16050 21876 16056
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21376 14498 21404 14554
rect 20824 14470 21036 14498
rect 21284 14470 21404 14498
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20626 13560 20682 13569
rect 20626 13495 20682 13504
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20732 12782 20760 13398
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20732 11830 20760 12718
rect 20824 12594 20852 14470
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21100 13394 21128 14282
rect 21192 13938 21220 14350
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 21192 13297 21220 13874
rect 21178 13288 21234 13297
rect 21178 13223 21234 13232
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20902 12608 20958 12617
rect 20824 12566 20902 12594
rect 20902 12543 20958 12552
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20456 11354 20484 11766
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20352 11008 20404 11014
rect 20352 10950 20404 10956
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20258 10296 20314 10305
rect 20258 10231 20314 10240
rect 20272 10198 20300 10231
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20180 9674 20208 9998
rect 20180 9646 20300 9674
rect 20364 9654 20392 10950
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8673 20024 8910
rect 19982 8664 20038 8673
rect 19982 8599 20038 8608
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 8022 19472 8366
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19260 5574 19288 6190
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 19260 2310 19288 5510
rect 19444 4214 19472 6870
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19628 4593 19656 4626
rect 19614 4584 19670 4593
rect 19614 4519 19670 4528
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19340 3528 19392 3534
rect 19338 3496 19340 3505
rect 19392 3496 19394 3505
rect 19338 3431 19394 3440
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19352 800 19380 3334
rect 19444 2990 19472 4150
rect 19996 3670 20024 8599
rect 20180 7834 20208 9522
rect 20272 8974 20300 9646
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8498 20300 8910
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20088 7806 20208 7834
rect 20088 4690 20116 7806
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 7546 20208 7686
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20272 6458 20300 8298
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20364 5778 20392 9318
rect 20456 9042 20484 10542
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20548 10062 20576 10406
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20456 4457 20484 8842
rect 20548 8430 20576 9998
rect 20640 8634 20668 11154
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 9994 20760 11018
rect 20824 9994 20852 11494
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20536 8424 20588 8430
rect 20588 8372 20668 8378
rect 20536 8366 20668 8372
rect 20548 8350 20668 8366
rect 20640 7954 20668 8350
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20640 7342 20668 7890
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 6390 20668 7278
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20732 4826 20760 9318
rect 20824 6882 20852 9930
rect 20916 9042 20944 12543
rect 21008 11898 21036 13126
rect 21192 12850 21220 13223
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21178 12472 21234 12481
rect 21284 12458 21312 14470
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21744 13394 21772 13806
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12986 21404 13126
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21468 12782 21496 13330
rect 21744 12918 21772 13330
rect 21732 12912 21784 12918
rect 21732 12854 21784 12860
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21234 12430 21312 12458
rect 21836 12442 21864 16050
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 22204 14498 22232 14826
rect 22112 14470 22232 14498
rect 22112 14278 22140 14470
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21928 13512 21956 14214
rect 22020 14074 22048 14214
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22296 13954 22324 18702
rect 22388 17746 22416 20470
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 18834 22600 19110
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22388 17542 22416 17682
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22388 16250 22416 17478
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22480 16096 22508 18022
rect 22388 16068 22508 16096
rect 22388 15434 22416 16068
rect 22664 16046 22692 18022
rect 22756 16522 22784 18566
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 22848 17134 22876 17750
rect 22940 17746 22968 19722
rect 23308 19310 23336 20334
rect 23400 19786 23428 20470
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23492 19718 23520 21286
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23584 19310 23612 21898
rect 23756 21412 23808 21418
rect 23756 21354 23808 21360
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22848 16522 22876 17070
rect 22940 16726 22968 17682
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22468 15972 22520 15978
rect 22468 15914 22520 15920
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22480 15162 22508 15914
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22388 14346 22416 14894
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22572 14074 22600 15030
rect 22664 14074 22692 15030
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22650 13968 22706 13977
rect 22100 13932 22152 13938
rect 22296 13926 22600 13954
rect 22100 13874 22152 13880
rect 22112 13841 22140 13874
rect 22098 13832 22154 13841
rect 22098 13767 22154 13776
rect 22008 13524 22060 13530
rect 21928 13484 22008 13512
rect 22008 13466 22060 13472
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 21824 12436 21876 12442
rect 21178 12407 21234 12416
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20916 7002 20944 7754
rect 21008 7274 21036 10950
rect 21086 10568 21142 10577
rect 21086 10503 21088 10512
rect 21140 10503 21142 10512
rect 21088 10474 21140 10480
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 20996 7268 21048 7274
rect 20996 7210 21048 7216
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20824 6854 20944 6882
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20442 4448 20498 4457
rect 20442 4383 20498 4392
rect 20732 4010 20760 4626
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 19800 3664 19852 3670
rect 19800 3606 19852 3612
rect 19984 3664 20036 3670
rect 19984 3606 20036 3612
rect 19812 3448 19840 3606
rect 19812 3420 20208 3448
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 20180 2854 20208 3420
rect 20824 3126 20852 6598
rect 20916 4078 20944 6854
rect 21100 5642 21128 9862
rect 21192 8566 21220 12407
rect 21824 12378 21876 12384
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 12102 21312 12174
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 22296 11898 22324 13194
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22376 12776 22428 12782
rect 22480 12753 22508 13126
rect 22376 12718 22428 12724
rect 22466 12744 22522 12753
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21284 10674 21312 10746
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21376 10470 21404 10746
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21180 8560 21232 8566
rect 21180 8502 21232 8508
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 20994 4584 21050 4593
rect 20994 4519 21050 4528
rect 21008 4146 21036 4519
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 21100 3369 21128 3538
rect 21086 3360 21142 3369
rect 21086 3295 21142 3304
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 21192 2446 21220 8026
rect 21284 7410 21312 8298
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 5574 21312 6258
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21100 2038 21128 2314
rect 21088 2032 21140 2038
rect 21088 1974 21140 1980
rect 21284 800 21312 5510
rect 21376 3194 21404 10406
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21468 9926 21496 10202
rect 21560 10130 21588 10950
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21468 7206 21496 9522
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21468 5710 21496 6598
rect 21560 5846 21588 8570
rect 21652 8537 21680 11222
rect 21822 10296 21878 10305
rect 21822 10231 21824 10240
rect 21876 10231 21878 10240
rect 21824 10202 21876 10208
rect 21928 10198 21956 11698
rect 22008 10736 22060 10742
rect 22008 10678 22060 10684
rect 21916 10192 21968 10198
rect 21836 10140 21916 10146
rect 21836 10134 21968 10140
rect 21836 10118 21956 10134
rect 21836 8634 21864 10118
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21638 8528 21694 8537
rect 21638 8463 21694 8472
rect 21822 8528 21878 8537
rect 21822 8463 21824 8472
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21652 5166 21680 8463
rect 21876 8463 21878 8472
rect 21824 8434 21876 8440
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21836 7478 21864 7754
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21744 5302 21772 5510
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21468 3466 21496 4966
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 4146 21588 4422
rect 21836 4214 21864 6938
rect 21928 6934 21956 9998
rect 22020 7834 22048 10678
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 9761 22140 10406
rect 22098 9752 22154 9761
rect 22098 9687 22154 9696
rect 22388 9178 22416 12718
rect 22466 12679 22522 12688
rect 22572 11830 22600 13926
rect 22650 13903 22652 13912
rect 22704 13903 22706 13912
rect 22652 13874 22704 13880
rect 22664 13705 22692 13874
rect 22650 13696 22706 13705
rect 22650 13631 22706 13640
rect 22848 13462 22876 15370
rect 22928 14816 22980 14822
rect 22926 14784 22928 14793
rect 22980 14784 22982 14793
rect 22926 14719 22982 14728
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22940 13258 22968 13466
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 12306 22876 12582
rect 23032 12442 23060 17546
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23308 16046 23336 16934
rect 23492 16522 23520 17070
rect 23584 17066 23612 19246
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 23572 17060 23624 17066
rect 23572 17002 23624 17008
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22756 11234 22784 11834
rect 22480 11206 22784 11234
rect 22480 11150 22508 11206
rect 22756 11150 22784 11206
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22112 8129 22140 8842
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22388 8430 22416 8774
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22284 8356 22336 8362
rect 22284 8298 22336 8304
rect 22098 8120 22154 8129
rect 22098 8055 22154 8064
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22020 7806 22140 7834
rect 22112 7290 22140 7806
rect 22204 7750 22232 7890
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22112 7274 22232 7290
rect 22112 7268 22244 7274
rect 22112 7262 22192 7268
rect 22192 7210 22244 7216
rect 22296 7154 22324 8298
rect 22204 7126 22324 7154
rect 21916 6928 21968 6934
rect 21916 6870 21968 6876
rect 22006 6896 22062 6905
rect 22006 6831 22062 6840
rect 22100 6860 22152 6866
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21928 5234 21956 6666
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21914 4312 21970 4321
rect 21914 4247 21916 4256
rect 21968 4247 21970 4256
rect 21916 4218 21968 4224
rect 21824 4208 21876 4214
rect 21824 4150 21876 4156
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21836 3534 21864 3946
rect 22020 3584 22048 6831
rect 22100 6802 22152 6808
rect 22112 6458 22140 6802
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22112 4622 22140 6394
rect 22204 5914 22232 7126
rect 22284 6384 22336 6390
rect 22284 6326 22336 6332
rect 22296 6254 22324 6326
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22112 4298 22140 4558
rect 22112 4282 22508 4298
rect 22112 4276 22520 4282
rect 22112 4270 22468 4276
rect 22112 3602 22140 4270
rect 22468 4218 22520 4224
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22204 3602 22232 3674
rect 22466 3632 22522 3641
rect 21928 3556 22048 3584
rect 22100 3596 22152 3602
rect 21824 3528 21876 3534
rect 21730 3496 21786 3505
rect 21456 3460 21508 3466
rect 21824 3470 21876 3476
rect 21730 3431 21786 3440
rect 21456 3402 21508 3408
rect 21744 3398 21772 3431
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21468 2854 21496 3130
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21928 2514 21956 3556
rect 22100 3538 22152 3544
rect 22192 3596 22244 3602
rect 22466 3567 22522 3576
rect 22192 3538 22244 3544
rect 22112 2514 22140 3538
rect 22480 3466 22508 3567
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22204 3097 22232 3130
rect 22468 3120 22520 3126
rect 22190 3088 22246 3097
rect 22190 3023 22246 3032
rect 22466 3088 22468 3097
rect 22520 3088 22522 3097
rect 22466 3023 22522 3032
rect 21916 2508 21968 2514
rect 21916 2450 21968 2456
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 21928 1970 21956 2450
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 22572 800 22600 3674
rect 22664 2922 22692 11086
rect 22756 10742 22784 11086
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22756 10198 22784 10678
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22742 8664 22798 8673
rect 22742 8599 22798 8608
rect 22756 8566 22784 8599
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22848 8362 22876 12242
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22940 12073 22968 12106
rect 22926 12064 22982 12073
rect 22926 11999 22982 12008
rect 23124 11914 23152 15846
rect 23308 15706 23336 15982
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23308 14958 23336 15642
rect 23492 15434 23520 15982
rect 23584 15706 23612 16118
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23216 14482 23244 14826
rect 23676 14482 23704 18294
rect 23768 18222 23796 21354
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23952 15722 23980 22066
rect 24032 18692 24084 18698
rect 24032 18634 24084 18640
rect 24044 18426 24072 18634
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24136 18358 24164 30194
rect 24412 23866 24440 34478
rect 24596 29850 24624 37198
rect 27344 37188 27396 37194
rect 27344 37130 27396 37136
rect 27356 36922 27384 37130
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27448 36553 27476 37198
rect 27724 37126 27752 39200
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 28356 36780 28408 36786
rect 28356 36722 28408 36728
rect 27434 36544 27490 36553
rect 27434 36479 27490 36488
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 25596 29504 25648 29510
rect 25596 29446 25648 29452
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 23952 15694 24072 15722
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23400 14198 23612 14226
rect 23400 14074 23428 14198
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23584 14006 23612 14198
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23664 13864 23716 13870
rect 23768 13841 23796 15574
rect 23940 14952 23992 14958
rect 23938 14920 23940 14929
rect 23992 14920 23994 14929
rect 23938 14855 23994 14864
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23860 14414 23888 14554
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23664 13806 23716 13812
rect 23754 13832 23810 13841
rect 23572 13456 23624 13462
rect 23572 13398 23624 13404
rect 23584 13274 23612 13398
rect 23492 13246 23612 13274
rect 23492 12850 23520 13246
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23676 12782 23704 13806
rect 23754 13767 23810 13776
rect 23768 13326 23796 13767
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 24044 12850 24072 15694
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23388 12708 23440 12714
rect 23440 12668 23520 12696
rect 23388 12650 23440 12656
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23124 11886 23244 11914
rect 23400 11898 23428 12174
rect 23112 11824 23164 11830
rect 23032 11772 23112 11778
rect 23032 11766 23164 11772
rect 23032 11750 23152 11766
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22940 10674 22968 11630
rect 23032 11393 23060 11750
rect 23216 11506 23244 11886
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23124 11478 23244 11506
rect 23018 11384 23074 11393
rect 23018 11319 23074 11328
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 22940 9042 22968 10610
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22940 8498 22968 8978
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 23032 8378 23060 11319
rect 23124 10742 23152 11478
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23124 8401 23152 8910
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 22940 8350 23060 8378
rect 23110 8392 23166 8401
rect 22742 7576 22798 7585
rect 22742 7511 22798 7520
rect 22756 7478 22784 7511
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22756 7342 22784 7414
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22940 6118 22968 8350
rect 23110 8327 23166 8336
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23124 6610 23152 8327
rect 23216 6798 23244 11290
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23204 6656 23256 6662
rect 23124 6604 23204 6610
rect 23124 6598 23256 6604
rect 23032 6254 23060 6598
rect 23124 6582 23244 6598
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 23216 6202 23244 6582
rect 23308 6390 23336 11222
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23400 10033 23428 10406
rect 23386 10024 23442 10033
rect 23386 9959 23442 9968
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23400 7546 23428 8026
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23492 6338 23520 12668
rect 23768 12434 23796 12786
rect 23768 12406 23888 12434
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23676 11218 23704 12038
rect 23768 11801 23796 12038
rect 23754 11792 23810 11801
rect 23754 11727 23810 11736
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23584 7206 23612 11018
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23676 8430 23704 10678
rect 23768 10452 23796 11727
rect 23860 10554 23888 12406
rect 24044 12102 24072 12786
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 23860 10526 24072 10554
rect 23768 10424 23980 10452
rect 23952 10198 23980 10424
rect 23940 10192 23992 10198
rect 23940 10134 23992 10140
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23676 7342 23704 7890
rect 23768 7818 23796 9862
rect 23848 9512 23900 9518
rect 23846 9480 23848 9489
rect 23900 9480 23902 9489
rect 23846 9415 23902 9424
rect 23952 8106 23980 10134
rect 24044 9926 24072 10526
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9382 24072 9862
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24044 8906 24072 9318
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 23860 8078 23980 8106
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23754 6760 23810 6769
rect 23754 6695 23810 6704
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23676 6458 23704 6598
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23492 6310 23704 6338
rect 23216 6174 23336 6202
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23204 5296 23256 5302
rect 23124 5244 23204 5250
rect 23124 5238 23256 5244
rect 23124 5222 23244 5238
rect 23124 5030 23152 5222
rect 23112 5024 23164 5030
rect 22834 4992 22890 5001
rect 23112 4966 23164 4972
rect 22834 4927 22890 4936
rect 22848 4554 22876 4927
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 23308 3913 23336 6174
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23400 5030 23428 5646
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23400 4282 23428 4966
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23492 4214 23520 6054
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23676 5522 23704 6310
rect 23768 5710 23796 6695
rect 23860 6458 23888 8078
rect 24136 7426 24164 18158
rect 24228 16726 24256 18158
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24320 17134 24348 17478
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24216 16720 24268 16726
rect 24216 16662 24268 16668
rect 24308 16176 24360 16182
rect 24360 16124 24440 16130
rect 24308 16118 24440 16124
rect 24320 16102 24440 16118
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24320 15910 24348 15982
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24320 15094 24348 15846
rect 24412 15502 24440 16102
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24214 12880 24270 12889
rect 24214 12815 24216 12824
rect 24268 12815 24270 12824
rect 24216 12786 24268 12792
rect 24412 12434 24440 15438
rect 24504 13705 24532 29446
rect 25504 27328 25556 27334
rect 25504 27270 25556 27276
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 22094 24900 23462
rect 24872 22066 25084 22094
rect 24952 20936 25004 20942
rect 24950 20904 24952 20913
rect 25004 20904 25006 20913
rect 24950 20839 25006 20848
rect 24584 19780 24636 19786
rect 24584 19722 24636 19728
rect 24596 19310 24624 19722
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 24596 16726 24624 17002
rect 24584 16720 24636 16726
rect 24584 16662 24636 16668
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24596 14958 24624 15506
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24688 15162 24716 15302
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24490 13696 24546 13705
rect 24490 13631 24546 13640
rect 24504 13326 24532 13631
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24780 12753 24808 18226
rect 24872 17338 24900 18634
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24964 17270 24992 18566
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 25056 17134 25084 22066
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25240 19922 25268 20742
rect 25332 20466 25360 21286
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25332 18154 25360 20402
rect 25516 19446 25544 27270
rect 25608 22094 25636 29446
rect 26620 24818 26648 35022
rect 27172 32910 27200 35634
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 27172 26586 27200 32846
rect 27160 26580 27212 26586
rect 27160 26522 27212 26528
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26620 24614 26648 24754
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26620 22642 26648 24550
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 25608 22066 25820 22094
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25516 18222 25544 19382
rect 25596 19236 25648 19242
rect 25596 19178 25648 19184
rect 25608 18970 25636 19178
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18358 25636 18566
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25320 18148 25372 18154
rect 25320 18090 25372 18096
rect 25332 17762 25360 18090
rect 25332 17734 25452 17762
rect 25792 17746 25820 22066
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25884 20466 25912 20742
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 25884 20058 25912 20402
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25872 20052 25924 20058
rect 25872 19994 25924 20000
rect 25976 19786 26004 20198
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 25872 19168 25924 19174
rect 25872 19110 25924 19116
rect 25884 18698 25912 19110
rect 25964 18964 26016 18970
rect 25964 18906 26016 18912
rect 25872 18692 25924 18698
rect 25872 18634 25924 18640
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 25228 17060 25280 17066
rect 25228 17002 25280 17008
rect 25044 16516 25096 16522
rect 25044 16458 25096 16464
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24872 13530 24900 15302
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24766 12744 24822 12753
rect 24584 12708 24636 12714
rect 24766 12679 24822 12688
rect 24584 12650 24636 12656
rect 24320 12406 24440 12434
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24228 10062 24256 10950
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 24228 8566 24256 9318
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24320 8022 24348 12406
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24504 9042 24532 9522
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 23952 7398 24164 7426
rect 24216 7472 24268 7478
rect 24320 7460 24348 7958
rect 24268 7432 24348 7460
rect 24216 7414 24268 7420
rect 23952 7342 23980 7398
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 23952 6730 23980 7278
rect 23940 6724 23992 6730
rect 23940 6666 23992 6672
rect 23952 6633 23980 6666
rect 23938 6624 23994 6633
rect 23938 6559 23994 6568
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23860 5778 23888 6394
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23388 3936 23440 3942
rect 23294 3904 23350 3913
rect 23388 3878 23440 3884
rect 23294 3839 23350 3848
rect 23400 3777 23428 3878
rect 23386 3768 23442 3777
rect 23584 3738 23612 5510
rect 23676 5494 23888 5522
rect 23860 4078 23888 5494
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23386 3703 23442 3712
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 24044 2854 24072 7278
rect 24412 6866 24440 8298
rect 24504 7954 24532 8978
rect 24492 7948 24544 7954
rect 24492 7890 24544 7896
rect 24504 6866 24532 7890
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24596 6338 24624 12650
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24780 12170 24808 12378
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24674 11112 24730 11121
rect 24674 11047 24676 11056
rect 24728 11047 24730 11056
rect 24676 11018 24728 11024
rect 24872 10713 24900 13330
rect 24964 11370 24992 13738
rect 25056 11898 25084 16458
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25148 12646 25176 15370
rect 25240 14074 25268 17002
rect 25424 16522 25452 17734
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25608 17270 25636 17546
rect 25596 17264 25648 17270
rect 25596 17206 25648 17212
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 25596 17060 25648 17066
rect 25596 17002 25648 17008
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 16182 25452 16458
rect 25608 16454 25636 17002
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 25504 15632 25556 15638
rect 25504 15574 25556 15580
rect 25412 15428 25464 15434
rect 25412 15370 25464 15376
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25332 13530 25360 14214
rect 25424 13870 25452 15370
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25332 12434 25360 12582
rect 25148 12406 25360 12434
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25044 11552 25096 11558
rect 25148 11506 25176 12406
rect 25424 12322 25452 12786
rect 25332 12294 25452 12322
rect 25332 11937 25360 12294
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25318 11928 25374 11937
rect 25318 11863 25374 11872
rect 25228 11756 25280 11762
rect 25424 11744 25452 12174
rect 25280 11716 25452 11744
rect 25228 11698 25280 11704
rect 25318 11656 25374 11665
rect 25318 11591 25374 11600
rect 25096 11500 25176 11506
rect 25044 11494 25176 11500
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25056 11478 25176 11494
rect 24964 11342 25084 11370
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24964 10810 24992 10950
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24858 10704 24914 10713
rect 24858 10639 24914 10648
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24688 9602 24716 9998
rect 24780 9926 24808 10406
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24872 9994 24900 10134
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24688 9574 24808 9602
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24688 8294 24716 8570
rect 24780 8378 24808 9574
rect 24780 8350 24900 8378
rect 24872 8294 24900 8350
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24860 8288 24912 8294
rect 24860 8230 24912 8236
rect 24872 7954 24900 8230
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24596 6310 24716 6338
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24596 5778 24624 6190
rect 24688 5817 24716 6310
rect 24674 5808 24730 5817
rect 24584 5772 24636 5778
rect 24674 5743 24730 5752
rect 24584 5714 24636 5720
rect 24398 5400 24454 5409
rect 24398 5335 24454 5344
rect 24308 5024 24360 5030
rect 24308 4966 24360 4972
rect 24320 4826 24348 4966
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24306 4720 24362 4729
rect 24306 4655 24308 4664
rect 24360 4655 24362 4664
rect 24308 4626 24360 4632
rect 24122 4584 24178 4593
rect 24122 4519 24178 4528
rect 24136 4486 24164 4519
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 24412 3466 24440 5335
rect 24596 5234 24624 5714
rect 24780 5642 24808 6802
rect 24964 6390 24992 7686
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 24596 4690 24624 5170
rect 24872 4690 24900 5850
rect 24584 4684 24636 4690
rect 24584 4626 24636 4632
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 24596 3738 24624 4626
rect 24858 4584 24914 4593
rect 24858 4519 24914 4528
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24596 3602 24624 3674
rect 24872 3602 24900 4519
rect 25056 4078 25084 11342
rect 25148 5817 25176 11478
rect 25240 10169 25268 11494
rect 25226 10160 25282 10169
rect 25226 10095 25282 10104
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25240 9178 25268 9590
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25332 9058 25360 11591
rect 25516 10810 25544 15574
rect 25608 14346 25636 16390
rect 25700 14958 25728 17070
rect 25792 16658 25820 17682
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25792 16046 25820 16594
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 25872 16040 25924 16046
rect 25872 15982 25924 15988
rect 25884 15638 25912 15982
rect 25976 15638 26004 18906
rect 26620 18834 26648 22374
rect 27436 20528 27488 20534
rect 27436 20470 27488 20476
rect 27160 20324 27212 20330
rect 27160 20266 27212 20272
rect 27172 19786 27200 20266
rect 27068 19780 27120 19786
rect 27068 19722 27120 19728
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27080 19514 27108 19722
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 27080 18970 27108 19246
rect 27068 18964 27120 18970
rect 27068 18906 27120 18912
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26620 17542 26648 18770
rect 26700 18760 26752 18766
rect 26698 18728 26700 18737
rect 26752 18728 26754 18737
rect 26698 18663 26754 18672
rect 26712 18426 26740 18663
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 27080 18086 27108 18906
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26620 16726 26648 17138
rect 26976 16992 27028 16998
rect 26976 16934 27028 16940
rect 26608 16720 26660 16726
rect 26608 16662 26660 16668
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 25780 15088 25832 15094
rect 25780 15030 25832 15036
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25792 14618 25820 15030
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 25780 14612 25832 14618
rect 25780 14554 25832 14560
rect 26240 14544 26292 14550
rect 26240 14486 26292 14492
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 26252 14249 26280 14486
rect 26238 14240 26294 14249
rect 26238 14175 26294 14184
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 25976 13462 26004 13806
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 25688 13320 25740 13326
rect 25740 13280 25820 13308
rect 25688 13262 25740 13268
rect 25594 12472 25650 12481
rect 25594 12407 25650 12416
rect 25608 12322 25636 12407
rect 25608 12294 25728 12322
rect 25700 12238 25728 12294
rect 25792 12288 25820 13280
rect 25976 12782 26004 13398
rect 26252 13258 26280 13670
rect 26344 13326 26372 14894
rect 26436 14890 26464 16594
rect 26620 16266 26648 16662
rect 26988 16522 27016 16934
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 27068 16516 27120 16522
rect 27068 16458 27120 16464
rect 26528 16238 26648 16266
rect 26528 15201 26556 16238
rect 26608 16176 26660 16182
rect 26608 16118 26660 16124
rect 26514 15192 26570 15201
rect 26514 15127 26570 15136
rect 26424 14884 26476 14890
rect 26424 14826 26476 14832
rect 26528 14113 26556 15127
rect 26514 14104 26570 14113
rect 26514 14039 26570 14048
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26056 12912 26108 12918
rect 26056 12854 26108 12860
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25792 12260 26004 12288
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25778 12200 25834 12209
rect 25596 12164 25648 12170
rect 25778 12135 25780 12144
rect 25596 12106 25648 12112
rect 25832 12135 25834 12144
rect 25780 12106 25832 12112
rect 25608 11558 25636 12106
rect 25870 11928 25926 11937
rect 25870 11863 25926 11872
rect 25688 11756 25740 11762
rect 25740 11716 25820 11744
rect 25688 11698 25740 11704
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 10736 25464 10742
rect 25412 10678 25464 10684
rect 25424 9654 25452 10678
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25240 9030 25360 9058
rect 25516 9042 25544 10746
rect 25504 9036 25556 9042
rect 25134 5808 25190 5817
rect 25134 5743 25190 5752
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 25240 3890 25268 9030
rect 25504 8978 25556 8984
rect 25608 7478 25636 11290
rect 25792 11150 25820 11716
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25700 9654 25728 10202
rect 25792 9761 25820 11086
rect 25778 9752 25834 9761
rect 25778 9687 25834 9696
rect 25688 9648 25740 9654
rect 25686 9616 25688 9625
rect 25740 9616 25742 9625
rect 25792 9586 25820 9687
rect 25686 9551 25742 9560
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25884 8537 25912 11863
rect 25870 8528 25926 8537
rect 25870 8463 25926 8472
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25596 7472 25648 7478
rect 25596 7414 25648 7420
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25516 5642 25544 7346
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 25056 3862 25268 3890
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24320 2990 24348 3334
rect 24492 3052 24544 3058
rect 24596 3040 24624 3538
rect 25056 3505 25084 3862
rect 25228 3596 25280 3602
rect 25148 3556 25228 3584
rect 25042 3496 25098 3505
rect 25148 3466 25176 3556
rect 25228 3538 25280 3544
rect 25042 3431 25098 3440
rect 25136 3460 25188 3466
rect 25136 3402 25188 3408
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24544 3012 24624 3040
rect 24492 2994 24544 3000
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24032 2848 24084 2854
rect 24412 2825 24440 2926
rect 24032 2790 24084 2796
rect 24398 2816 24454 2825
rect 24398 2751 24454 2760
rect 24674 2816 24730 2825
rect 24674 2751 24730 2760
rect 24688 2106 24716 2751
rect 24676 2100 24728 2106
rect 24676 2042 24728 2048
rect 24504 870 24624 898
rect 24504 800 24532 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 7746 200 7802 800
rect 9678 200 9734 800
rect 10966 200 11022 800
rect 12898 200 12954 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 24490 200 24546 800
rect 24596 762 24624 870
rect 24780 762 24808 3334
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24872 2990 24900 3062
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 25700 2774 25728 8298
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25884 5302 25912 7890
rect 25976 5914 26004 12260
rect 26068 10810 26096 12854
rect 26148 12708 26200 12714
rect 26148 12650 26200 12656
rect 26160 12306 26188 12650
rect 26252 12434 26280 13194
rect 26332 12776 26384 12782
rect 26330 12744 26332 12753
rect 26384 12744 26386 12753
rect 26330 12679 26386 12688
rect 26252 12406 26372 12434
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26148 12164 26200 12170
rect 26148 12106 26200 12112
rect 26160 11014 26188 12106
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 26056 10804 26108 10810
rect 26056 10746 26108 10752
rect 26252 9466 26280 11698
rect 26160 9438 26280 9466
rect 26056 9104 26108 9110
rect 26056 9046 26108 9052
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 25962 5808 26018 5817
rect 25962 5743 26018 5752
rect 25976 5642 26004 5743
rect 25964 5636 26016 5642
rect 25964 5578 26016 5584
rect 25872 5296 25924 5302
rect 25872 5238 25924 5244
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 25976 4729 26004 4966
rect 25962 4720 26018 4729
rect 25962 4655 26018 4664
rect 25962 4448 26018 4457
rect 25962 4383 26018 4392
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 25884 3602 25912 3946
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 25608 2746 25728 2774
rect 25608 2038 25636 2746
rect 25976 2514 26004 4383
rect 26068 4214 26096 9046
rect 26160 9042 26188 9438
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 26252 8974 26280 9318
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 26160 7750 26188 7822
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26252 6905 26280 8366
rect 26238 6896 26294 6905
rect 26238 6831 26294 6840
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26252 5914 26280 6394
rect 26240 5908 26292 5914
rect 26240 5850 26292 5856
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26252 5001 26280 5170
rect 26238 4992 26294 5001
rect 26238 4927 26294 4936
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 26056 4208 26108 4214
rect 26056 4150 26108 4156
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 26068 2378 26096 4014
rect 26252 3398 26280 4490
rect 26344 4146 26372 12406
rect 26436 11898 26464 13942
rect 26516 13728 26568 13734
rect 26514 13696 26516 13705
rect 26568 13696 26570 13705
rect 26514 13631 26570 13640
rect 26620 12238 26648 16118
rect 27080 15910 27108 16458
rect 27068 15904 27120 15910
rect 27068 15846 27120 15852
rect 26884 15156 26936 15162
rect 26884 15098 26936 15104
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26804 14618 26832 14758
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26790 14104 26846 14113
rect 26790 14039 26846 14048
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26712 10849 26740 11086
rect 26698 10840 26754 10849
rect 26698 10775 26754 10784
rect 26712 10742 26740 10775
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26436 8430 26464 10610
rect 26700 10532 26752 10538
rect 26700 10474 26752 10480
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26620 9518 26648 9998
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 26528 8566 26556 9386
rect 26620 9042 26648 9454
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26620 8634 26648 8842
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26528 7750 26556 8502
rect 26712 8294 26740 10474
rect 26804 9489 26832 14039
rect 26896 14006 26924 15098
rect 27068 14476 27120 14482
rect 26988 14436 27068 14464
rect 26988 14346 27016 14436
rect 27068 14418 27120 14424
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 26884 10668 26936 10674
rect 26884 10610 26936 10616
rect 26790 9480 26846 9489
rect 26790 9415 26846 9424
rect 26700 8288 26752 8294
rect 26700 8230 26752 8236
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26712 7478 26740 7686
rect 26700 7472 26752 7478
rect 26700 7414 26752 7420
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26332 4140 26384 4146
rect 26332 4082 26384 4088
rect 26436 3942 26464 5306
rect 26620 4690 26648 6734
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26712 6633 26740 6666
rect 26698 6624 26754 6633
rect 26698 6559 26754 6568
rect 26804 5166 26832 9415
rect 26896 5302 26924 10610
rect 26988 8906 27016 13874
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 27080 12850 27108 13126
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27080 12714 27108 12786
rect 27068 12708 27120 12714
rect 27068 12650 27120 12656
rect 27066 12336 27122 12345
rect 27066 12271 27068 12280
rect 27120 12271 27122 12280
rect 27068 12242 27120 12248
rect 27172 10538 27200 18702
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27264 16250 27292 18022
rect 27356 17814 27384 18226
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27342 16144 27398 16153
rect 27342 16079 27344 16088
rect 27396 16079 27398 16088
rect 27344 16050 27396 16056
rect 27356 15910 27384 16050
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27448 15178 27476 20470
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27632 18222 27660 19654
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27632 17626 27660 18158
rect 27724 17746 27752 18566
rect 28368 17882 28396 36722
rect 28460 35834 28488 37198
rect 29656 37126 29684 39200
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 28448 35828 28500 35834
rect 28448 35770 28500 35776
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 29840 31142 29868 31282
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 29736 29572 29788 29578
rect 29736 29514 29788 29520
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28828 18086 28856 18362
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28356 17876 28408 17882
rect 28356 17818 28408 17824
rect 27896 17808 27948 17814
rect 27896 17750 27948 17756
rect 27712 17740 27764 17746
rect 27712 17682 27764 17688
rect 27632 17610 27752 17626
rect 27528 17604 27580 17610
rect 27632 17604 27764 17610
rect 27632 17598 27712 17604
rect 27528 17546 27580 17552
rect 27712 17546 27764 17552
rect 27540 17354 27568 17546
rect 27540 17338 27660 17354
rect 27540 17332 27672 17338
rect 27540 17326 27620 17332
rect 27620 17274 27672 17280
rect 27908 16250 27936 17750
rect 28828 17202 28856 18022
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17202 29040 17478
rect 28816 17196 28868 17202
rect 28816 17138 28868 17144
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 28632 17128 28684 17134
rect 28632 17070 28684 17076
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28184 16250 28212 16458
rect 27896 16244 27948 16250
rect 27896 16186 27948 16192
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 27528 15972 27580 15978
rect 27528 15914 27580 15920
rect 27540 15434 27568 15914
rect 27908 15570 27936 16186
rect 28080 15632 28132 15638
rect 28080 15574 28132 15580
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27448 15150 27752 15178
rect 27620 15088 27672 15094
rect 27620 15030 27672 15036
rect 27344 14952 27396 14958
rect 27250 14920 27306 14929
rect 27396 14900 27568 14906
rect 27344 14894 27568 14900
rect 27356 14878 27568 14894
rect 27250 14855 27306 14864
rect 27264 14346 27292 14855
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27540 13394 27568 14878
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27448 12986 27476 13330
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27448 12646 27476 12786
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27344 12096 27396 12102
rect 27250 12064 27306 12073
rect 27396 12056 27568 12084
rect 27344 12038 27396 12044
rect 27250 11999 27306 12008
rect 27264 11898 27292 11999
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 27540 11762 27568 12056
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27356 11665 27384 11698
rect 27342 11656 27398 11665
rect 27342 11591 27398 11600
rect 27356 11286 27384 11591
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 10606 27292 10950
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27068 10056 27120 10062
rect 27068 9998 27120 10004
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 26988 6118 27016 8842
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 27080 5370 27108 9998
rect 27356 9761 27384 11086
rect 27632 10266 27660 15030
rect 27724 14958 27752 15150
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 27712 13252 27764 13258
rect 27712 13194 27764 13200
rect 27724 12481 27752 13194
rect 27710 12472 27766 12481
rect 27710 12407 27766 12416
rect 27816 11898 27844 15370
rect 28092 14414 28120 15574
rect 28276 15502 28304 16594
rect 28356 16448 28408 16454
rect 28356 16390 28408 16396
rect 28368 16114 28396 16390
rect 28644 16114 28672 17070
rect 28724 16992 28776 16998
rect 28724 16934 28776 16940
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28632 15564 28684 15570
rect 28632 15506 28684 15512
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28172 14816 28224 14822
rect 28170 14784 28172 14793
rect 28224 14784 28226 14793
rect 28170 14719 28226 14728
rect 28276 14618 28304 15438
rect 28540 15428 28592 15434
rect 28540 15370 28592 15376
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 27896 14000 27948 14006
rect 27896 13942 27948 13948
rect 27804 11892 27856 11898
rect 27804 11834 27856 11840
rect 27908 11354 27936 13942
rect 28092 13870 28120 14350
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28092 13394 28120 13806
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27988 13252 28040 13258
rect 27988 13194 28040 13200
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 28000 10810 28028 13194
rect 28078 12472 28134 12481
rect 28078 12407 28134 12416
rect 27988 10804 28040 10810
rect 27988 10746 28040 10752
rect 28092 10742 28120 12407
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 28080 10736 28132 10742
rect 28080 10678 28132 10684
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 27342 9752 27398 9761
rect 27342 9687 27398 9696
rect 27356 9586 27384 9687
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27160 9444 27212 9450
rect 27160 9386 27212 9392
rect 27172 7818 27200 9386
rect 27356 8498 27384 9522
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27160 7812 27212 7818
rect 27160 7754 27212 7760
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27264 7002 27292 7142
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 27252 6656 27304 6662
rect 27252 6598 27304 6604
rect 27264 6118 27292 6598
rect 27540 6254 27568 7142
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27068 5364 27120 5370
rect 27068 5306 27120 5312
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 26792 5160 26844 5166
rect 26792 5102 26844 5108
rect 26698 4856 26754 4865
rect 26698 4791 26754 4800
rect 26712 4690 26740 4791
rect 26608 4684 26660 4690
rect 26608 4626 26660 4632
rect 26700 4684 26752 4690
rect 26700 4626 26752 4632
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26528 4282 26556 4558
rect 26606 4312 26662 4321
rect 26516 4276 26568 4282
rect 26606 4247 26608 4256
rect 26516 4218 26568 4224
rect 26660 4247 26662 4256
rect 26608 4218 26660 4224
rect 26896 4078 26924 5238
rect 27264 5166 27292 6054
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 27252 5160 27304 5166
rect 27252 5102 27304 5108
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26988 4593 27016 4626
rect 26974 4584 27030 4593
rect 27356 4554 27384 5510
rect 27632 4622 27660 9930
rect 27712 9920 27764 9926
rect 27712 9862 27764 9868
rect 27724 8634 27752 9862
rect 27802 9616 27858 9625
rect 27802 9551 27804 9560
rect 27856 9551 27858 9560
rect 27804 9522 27856 9528
rect 27908 9518 27936 9998
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27816 9042 27844 9318
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27710 8528 27766 8537
rect 27710 8463 27712 8472
rect 27764 8463 27766 8472
rect 27712 8434 27764 8440
rect 27908 7410 27936 9454
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 27804 6384 27856 6390
rect 27802 6352 27804 6361
rect 27856 6352 27858 6361
rect 27908 6322 27936 7346
rect 27802 6287 27858 6296
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 27908 5234 27936 6258
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 28000 5137 28028 9862
rect 28078 8120 28134 8129
rect 28078 8055 28134 8064
rect 28092 8022 28120 8055
rect 28080 8016 28132 8022
rect 28080 7958 28132 7964
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 28092 6798 28120 7346
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 28092 5409 28120 6598
rect 28078 5400 28134 5409
rect 28078 5335 28134 5344
rect 27986 5128 28042 5137
rect 27986 5063 28042 5072
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 26974 4519 27030 4528
rect 27344 4548 27396 4554
rect 27344 4490 27396 4496
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26424 3732 26476 3738
rect 26424 3674 26476 3680
rect 26344 3534 26372 3674
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26148 3120 26200 3126
rect 26146 3088 26148 3097
rect 26200 3088 26202 3097
rect 26146 3023 26202 3032
rect 26344 2514 26372 3470
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 26056 2372 26108 2378
rect 26056 2314 26108 2320
rect 25596 2032 25648 2038
rect 25596 1974 25648 1980
rect 26436 800 26464 3674
rect 26804 3534 26832 3878
rect 27632 3738 27660 4422
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 26804 3194 26832 3470
rect 27068 3460 27120 3466
rect 26988 3420 27068 3448
rect 26884 3392 26936 3398
rect 26988 3380 27016 3420
rect 27068 3402 27120 3408
rect 27344 3460 27396 3466
rect 27724 3448 27752 3674
rect 27396 3420 27752 3448
rect 27344 3402 27396 3408
rect 26936 3352 27016 3380
rect 26884 3334 26936 3340
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 26620 2990 26648 3130
rect 27620 3120 27672 3126
rect 27618 3088 27620 3097
rect 27672 3088 27674 3097
rect 27618 3023 27674 3032
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 27712 2848 27764 2854
rect 27816 2825 27844 4558
rect 27712 2790 27764 2796
rect 27802 2816 27858 2825
rect 27724 800 27752 2790
rect 27802 2751 27858 2760
rect 28184 2530 28212 11698
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28276 3777 28304 11086
rect 28368 9994 28396 14350
rect 28446 14240 28502 14249
rect 28446 14175 28502 14184
rect 28460 13870 28488 14175
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28460 11898 28488 12038
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28460 11082 28488 11698
rect 28552 11150 28580 15370
rect 28644 15162 28672 15506
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28736 15042 28764 16934
rect 28644 15014 28764 15042
rect 28644 11626 28672 15014
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28632 11620 28684 11626
rect 28632 11562 28684 11568
rect 28736 11286 28764 12786
rect 28828 12434 28856 17138
rect 29012 15609 29040 17138
rect 28998 15600 29054 15609
rect 29104 15570 29132 20402
rect 29748 17762 29776 29514
rect 29840 20942 29868 31078
rect 29932 30326 29960 37198
rect 30944 37126 30972 39200
rect 31024 37256 31076 37262
rect 31024 37198 31076 37204
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 31036 36922 31064 37198
rect 32876 37108 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 33140 37120 33192 37126
rect 32876 37080 33140 37108
rect 34440 37108 34468 39222
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 35530 38176 35586 38185
rect 35530 38111 35586 38120
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 33140 37062 33192 37068
rect 34520 37062 34572 37068
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 34520 35692 34572 35698
rect 34520 35634 34572 35640
rect 29920 30320 29972 30326
rect 29920 30262 29972 30268
rect 34532 27470 34560 35634
rect 34808 29850 34836 37198
rect 35544 36922 35572 38111
rect 36096 37346 36124 39200
rect 36096 37318 36216 37346
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 35532 36916 35584 36922
rect 35532 36858 35584 36864
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35900 36712 35952 36718
rect 35900 36654 35952 36660
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35532 36168 35584 36174
rect 35530 36136 35532 36145
rect 35808 36168 35860 36174
rect 35584 36136 35586 36145
rect 35808 36110 35860 36116
rect 35530 36071 35586 36080
rect 35820 35698 35848 36110
rect 35808 35692 35860 35698
rect 35808 35634 35860 35640
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35808 31816 35860 31822
rect 35808 31758 35860 31764
rect 35820 31385 35848 31758
rect 35912 31482 35940 36654
rect 35900 31476 35952 31482
rect 35900 31418 35952 31424
rect 35806 31376 35862 31385
rect 35806 31311 35862 31320
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35348 27940 35400 27946
rect 35348 27882 35400 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 32508 19514 32536 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34244 21140 34296 21146
rect 34244 21082 34296 21088
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32324 18426 32352 19314
rect 32312 18420 32364 18426
rect 32312 18362 32364 18368
rect 29748 17734 29868 17762
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 28998 15535 29054 15544
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 29104 15162 29132 15506
rect 29092 15156 29144 15162
rect 29092 15098 29144 15104
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 29012 14414 29040 14894
rect 29000 14408 29052 14414
rect 29000 14350 29052 14356
rect 29104 14006 29132 15098
rect 29092 14000 29144 14006
rect 29092 13942 29144 13948
rect 29196 13394 29224 17206
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29288 14958 29316 15302
rect 29276 14952 29328 14958
rect 29276 14894 29328 14900
rect 29460 13864 29512 13870
rect 29460 13806 29512 13812
rect 29184 13388 29236 13394
rect 29184 13330 29236 13336
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28828 12406 28948 12434
rect 28816 11824 28868 11830
rect 28814 11792 28816 11801
rect 28868 11792 28870 11801
rect 28814 11727 28870 11736
rect 28724 11280 28776 11286
rect 28724 11222 28776 11228
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28448 11076 28500 11082
rect 28448 11018 28500 11024
rect 28356 9988 28408 9994
rect 28356 9930 28408 9936
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28368 7886 28396 8434
rect 28460 8362 28488 11018
rect 28644 11014 28672 11086
rect 28632 11008 28684 11014
rect 28632 10950 28684 10956
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28552 8401 28580 9318
rect 28538 8392 28594 8401
rect 28448 8356 28500 8362
rect 28538 8327 28594 8336
rect 28448 8298 28500 8304
rect 28460 7970 28488 8298
rect 28460 7942 28580 7970
rect 28552 7886 28580 7942
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28552 7410 28580 7822
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28552 6934 28580 7142
rect 28540 6928 28592 6934
rect 28540 6870 28592 6876
rect 28644 4622 28672 10950
rect 28736 10849 28764 11222
rect 28722 10840 28778 10849
rect 28722 10775 28778 10784
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28736 10198 28764 10542
rect 28724 10192 28776 10198
rect 28724 10134 28776 10140
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28736 8498 28764 9930
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28828 6798 28856 8366
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28736 5098 28764 6598
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28724 5092 28776 5098
rect 28724 5034 28776 5040
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28724 4480 28776 4486
rect 28722 4448 28724 4457
rect 28776 4448 28778 4457
rect 28722 4383 28778 4392
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28632 4072 28684 4078
rect 28632 4014 28684 4020
rect 28262 3768 28318 3777
rect 28552 3738 28580 4014
rect 28262 3703 28318 3712
rect 28540 3732 28592 3738
rect 28540 3674 28592 3680
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28356 3460 28408 3466
rect 28356 3402 28408 3408
rect 28368 3194 28396 3402
rect 28460 3369 28488 3470
rect 28446 3360 28502 3369
rect 28446 3295 28502 3304
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 28644 2650 28672 4014
rect 28828 3466 28856 5102
rect 28816 3460 28868 3466
rect 28816 3402 28868 3408
rect 28828 3126 28856 3402
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28184 2514 28672 2530
rect 28184 2508 28684 2514
rect 28184 2502 28632 2508
rect 28632 2450 28684 2456
rect 28828 2310 28856 3062
rect 28920 2514 28948 12406
rect 29012 11626 29040 13262
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29000 11620 29052 11626
rect 29000 11562 29052 11568
rect 29000 11280 29052 11286
rect 29000 11222 29052 11228
rect 29012 9586 29040 11222
rect 29104 9994 29132 12378
rect 29182 11384 29238 11393
rect 29182 11319 29238 11328
rect 29196 11150 29224 11319
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29196 10062 29224 10610
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29092 9988 29144 9994
rect 29092 9930 29144 9936
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29012 7954 29040 9522
rect 29196 9042 29224 9998
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29184 8900 29236 8906
rect 29184 8842 29236 8848
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 29012 7410 29040 7890
rect 29196 7546 29224 8842
rect 29288 8838 29316 12786
rect 29368 11620 29420 11626
rect 29368 11562 29420 11568
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29380 7818 29408 11562
rect 29368 7812 29420 7818
rect 29368 7754 29420 7760
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29012 6798 29040 7346
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 29012 4826 29040 4966
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29012 3942 29040 4082
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 28998 3632 29054 3641
rect 28998 3567 29054 3576
rect 29012 3398 29040 3567
rect 29000 3392 29052 3398
rect 29000 3334 29052 3340
rect 29000 3120 29052 3126
rect 28998 3088 29000 3097
rect 29052 3088 29054 3097
rect 28998 3023 29054 3032
rect 28908 2508 28960 2514
rect 28908 2450 28960 2456
rect 29104 2378 29132 6054
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29196 2582 29224 5510
rect 29472 5098 29500 13806
rect 29644 13728 29696 13734
rect 29644 13670 29696 13676
rect 29656 13258 29684 13670
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29748 12986 29776 17274
rect 29840 16794 29868 17734
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29840 15910 29868 16730
rect 30300 16658 30328 16934
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30288 16516 30340 16522
rect 30288 16458 30340 16464
rect 30300 16250 30328 16458
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 30288 16244 30340 16250
rect 30288 16186 30340 16192
rect 31128 16114 31156 16390
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 29932 15502 29960 15982
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 29828 15360 29880 15366
rect 29828 15302 29880 15308
rect 29840 15026 29868 15302
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 29828 12164 29880 12170
rect 29828 12106 29880 12112
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 29564 11150 29592 11698
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29656 9654 29684 12106
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29564 9110 29592 9590
rect 29552 9104 29604 9110
rect 29552 9046 29604 9052
rect 29564 7410 29592 9046
rect 29656 8838 29684 9590
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29564 6322 29592 7346
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29460 5092 29512 5098
rect 29460 5034 29512 5040
rect 29656 4214 29684 6054
rect 29644 4208 29696 4214
rect 29644 4150 29696 4156
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29564 3058 29592 3878
rect 29748 3670 29776 11698
rect 29840 11354 29868 12106
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29932 8922 29960 15438
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 30024 10674 30052 14758
rect 30484 14482 30512 15302
rect 31128 14890 31156 16050
rect 31116 14884 31168 14890
rect 31116 14826 31168 14832
rect 31760 14816 31812 14822
rect 31760 14758 31812 14764
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 31772 14414 31800 14758
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 31760 14408 31812 14414
rect 31760 14350 31812 14356
rect 30104 14340 30156 14346
rect 30104 14282 30156 14288
rect 30116 14006 30144 14282
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30484 14074 30512 14214
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30104 14000 30156 14006
rect 30104 13942 30156 13948
rect 30378 13968 30434 13977
rect 30378 13903 30380 13912
rect 30432 13903 30434 13912
rect 30380 13874 30432 13880
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12986 30328 13194
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30392 12152 30420 13398
rect 30472 12844 30524 12850
rect 30472 12786 30524 12792
rect 30484 12374 30512 12786
rect 30472 12368 30524 12374
rect 30472 12310 30524 12316
rect 30472 12164 30524 12170
rect 30392 12124 30472 12152
rect 30472 12106 30524 12112
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30116 11150 30144 11494
rect 30104 11144 30156 11150
rect 30104 11086 30156 11092
rect 30012 10668 30064 10674
rect 30012 10610 30064 10616
rect 29840 8498 29868 8910
rect 29932 8894 30052 8922
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 29840 7886 29868 8434
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 29932 3534 29960 8774
rect 30024 8566 30052 8894
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 30116 5302 30144 11086
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 30208 10130 30236 10610
rect 30380 10464 30432 10470
rect 30380 10406 30432 10412
rect 30392 10198 30420 10406
rect 30380 10192 30432 10198
rect 30380 10134 30432 10140
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 30392 9994 30420 10134
rect 30196 9988 30248 9994
rect 30196 9930 30248 9936
rect 30380 9988 30432 9994
rect 30380 9930 30432 9936
rect 30208 9042 30236 9930
rect 30576 9738 30604 14350
rect 31116 14272 31168 14278
rect 31116 14214 31168 14220
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30656 12640 30708 12646
rect 30656 12582 30708 12588
rect 30668 12322 30696 12582
rect 30760 12434 30788 12786
rect 30932 12708 30984 12714
rect 30932 12650 30984 12656
rect 30944 12442 30972 12650
rect 30932 12436 30984 12442
rect 30760 12406 30880 12434
rect 30668 12294 30788 12322
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30484 9710 30604 9738
rect 30196 9036 30248 9042
rect 30196 8978 30248 8984
rect 30288 8968 30340 8974
rect 30288 8910 30340 8916
rect 30300 7954 30328 8910
rect 30288 7948 30340 7954
rect 30288 7890 30340 7896
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30300 6322 30328 6734
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30300 5710 30328 6258
rect 30288 5704 30340 5710
rect 30288 5646 30340 5652
rect 30104 5296 30156 5302
rect 30104 5238 30156 5244
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 30024 4146 30052 5170
rect 30392 4185 30420 7142
rect 30378 4176 30434 4185
rect 30012 4140 30064 4146
rect 30378 4111 30434 4120
rect 30012 4082 30064 4088
rect 30484 4010 30512 9710
rect 30668 9654 30696 12106
rect 30564 9648 30616 9654
rect 30564 9590 30616 9596
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30576 4826 30604 9590
rect 30760 6769 30788 12294
rect 30746 6760 30802 6769
rect 30746 6695 30802 6704
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30472 4004 30524 4010
rect 30472 3946 30524 3952
rect 30760 3913 30788 4082
rect 30746 3904 30802 3913
rect 30746 3839 30802 3848
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29748 3398 29776 3470
rect 29736 3392 29788 3398
rect 29736 3334 29788 3340
rect 30852 3126 30880 12406
rect 30932 12378 30984 12384
rect 30944 10062 30972 12378
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 30840 3120 30892 3126
rect 30840 3062 30892 3068
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29184 2576 29236 2582
rect 29184 2518 29236 2524
rect 29092 2372 29144 2378
rect 29092 2314 29144 2320
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 29656 800 29684 2994
rect 31036 2854 31064 3334
rect 31128 2854 31156 14214
rect 31576 13796 31628 13802
rect 31576 13738 31628 13744
rect 31588 13530 31616 13738
rect 31576 13524 31628 13530
rect 31576 13466 31628 13472
rect 31588 13190 31616 13466
rect 31576 13184 31628 13190
rect 31576 13126 31628 13132
rect 31576 12980 31628 12986
rect 31576 12922 31628 12928
rect 31588 12782 31616 12922
rect 31576 12776 31628 12782
rect 31576 12718 31628 12724
rect 31588 12442 31616 12718
rect 31576 12436 31628 12442
rect 31576 12378 31628 12384
rect 31772 12170 31800 14350
rect 31760 12164 31812 12170
rect 31760 12106 31812 12112
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 31680 11150 31708 11494
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 31760 8900 31812 8906
rect 31760 8842 31812 8848
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31312 8090 31340 8230
rect 31300 8084 31352 8090
rect 31300 8026 31352 8032
rect 31772 5914 31800 8842
rect 31852 6724 31904 6730
rect 31852 6666 31904 6672
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 31220 3738 31248 5646
rect 31392 4276 31444 4282
rect 31392 4218 31444 4224
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31208 3732 31260 3738
rect 31208 3674 31260 3680
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 31116 2848 31168 2854
rect 31116 2790 31168 2796
rect 30576 2514 30604 2790
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 31312 2446 31340 3878
rect 31404 3738 31432 4218
rect 31760 4208 31812 4214
rect 31864 4196 31892 6666
rect 31812 4168 31892 4196
rect 31760 4150 31812 4156
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 31772 3534 31800 4150
rect 32048 3738 32076 9658
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 32036 3528 32088 3534
rect 32220 3528 32272 3534
rect 32088 3488 32220 3516
rect 32036 3470 32088 3476
rect 32220 3470 32272 3476
rect 31576 3460 31628 3466
rect 31576 3402 31628 3408
rect 31588 2922 31616 3402
rect 32416 3194 32444 12038
rect 32496 7880 32548 7886
rect 32496 7822 32548 7828
rect 32508 6798 32536 7822
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32508 3602 32536 6734
rect 32496 3596 32548 3602
rect 32496 3538 32548 3544
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 32404 3188 32456 3194
rect 32404 3130 32456 3136
rect 32968 3058 32996 3470
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 31576 2916 31628 2922
rect 31576 2858 31628 2864
rect 32864 2916 32916 2922
rect 32864 2858 32916 2864
rect 32876 2446 32904 2858
rect 34256 2650 34284 21082
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 12986 35388 27882
rect 35808 26512 35860 26518
rect 35808 26454 35860 26460
rect 35820 25945 35848 26454
rect 35806 25936 35862 25945
rect 35806 25871 35862 25880
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 35912 19446 35940 20878
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 36004 15162 36032 36722
rect 36096 35834 36124 37198
rect 36188 37126 36216 37318
rect 36176 37120 36228 37126
rect 36176 37062 36228 37068
rect 37384 36922 37412 39200
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 36084 35828 36136 35834
rect 36084 35770 36136 35776
rect 36360 35080 36412 35086
rect 36360 35022 36412 35028
rect 36372 34785 36400 35022
rect 36358 34776 36414 34785
rect 36358 34711 36360 34720
rect 36412 34711 36414 34720
rect 36360 34682 36412 34688
rect 36084 34536 36136 34542
rect 36084 34478 36136 34484
rect 36096 31958 36124 34478
rect 36360 32904 36412 32910
rect 36360 32846 36412 32852
rect 36372 32745 36400 32846
rect 36358 32736 36414 32745
rect 36358 32671 36414 32680
rect 36372 32570 36400 32671
rect 36360 32564 36412 32570
rect 36360 32506 36412 32512
rect 36084 31952 36136 31958
rect 36084 31894 36136 31900
rect 36360 29572 36412 29578
rect 36360 29514 36412 29520
rect 36372 29345 36400 29514
rect 36358 29336 36414 29345
rect 36358 29271 36360 29280
rect 36412 29271 36414 29280
rect 36360 29242 36412 29248
rect 36268 28076 36320 28082
rect 36268 28018 36320 28024
rect 36280 27985 36308 28018
rect 36266 27976 36322 27985
rect 36266 27911 36322 27920
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 36096 20602 36124 26318
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 36084 20596 36136 20602
rect 36084 20538 36136 20544
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 36096 15706 36124 19314
rect 36084 15700 36136 15706
rect 36084 15642 36136 15648
rect 36188 15162 36216 24006
rect 36372 23905 36400 24142
rect 36358 23896 36414 23905
rect 36358 23831 36414 23840
rect 36266 22536 36322 22545
rect 36266 22471 36268 22480
rect 36320 22471 36322 22480
rect 36268 22442 36320 22448
rect 36268 20800 36320 20806
rect 36268 20742 36320 20748
rect 36280 20505 36308 20742
rect 36266 20496 36322 20505
rect 36266 20431 36322 20440
rect 36268 19168 36320 19174
rect 36266 19136 36268 19145
rect 36320 19136 36322 19145
rect 36266 19071 36322 19080
rect 36266 17096 36322 17105
rect 36266 17031 36268 17040
rect 36320 17031 36322 17040
rect 36268 17002 36320 17008
rect 36268 15904 36320 15910
rect 36268 15846 36320 15852
rect 36280 15745 36308 15846
rect 36266 15736 36322 15745
rect 36266 15671 36322 15680
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 35900 13184 35952 13190
rect 35900 13126 35952 13132
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35532 11076 35584 11082
rect 35532 11018 35584 11024
rect 35544 10810 35572 11018
rect 35532 10804 35584 10810
rect 35532 10746 35584 10752
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35912 7478 35940 13126
rect 36004 10674 36032 14010
rect 36188 13394 36216 14962
rect 36360 13932 36412 13938
rect 36360 13874 36412 13880
rect 36372 13705 36400 13874
rect 36358 13696 36414 13705
rect 36358 13631 36414 13640
rect 36176 13388 36228 13394
rect 36176 13330 36228 13336
rect 36084 11620 36136 11626
rect 36084 11562 36136 11568
rect 36096 11257 36124 11562
rect 36082 11248 36138 11257
rect 36082 11183 36138 11192
rect 35992 10668 36044 10674
rect 35992 10610 36044 10616
rect 36004 9586 36032 10610
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 36084 9376 36136 9382
rect 36084 9318 36136 9324
rect 36096 8498 36124 9318
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35820 6905 35848 7346
rect 35806 6896 35862 6905
rect 35806 6831 35862 6840
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36188 5234 36216 13330
rect 36268 11756 36320 11762
rect 36268 11698 36320 11704
rect 36280 11665 36308 11698
rect 36266 11656 36322 11665
rect 36266 11591 36322 11600
rect 36268 10464 36320 10470
rect 36268 10406 36320 10412
rect 36280 10305 36308 10406
rect 36266 10296 36322 10305
rect 36266 10231 36322 10240
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36280 8265 36308 8298
rect 36266 8256 36322 8265
rect 36266 8191 36322 8200
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 36360 5160 36412 5166
rect 36360 5102 36412 5108
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36372 4865 36400 5102
rect 36358 4856 36414 4865
rect 36358 4791 36360 4800
rect 36412 4791 36414 4800
rect 36360 4762 36412 4768
rect 35898 4040 35954 4049
rect 35898 3975 35900 3984
rect 35952 3975 35954 3984
rect 35900 3946 35952 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35348 3664 35400 3670
rect 35348 3606 35400 3612
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 34256 2446 34284 2586
rect 35360 2446 35388 3606
rect 35912 3534 35940 3946
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36266 3496 36322 3505
rect 36266 3431 36322 3440
rect 36280 3398 36308 3431
rect 36268 3392 36320 3398
rect 36268 3334 36320 3340
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 34244 2440 34296 2446
rect 34244 2382 34296 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30944 800 30972 2246
rect 32876 800 32904 2382
rect 34428 2304 34480 2310
rect 34428 2246 34480 2252
rect 34164 870 34284 898
rect 34164 800 34192 870
rect 24596 734 24808 762
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 29642 200 29698 800
rect 30930 200 30986 800
rect 32862 200 32918 800
rect 34150 200 34206 800
rect 34256 762 34284 870
rect 34440 762 34468 2246
rect 34256 734 34468 762
rect 36004 105 36032 2994
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 36096 800 36124 2246
rect 36280 1465 36308 2994
rect 36266 1456 36322 1465
rect 36266 1391 36322 1400
rect 36082 200 36138 800
rect 35990 96 36046 105
rect 35990 31 36046 40
<< via2 >>
rect 2778 39480 2834 39536
rect 2410 38120 2466 38176
rect 1674 36100 1730 36136
rect 1674 36080 1676 36100
rect 1676 36080 1728 36100
rect 1728 36080 1730 36100
rect 1674 34720 1730 34776
rect 1674 32680 1730 32736
rect 1582 31356 1584 31376
rect 1584 31356 1636 31376
rect 1636 31356 1638 31376
rect 1582 31320 1638 31356
rect 1582 29300 1638 29336
rect 1582 29280 1584 29300
rect 1584 29280 1636 29300
rect 1636 29280 1638 29300
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1674 25880 1730 25936
rect 1582 23860 1638 23896
rect 1582 23840 1584 23860
rect 1584 23840 1636 23860
rect 1636 23840 1638 23860
rect 1674 22500 1730 22536
rect 1674 22480 1676 22500
rect 1676 22480 1728 22500
rect 1728 22480 1730 22500
rect 1582 20440 1638 20496
rect 1582 19080 1638 19136
rect 1674 17040 1730 17096
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1674 15680 1730 15736
rect 1674 13676 1676 13696
rect 1676 13676 1728 13696
rect 1728 13676 1730 13696
rect 1674 13640 1730 13676
rect 1674 11620 1730 11656
rect 1674 11600 1676 11620
rect 1676 11600 1728 11620
rect 1728 11600 1730 11620
rect 1674 10240 1730 10296
rect 1582 8200 1638 8256
rect 1582 6840 1638 6896
rect 1858 8356 1914 8392
rect 1858 8336 1860 8356
rect 1860 8336 1912 8356
rect 1912 8336 1914 8356
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2410 15952 2466 16008
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1582 4820 1638 4856
rect 1582 4800 1584 4820
rect 1584 4800 1636 4820
rect 1636 4800 1638 4820
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1674 3440 1730 3496
rect 2410 3052 2466 3088
rect 2410 3032 2412 3052
rect 2412 3032 2464 3052
rect 2464 3032 2466 3052
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 15658 37068 15660 37088
rect 15660 37068 15712 37088
rect 15712 37068 15714 37088
rect 15658 37032 15714 37068
rect 10782 12688 10838 12744
rect 10046 11192 10102 11248
rect 10506 10684 10508 10704
rect 10508 10684 10560 10704
rect 10560 10684 10562 10704
rect 10506 10648 10562 10684
rect 11150 11736 11206 11792
rect 10966 9324 10968 9344
rect 10968 9324 11020 9344
rect 11020 9324 11022 9344
rect 10966 9288 11022 9324
rect 2778 1400 2834 1456
rect 11610 15544 11666 15600
rect 12622 16108 12678 16144
rect 12622 16088 12624 16108
rect 12624 16088 12676 16108
rect 12676 16088 12678 16108
rect 11702 14356 11704 14376
rect 11704 14356 11756 14376
rect 11756 14356 11758 14376
rect 11702 14320 11758 14356
rect 11426 12860 11428 12880
rect 11428 12860 11480 12880
rect 11480 12860 11482 12880
rect 11426 12824 11482 12860
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 13726 16632 13782 16688
rect 13634 15408 13690 15464
rect 13542 14900 13544 14920
rect 13544 14900 13596 14920
rect 13596 14900 13598 14920
rect 13542 14864 13598 14900
rect 11610 12280 11666 12336
rect 11794 12280 11850 12336
rect 12898 12860 12900 12880
rect 12900 12860 12952 12880
rect 12952 12860 12954 12880
rect 12898 12824 12954 12860
rect 12530 12708 12586 12744
rect 12530 12688 12532 12708
rect 12532 12688 12584 12708
rect 12584 12688 12586 12708
rect 12254 12316 12256 12336
rect 12256 12316 12308 12336
rect 12308 12316 12310 12336
rect 12254 12280 12310 12316
rect 10874 2488 10930 2544
rect 10782 2372 10838 2408
rect 10782 2352 10784 2372
rect 10784 2352 10836 2372
rect 10836 2352 10838 2372
rect 11794 3440 11850 3496
rect 14370 16904 14426 16960
rect 14186 16088 14242 16144
rect 14002 13388 14058 13424
rect 14002 13368 14004 13388
rect 14004 13368 14056 13388
rect 14056 13368 14058 13388
rect 14002 9696 14058 9752
rect 14002 9288 14058 9344
rect 14002 8492 14058 8528
rect 14002 8472 14004 8492
rect 14004 8472 14056 8492
rect 14056 8472 14058 8492
rect 13726 6316 13782 6352
rect 13726 6296 13728 6316
rect 13728 6296 13780 6316
rect 13780 6296 13782 6316
rect 14462 14900 14464 14920
rect 14464 14900 14516 14920
rect 14516 14900 14518 14920
rect 14462 14864 14518 14900
rect 14278 12008 14334 12064
rect 13634 5636 13690 5672
rect 13634 5616 13636 5636
rect 13636 5616 13688 5636
rect 13688 5616 13690 5636
rect 13174 4800 13230 4856
rect 12990 4664 13046 4720
rect 13542 3576 13598 3632
rect 14554 9868 14556 9888
rect 14556 9868 14608 9888
rect 14608 9868 14610 9888
rect 14554 9832 14610 9868
rect 14830 10684 14832 10704
rect 14832 10684 14884 10704
rect 14884 10684 14886 10704
rect 14830 10648 14886 10684
rect 14830 10376 14886 10432
rect 15014 10376 15070 10432
rect 14738 8744 14794 8800
rect 14278 3476 14280 3496
rect 14280 3476 14332 3496
rect 14332 3476 14334 3496
rect 14278 3440 14334 3476
rect 12070 2896 12126 2952
rect 12714 2896 12770 2952
rect 13450 2896 13506 2952
rect 12438 2796 12440 2816
rect 12440 2796 12492 2816
rect 12492 2796 12494 2816
rect 12438 2760 12494 2796
rect 14462 2760 14518 2816
rect 13634 2624 13690 2680
rect 15566 13388 15622 13424
rect 15566 13368 15568 13388
rect 15568 13368 15620 13388
rect 15620 13368 15622 13388
rect 16026 17040 16082 17096
rect 16210 14320 16266 14376
rect 15658 9560 15714 9616
rect 15842 10648 15898 10704
rect 16026 10412 16028 10432
rect 16028 10412 16080 10432
rect 16080 10412 16082 10432
rect 16026 10376 16082 10412
rect 15934 8628 15990 8664
rect 15934 8608 15936 8628
rect 15936 8608 15988 8628
rect 15988 8608 15990 8628
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 16946 16652 17002 16688
rect 16946 16632 16948 16652
rect 16948 16632 17000 16652
rect 17000 16632 17002 16652
rect 15566 5072 15622 5128
rect 17222 15428 17278 15464
rect 17222 15408 17224 15428
rect 17224 15408 17276 15428
rect 17276 15408 17278 15428
rect 16670 9560 16726 9616
rect 16302 5752 16358 5808
rect 15014 3168 15070 3224
rect 16486 5244 16488 5264
rect 16488 5244 16540 5264
rect 16540 5244 16542 5264
rect 16486 5208 16542 5244
rect 18142 16904 18198 16960
rect 18510 15972 18566 16008
rect 18510 15952 18512 15972
rect 18512 15952 18564 15972
rect 18564 15952 18566 15972
rect 17130 12552 17186 12608
rect 17314 12416 17370 12472
rect 17038 9444 17094 9480
rect 17038 9424 17040 9444
rect 17040 9424 17092 9444
rect 17092 9424 17094 9444
rect 16854 8744 16910 8800
rect 18142 12824 18198 12880
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18878 17060 18934 17096
rect 18878 17040 18880 17060
rect 18880 17040 18932 17060
rect 18932 17040 18934 17060
rect 17682 9968 17738 10024
rect 17774 8628 17830 8664
rect 17774 8608 17776 8628
rect 17776 8608 17828 8628
rect 17828 8608 17830 8628
rect 18326 9832 18382 9888
rect 19338 16088 19394 16144
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19338 14220 19340 14240
rect 19340 14220 19392 14240
rect 19392 14220 19394 14240
rect 19338 14184 19394 14220
rect 19338 13268 19340 13288
rect 19340 13268 19392 13288
rect 19392 13268 19394 13288
rect 19338 13232 19394 13268
rect 18602 9288 18658 9344
rect 18234 4700 18236 4720
rect 18236 4700 18288 4720
rect 18288 4700 18290 4720
rect 18234 4664 18290 4700
rect 18510 4156 18512 4176
rect 18512 4156 18564 4176
rect 18564 4156 18566 4176
rect 18510 4120 18566 4156
rect 18878 9424 18934 9480
rect 18786 4820 18842 4856
rect 18786 4800 18788 4820
rect 18788 4800 18840 4820
rect 18840 4800 18842 4820
rect 16578 2896 16634 2952
rect 19246 12300 19302 12336
rect 19246 12280 19248 12300
rect 19248 12280 19300 12300
rect 19300 12280 19302 12300
rect 18970 3440 19026 3496
rect 18878 3032 18934 3088
rect 19246 12044 19248 12064
rect 19248 12044 19300 12064
rect 19300 12044 19302 12064
rect 19246 12008 19302 12044
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19890 12824 19946 12880
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20810 17620 20812 17640
rect 20812 17620 20864 17640
rect 20864 17620 20866 17640
rect 20810 17584 20866 17620
rect 20350 16108 20406 16144
rect 20350 16088 20352 16108
rect 20352 16088 20404 16108
rect 20404 16088 20406 16108
rect 20166 12688 20222 12744
rect 20350 13368 20406 13424
rect 20258 12280 20314 12336
rect 19246 10684 19248 10704
rect 19248 10684 19300 10704
rect 19300 10684 19302 10704
rect 19246 10648 19302 10684
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19614 10532 19670 10568
rect 19614 10512 19616 10532
rect 19616 10512 19668 10532
rect 19668 10512 19670 10532
rect 19982 10240 20038 10296
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20810 15136 20866 15192
rect 21822 18708 21824 18728
rect 21824 18708 21876 18728
rect 21876 18708 21878 18728
rect 21822 18672 21878 18708
rect 21270 15680 21326 15736
rect 21086 14864 21142 14920
rect 21822 16108 21878 16144
rect 21822 16088 21824 16108
rect 21824 16088 21876 16108
rect 21876 16088 21878 16108
rect 20626 13504 20682 13560
rect 21178 13232 21234 13288
rect 20902 12552 20958 12608
rect 20258 10240 20314 10296
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19982 8608 20038 8664
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19614 4528 19670 4584
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19338 3476 19340 3496
rect 19340 3476 19392 3496
rect 19392 3476 19394 3496
rect 19338 3440 19394 3476
rect 21178 12416 21234 12472
rect 22098 13776 22154 13832
rect 21086 10532 21142 10568
rect 21086 10512 21088 10532
rect 21088 10512 21140 10532
rect 21140 10512 21142 10532
rect 20442 4392 20498 4448
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20994 4528 21050 4584
rect 21086 3304 21142 3360
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21822 10260 21878 10296
rect 21822 10240 21824 10260
rect 21824 10240 21876 10260
rect 21876 10240 21878 10260
rect 21638 8472 21694 8528
rect 21822 8492 21878 8528
rect 21822 8472 21824 8492
rect 21824 8472 21876 8492
rect 21876 8472 21878 8492
rect 22098 9696 22154 9752
rect 22466 12688 22522 12744
rect 22650 13932 22706 13968
rect 22650 13912 22652 13932
rect 22652 13912 22704 13932
rect 22704 13912 22706 13932
rect 22650 13640 22706 13696
rect 22926 14764 22928 14784
rect 22928 14764 22980 14784
rect 22980 14764 22982 14784
rect 22926 14728 22982 14764
rect 22098 8064 22154 8120
rect 22006 6840 22062 6896
rect 21914 4276 21970 4312
rect 21914 4256 21916 4276
rect 21916 4256 21968 4276
rect 21968 4256 21970 4276
rect 21730 3440 21786 3496
rect 22466 3576 22522 3632
rect 22190 3032 22246 3088
rect 22466 3068 22468 3088
rect 22468 3068 22520 3088
rect 22520 3068 22522 3088
rect 22466 3032 22522 3068
rect 22742 8608 22798 8664
rect 22926 12008 22982 12064
rect 27434 36488 27490 36544
rect 23938 14900 23940 14920
rect 23940 14900 23992 14920
rect 23992 14900 23994 14920
rect 23938 14864 23994 14900
rect 23754 13776 23810 13832
rect 23018 11328 23074 11384
rect 22742 7520 22798 7576
rect 23110 8336 23166 8392
rect 23386 9968 23442 10024
rect 23754 11736 23810 11792
rect 23846 9460 23848 9480
rect 23848 9460 23900 9480
rect 23900 9460 23902 9480
rect 23846 9424 23902 9460
rect 23754 6704 23810 6760
rect 22834 4936 22890 4992
rect 24214 12844 24270 12880
rect 24214 12824 24216 12844
rect 24216 12824 24268 12844
rect 24268 12824 24270 12844
rect 24950 20884 24952 20904
rect 24952 20884 25004 20904
rect 25004 20884 25006 20904
rect 24950 20848 25006 20884
rect 24490 13640 24546 13696
rect 24766 12688 24822 12744
rect 23938 6568 23994 6624
rect 23294 3848 23350 3904
rect 23386 3712 23442 3768
rect 24674 11076 24730 11112
rect 24674 11056 24676 11076
rect 24676 11056 24728 11076
rect 24728 11056 24730 11076
rect 25318 11872 25374 11928
rect 25318 11600 25374 11656
rect 24858 10648 24914 10704
rect 24674 5752 24730 5808
rect 24398 5344 24454 5400
rect 24306 4684 24362 4720
rect 24306 4664 24308 4684
rect 24308 4664 24360 4684
rect 24360 4664 24362 4684
rect 24122 4528 24178 4584
rect 24858 4528 24914 4584
rect 25226 10104 25282 10160
rect 26698 18708 26700 18728
rect 26700 18708 26752 18728
rect 26752 18708 26754 18728
rect 26698 18672 26754 18708
rect 26238 14184 26294 14240
rect 25594 12416 25650 12472
rect 26514 15136 26570 15192
rect 26514 14048 26570 14104
rect 25778 12164 25834 12200
rect 25778 12144 25780 12164
rect 25780 12144 25832 12164
rect 25832 12144 25834 12164
rect 25870 11872 25926 11928
rect 25134 5752 25190 5808
rect 25778 9696 25834 9752
rect 25686 9596 25688 9616
rect 25688 9596 25740 9616
rect 25740 9596 25742 9616
rect 25686 9560 25742 9596
rect 25870 8472 25926 8528
rect 25042 3440 25098 3496
rect 24398 2760 24454 2816
rect 24674 2760 24730 2816
rect 26330 12724 26332 12744
rect 26332 12724 26384 12744
rect 26384 12724 26386 12744
rect 26330 12688 26386 12724
rect 25962 5752 26018 5808
rect 25962 4664 26018 4720
rect 25962 4392 26018 4448
rect 26238 6840 26294 6896
rect 26238 4936 26294 4992
rect 26514 13676 26516 13696
rect 26516 13676 26568 13696
rect 26568 13676 26570 13696
rect 26514 13640 26570 13676
rect 26790 14048 26846 14104
rect 26698 10784 26754 10840
rect 26790 9424 26846 9480
rect 26698 6568 26754 6624
rect 27066 12300 27122 12336
rect 27066 12280 27068 12300
rect 27068 12280 27120 12300
rect 27120 12280 27122 12300
rect 27342 16108 27398 16144
rect 27342 16088 27344 16108
rect 27344 16088 27396 16108
rect 27396 16088 27398 16108
rect 27250 14864 27306 14920
rect 27250 12008 27306 12064
rect 27342 11600 27398 11656
rect 27710 12416 27766 12472
rect 28170 14764 28172 14784
rect 28172 14764 28224 14784
rect 28224 14764 28226 14784
rect 28170 14728 28226 14764
rect 28078 12416 28134 12472
rect 27342 9696 27398 9752
rect 26698 4800 26754 4856
rect 26606 4276 26662 4312
rect 26606 4256 26608 4276
rect 26608 4256 26660 4276
rect 26660 4256 26662 4276
rect 26974 4528 27030 4584
rect 27802 9580 27858 9616
rect 27802 9560 27804 9580
rect 27804 9560 27856 9580
rect 27856 9560 27858 9580
rect 27710 8492 27766 8528
rect 27710 8472 27712 8492
rect 27712 8472 27764 8492
rect 27764 8472 27766 8492
rect 27802 6332 27804 6352
rect 27804 6332 27856 6352
rect 27856 6332 27858 6352
rect 27802 6296 27858 6332
rect 28078 8064 28134 8120
rect 28078 5344 28134 5400
rect 27986 5072 28042 5128
rect 26146 3068 26148 3088
rect 26148 3068 26200 3088
rect 26200 3068 26202 3088
rect 26146 3032 26202 3068
rect 27618 3068 27620 3088
rect 27620 3068 27672 3088
rect 27672 3068 27674 3088
rect 27618 3032 27674 3068
rect 27802 2760 27858 2816
rect 28446 14184 28502 14240
rect 28998 15544 29054 15600
rect 35530 38120 35586 38176
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35530 36116 35532 36136
rect 35532 36116 35584 36136
rect 35584 36116 35586 36136
rect 35530 36080 35586 36116
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35806 31320 35862 31376
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 28814 11772 28816 11792
rect 28816 11772 28868 11792
rect 28868 11772 28870 11792
rect 28814 11736 28870 11772
rect 28538 8336 28594 8392
rect 28722 10784 28778 10840
rect 28722 4428 28724 4448
rect 28724 4428 28776 4448
rect 28776 4428 28778 4448
rect 28722 4392 28778 4428
rect 28262 3712 28318 3768
rect 28446 3304 28502 3360
rect 29182 11328 29238 11384
rect 28998 3576 29054 3632
rect 28998 3068 29000 3088
rect 29000 3068 29052 3088
rect 29052 3068 29054 3088
rect 28998 3032 29054 3068
rect 30378 13932 30434 13968
rect 30378 13912 30380 13932
rect 30380 13912 30432 13932
rect 30432 13912 30434 13932
rect 30378 4120 30434 4176
rect 30746 6704 30802 6760
rect 30746 3848 30802 3904
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35806 25880 35862 25936
rect 36358 34740 36414 34776
rect 36358 34720 36360 34740
rect 36360 34720 36412 34740
rect 36412 34720 36414 34740
rect 36358 32680 36414 32736
rect 36358 29300 36414 29336
rect 36358 29280 36360 29300
rect 36360 29280 36412 29300
rect 36412 29280 36414 29300
rect 36266 27920 36322 27976
rect 36358 23840 36414 23896
rect 36266 22500 36322 22536
rect 36266 22480 36268 22500
rect 36268 22480 36320 22500
rect 36320 22480 36322 22500
rect 36266 20440 36322 20496
rect 36266 19116 36268 19136
rect 36268 19116 36320 19136
rect 36320 19116 36322 19136
rect 36266 19080 36322 19116
rect 36266 17060 36322 17096
rect 36266 17040 36268 17060
rect 36268 17040 36320 17060
rect 36320 17040 36322 17060
rect 36266 15680 36322 15736
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 36358 13640 36414 13696
rect 36082 11192 36138 11248
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35806 6840 35862 6896
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 36266 11600 36322 11656
rect 36266 10240 36322 10296
rect 36266 8200 36322 8256
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 36358 4820 36414 4856
rect 36358 4800 36360 4820
rect 36360 4800 36412 4820
rect 36412 4800 36414 4820
rect 35898 4004 35954 4040
rect 35898 3984 35900 4004
rect 35900 3984 35952 4004
rect 35952 3984 35954 4004
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36266 3440 36322 3496
rect 36266 1400 36322 1456
rect 35990 40 36046 96
<< metal3 >>
rect 200 39538 800 39568
rect 2773 39538 2839 39541
rect 200 39536 2839 39538
rect 200 39480 2778 39536
rect 2834 39480 2839 39536
rect 200 39478 2839 39480
rect 200 39448 800 39478
rect 2773 39475 2839 39478
rect 200 38178 800 38208
rect 2405 38178 2471 38181
rect 200 38176 2471 38178
rect 200 38120 2410 38176
rect 2466 38120 2471 38176
rect 200 38118 2471 38120
rect 200 38088 800 38118
rect 2405 38115 2471 38118
rect 35525 38178 35591 38181
rect 37200 38178 37800 38208
rect 35525 38176 37800 38178
rect 35525 38120 35530 38176
rect 35586 38120 37800 38176
rect 35525 38118 37800 38120
rect 35525 38115 35591 38118
rect 37200 38088 37800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 15653 37092 15719 37093
rect 15653 37090 15700 37092
rect 15608 37088 15700 37090
rect 15608 37032 15658 37088
rect 15608 37030 15700 37032
rect 15653 37028 15700 37030
rect 15764 37028 15770 37092
rect 15653 37027 15719 37028
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 27429 36548 27495 36549
rect 27429 36544 27476 36548
rect 27540 36546 27546 36548
rect 27429 36488 27434 36544
rect 27429 36484 27476 36488
rect 27540 36486 27586 36546
rect 27540 36484 27546 36486
rect 27429 36483 27495 36484
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 36048 800 36078
rect 1669 36075 1735 36078
rect 35525 36138 35591 36141
rect 37200 36138 37800 36168
rect 35525 36136 37800 36138
rect 35525 36080 35530 36136
rect 35586 36080 37800 36136
rect 35525 36078 37800 36080
rect 35525 36075 35591 36078
rect 37200 36048 37800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1669 34778 1735 34781
rect 200 34776 1735 34778
rect 200 34720 1674 34776
rect 1730 34720 1735 34776
rect 200 34718 1735 34720
rect 200 34688 800 34718
rect 1669 34715 1735 34718
rect 36353 34778 36419 34781
rect 37200 34778 37800 34808
rect 36353 34776 37800 34778
rect 36353 34720 36358 34776
rect 36414 34720 37800 34776
rect 36353 34718 37800 34720
rect 36353 34715 36419 34718
rect 37200 34688 37800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1669 32738 1735 32741
rect 200 32736 1735 32738
rect 200 32680 1674 32736
rect 1730 32680 1735 32736
rect 200 32678 1735 32680
rect 200 32648 800 32678
rect 1669 32675 1735 32678
rect 36353 32738 36419 32741
rect 37200 32738 37800 32768
rect 36353 32736 37800 32738
rect 36353 32680 36358 32736
rect 36414 32680 37800 32736
rect 36353 32678 37800 32680
rect 36353 32675 36419 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 37200 32648 37800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1577 31378 1643 31381
rect 200 31376 1643 31378
rect 200 31320 1582 31376
rect 1638 31320 1643 31376
rect 200 31318 1643 31320
rect 200 31288 800 31318
rect 1577 31315 1643 31318
rect 35801 31378 35867 31381
rect 37200 31378 37800 31408
rect 35801 31376 37800 31378
rect 35801 31320 35806 31376
rect 35862 31320 37800 31376
rect 35801 31318 37800 31320
rect 35801 31315 35867 31318
rect 37200 31288 37800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1577 29338 1643 29341
rect 200 29336 1643 29338
rect 200 29280 1582 29336
rect 1638 29280 1643 29336
rect 200 29278 1643 29280
rect 200 29248 800 29278
rect 1577 29275 1643 29278
rect 36353 29338 36419 29341
rect 37200 29338 37800 29368
rect 36353 29336 37800 29338
rect 36353 29280 36358 29336
rect 36414 29280 37800 29336
rect 36353 29278 37800 29280
rect 36353 29275 36419 29278
rect 37200 29248 37800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28008
rect 1669 27978 1735 27981
rect 200 27976 1735 27978
rect 200 27920 1674 27976
rect 1730 27920 1735 27976
rect 200 27918 1735 27920
rect 200 27888 800 27918
rect 1669 27915 1735 27918
rect 36261 27978 36327 27981
rect 37200 27978 37800 28008
rect 36261 27976 37800 27978
rect 36261 27920 36266 27976
rect 36322 27920 37800 27976
rect 36261 27918 37800 27920
rect 36261 27915 36327 27918
rect 37200 27888 37800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1669 25938 1735 25941
rect 200 25936 1735 25938
rect 200 25880 1674 25936
rect 1730 25880 1735 25936
rect 200 25878 1735 25880
rect 200 25848 800 25878
rect 1669 25875 1735 25878
rect 35801 25938 35867 25941
rect 37200 25938 37800 25968
rect 35801 25936 37800 25938
rect 35801 25880 35806 25936
rect 35862 25880 37800 25936
rect 35801 25878 37800 25880
rect 35801 25875 35867 25878
rect 37200 25848 37800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1577 23898 1643 23901
rect 200 23896 1643 23898
rect 200 23840 1582 23896
rect 1638 23840 1643 23896
rect 200 23838 1643 23840
rect 200 23808 800 23838
rect 1577 23835 1643 23838
rect 36353 23898 36419 23901
rect 37200 23898 37800 23928
rect 36353 23896 37800 23898
rect 36353 23840 36358 23896
rect 36414 23840 37800 23896
rect 36353 23838 37800 23840
rect 36353 23835 36419 23838
rect 37200 23808 37800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 36261 22538 36327 22541
rect 37200 22538 37800 22568
rect 36261 22536 37800 22538
rect 36261 22480 36266 22536
rect 36322 22480 37800 22536
rect 36261 22478 37800 22480
rect 36261 22475 36327 22478
rect 37200 22448 37800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 24945 20906 25011 20909
rect 25078 20906 25084 20908
rect 24945 20904 25084 20906
rect 24945 20848 24950 20904
rect 25006 20848 25084 20904
rect 24945 20846 25084 20848
rect 24945 20843 25011 20846
rect 25078 20844 25084 20846
rect 25148 20844 25154 20908
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1577 20498 1643 20501
rect 200 20496 1643 20498
rect 200 20440 1582 20496
rect 1638 20440 1643 20496
rect 200 20438 1643 20440
rect 200 20408 800 20438
rect 1577 20435 1643 20438
rect 36261 20498 36327 20501
rect 37200 20498 37800 20528
rect 36261 20496 37800 20498
rect 36261 20440 36266 20496
rect 36322 20440 37800 20496
rect 36261 20438 37800 20440
rect 36261 20435 36327 20438
rect 37200 20408 37800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 19138 800 19168
rect 1577 19138 1643 19141
rect 200 19136 1643 19138
rect 200 19080 1582 19136
rect 1638 19080 1643 19136
rect 200 19078 1643 19080
rect 200 19048 800 19078
rect 1577 19075 1643 19078
rect 36261 19138 36327 19141
rect 37200 19138 37800 19168
rect 36261 19136 37800 19138
rect 36261 19080 36266 19136
rect 36322 19080 37800 19136
rect 36261 19078 37800 19080
rect 36261 19075 36327 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 37200 19048 37800 19078
rect 34930 19007 35246 19008
rect 21817 18730 21883 18733
rect 26693 18730 26759 18733
rect 21817 18728 26759 18730
rect 21817 18672 21822 18728
rect 21878 18672 26698 18728
rect 26754 18672 26759 18728
rect 21817 18670 26759 18672
rect 21817 18667 21883 18670
rect 26693 18667 26759 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 20805 17644 20871 17645
rect 20805 17642 20852 17644
rect 20760 17640 20852 17642
rect 20760 17584 20810 17640
rect 20760 17582 20852 17584
rect 20805 17580 20852 17582
rect 20916 17580 20922 17644
rect 20805 17579 20871 17580
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 200 17098 800 17128
rect 1669 17098 1735 17101
rect 200 17096 1735 17098
rect 200 17040 1674 17096
rect 1730 17040 1735 17096
rect 200 17038 1735 17040
rect 200 17008 800 17038
rect 1669 17035 1735 17038
rect 16021 17098 16087 17101
rect 18873 17098 18939 17101
rect 16021 17096 18939 17098
rect 16021 17040 16026 17096
rect 16082 17040 18878 17096
rect 18934 17040 18939 17096
rect 16021 17038 18939 17040
rect 16021 17035 16087 17038
rect 18873 17035 18939 17038
rect 36261 17098 36327 17101
rect 37200 17098 37800 17128
rect 36261 17096 37800 17098
rect 36261 17040 36266 17096
rect 36322 17040 37800 17096
rect 36261 17038 37800 17040
rect 36261 17035 36327 17038
rect 37200 17008 37800 17038
rect 14365 16962 14431 16965
rect 18137 16962 18203 16965
rect 14365 16960 18203 16962
rect 14365 16904 14370 16960
rect 14426 16904 18142 16960
rect 18198 16904 18203 16960
rect 14365 16902 18203 16904
rect 14365 16899 14431 16902
rect 18137 16899 18203 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 13721 16690 13787 16693
rect 16941 16690 17007 16693
rect 13721 16688 17007 16690
rect 13721 16632 13726 16688
rect 13782 16632 16946 16688
rect 17002 16632 17007 16688
rect 13721 16630 17007 16632
rect 13721 16627 13787 16630
rect 16941 16627 17007 16630
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 12617 16146 12683 16149
rect 14181 16146 14247 16149
rect 12617 16144 14247 16146
rect 12617 16088 12622 16144
rect 12678 16088 14186 16144
rect 14242 16088 14247 16144
rect 12617 16086 14247 16088
rect 12617 16083 12683 16086
rect 14181 16083 14247 16086
rect 19333 16148 19399 16149
rect 19333 16144 19380 16148
rect 19444 16146 19450 16148
rect 20345 16146 20411 16149
rect 19444 16144 20411 16146
rect 19333 16088 19338 16144
rect 19444 16088 20350 16144
rect 20406 16088 20411 16144
rect 19333 16084 19380 16088
rect 19444 16086 20411 16088
rect 19444 16084 19450 16086
rect 19333 16083 19399 16084
rect 20345 16083 20411 16086
rect 21817 16146 21883 16149
rect 27337 16146 27403 16149
rect 21817 16144 27403 16146
rect 21817 16088 21822 16144
rect 21878 16088 27342 16144
rect 27398 16088 27403 16144
rect 21817 16086 27403 16088
rect 21817 16083 21883 16086
rect 27337 16083 27403 16086
rect 2405 16010 2471 16013
rect 18505 16010 18571 16013
rect 2405 16008 18571 16010
rect 2405 15952 2410 16008
rect 2466 15952 18510 16008
rect 18566 15952 18571 16008
rect 2405 15950 18571 15952
rect 2405 15947 2471 15950
rect 18505 15947 18571 15950
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 21265 15738 21331 15741
rect 21398 15738 21404 15740
rect 21265 15736 21404 15738
rect 21265 15680 21270 15736
rect 21326 15680 21404 15736
rect 21265 15678 21404 15680
rect 21265 15675 21331 15678
rect 21398 15676 21404 15678
rect 21468 15676 21474 15740
rect 36261 15738 36327 15741
rect 37200 15738 37800 15768
rect 36261 15736 37800 15738
rect 36261 15680 36266 15736
rect 36322 15680 37800 15736
rect 36261 15678 37800 15680
rect 36261 15675 36327 15678
rect 37200 15648 37800 15678
rect 11605 15602 11671 15605
rect 28993 15602 29059 15605
rect 11605 15600 29059 15602
rect 11605 15544 11610 15600
rect 11666 15544 28998 15600
rect 29054 15544 29059 15600
rect 11605 15542 29059 15544
rect 11605 15539 11671 15542
rect 28993 15539 29059 15542
rect 13629 15466 13695 15469
rect 17217 15466 17283 15469
rect 13629 15464 17283 15466
rect 13629 15408 13634 15464
rect 13690 15408 17222 15464
rect 17278 15408 17283 15464
rect 13629 15406 17283 15408
rect 13629 15403 13695 15406
rect 17217 15403 17283 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 20805 15194 20871 15197
rect 26509 15194 26575 15197
rect 20805 15192 26575 15194
rect 20805 15136 20810 15192
rect 20866 15136 26514 15192
rect 26570 15136 26575 15192
rect 20805 15134 26575 15136
rect 20805 15131 20871 15134
rect 26509 15131 26575 15134
rect 13537 14922 13603 14925
rect 14457 14922 14523 14925
rect 13537 14920 14523 14922
rect 13537 14864 13542 14920
rect 13598 14864 14462 14920
rect 14518 14864 14523 14920
rect 13537 14862 14523 14864
rect 13537 14859 13603 14862
rect 14457 14859 14523 14862
rect 21081 14922 21147 14925
rect 23933 14922 23999 14925
rect 27245 14922 27311 14925
rect 21081 14920 27311 14922
rect 21081 14864 21086 14920
rect 21142 14864 23938 14920
rect 23994 14864 27250 14920
rect 27306 14864 27311 14920
rect 21081 14862 27311 14864
rect 21081 14859 21147 14862
rect 23933 14859 23999 14862
rect 27245 14859 27311 14862
rect 22921 14786 22987 14789
rect 28165 14786 28231 14789
rect 22921 14784 28231 14786
rect 22921 14728 22926 14784
rect 22982 14728 28170 14784
rect 28226 14728 28231 14784
rect 22921 14726 28231 14728
rect 22921 14723 22987 14726
rect 28165 14723 28231 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 11697 14378 11763 14381
rect 16205 14378 16271 14381
rect 11697 14376 16271 14378
rect 11697 14320 11702 14376
rect 11758 14320 16210 14376
rect 16266 14320 16271 14376
rect 11697 14318 16271 14320
rect 11697 14315 11763 14318
rect 16205 14315 16271 14318
rect 19333 14244 19399 14245
rect 19333 14240 19380 14244
rect 19444 14242 19450 14244
rect 26233 14242 26299 14245
rect 28441 14242 28507 14245
rect 19333 14184 19338 14240
rect 19333 14180 19380 14184
rect 19444 14182 19490 14242
rect 26233 14240 28507 14242
rect 26233 14184 26238 14240
rect 26294 14184 28446 14240
rect 28502 14184 28507 14240
rect 26233 14182 28507 14184
rect 19444 14180 19450 14182
rect 19333 14179 19399 14180
rect 26233 14179 26299 14182
rect 28441 14179 28507 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 26509 14106 26575 14109
rect 26785 14106 26851 14109
rect 26509 14104 26851 14106
rect 26509 14048 26514 14104
rect 26570 14048 26790 14104
rect 26846 14048 26851 14104
rect 26509 14046 26851 14048
rect 26509 14043 26575 14046
rect 26785 14043 26851 14046
rect 22645 13970 22711 13973
rect 30373 13970 30439 13973
rect 22645 13968 30439 13970
rect 22645 13912 22650 13968
rect 22706 13912 30378 13968
rect 30434 13912 30439 13968
rect 22645 13910 30439 13912
rect 22645 13907 22711 13910
rect 30373 13907 30439 13910
rect 22093 13834 22159 13837
rect 23749 13834 23815 13837
rect 22093 13832 23815 13834
rect 22093 13776 22098 13832
rect 22154 13776 23754 13832
rect 23810 13776 23815 13832
rect 22093 13774 23815 13776
rect 22093 13771 22159 13774
rect 23749 13771 23815 13774
rect 200 13698 800 13728
rect 1669 13698 1735 13701
rect 200 13696 1735 13698
rect 200 13640 1674 13696
rect 1730 13640 1735 13696
rect 200 13638 1735 13640
rect 200 13608 800 13638
rect 1669 13635 1735 13638
rect 22502 13636 22508 13700
rect 22572 13698 22578 13700
rect 22645 13698 22711 13701
rect 22572 13696 22711 13698
rect 22572 13640 22650 13696
rect 22706 13640 22711 13696
rect 22572 13638 22711 13640
rect 22572 13636 22578 13638
rect 22645 13635 22711 13638
rect 24485 13698 24551 13701
rect 26509 13698 26575 13701
rect 24485 13696 26575 13698
rect 24485 13640 24490 13696
rect 24546 13640 26514 13696
rect 26570 13640 26575 13696
rect 24485 13638 26575 13640
rect 24485 13635 24551 13638
rect 26509 13635 26575 13638
rect 36353 13698 36419 13701
rect 37200 13698 37800 13728
rect 36353 13696 37800 13698
rect 36353 13640 36358 13696
rect 36414 13640 37800 13696
rect 36353 13638 37800 13640
rect 36353 13635 36419 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 37200 13608 37800 13638
rect 34930 13567 35246 13568
rect 20621 13562 20687 13565
rect 20486 13560 20687 13562
rect 20486 13504 20626 13560
rect 20682 13504 20687 13560
rect 20486 13502 20687 13504
rect 13997 13426 14063 13429
rect 15561 13426 15627 13429
rect 13997 13424 15627 13426
rect 13997 13368 14002 13424
rect 14058 13368 15566 13424
rect 15622 13368 15627 13424
rect 13997 13366 15627 13368
rect 13997 13363 14063 13366
rect 15561 13363 15627 13366
rect 20345 13426 20411 13429
rect 20486 13426 20546 13502
rect 20621 13499 20687 13502
rect 20345 13424 20546 13426
rect 20345 13368 20350 13424
rect 20406 13368 20546 13424
rect 20345 13366 20546 13368
rect 20345 13363 20411 13366
rect 19333 13290 19399 13293
rect 21173 13290 21239 13293
rect 19333 13288 21239 13290
rect 19333 13232 19338 13288
rect 19394 13232 21178 13288
rect 21234 13232 21239 13288
rect 19333 13230 21239 13232
rect 19333 13227 19399 13230
rect 21173 13227 21239 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 11421 12882 11487 12885
rect 12893 12882 12959 12885
rect 11421 12880 12959 12882
rect 11421 12824 11426 12880
rect 11482 12824 12898 12880
rect 12954 12824 12959 12880
rect 11421 12822 12959 12824
rect 11421 12819 11487 12822
rect 12893 12819 12959 12822
rect 18137 12882 18203 12885
rect 18270 12882 18276 12884
rect 18137 12880 18276 12882
rect 18137 12824 18142 12880
rect 18198 12824 18276 12880
rect 18137 12822 18276 12824
rect 18137 12819 18203 12822
rect 18270 12820 18276 12822
rect 18340 12820 18346 12884
rect 19885 12882 19951 12885
rect 24209 12882 24275 12885
rect 19885 12880 24275 12882
rect 19885 12824 19890 12880
rect 19946 12824 24214 12880
rect 24270 12824 24275 12880
rect 19885 12822 24275 12824
rect 19885 12819 19951 12822
rect 24209 12819 24275 12822
rect 10777 12746 10843 12749
rect 12525 12746 12591 12749
rect 10777 12744 12591 12746
rect 10777 12688 10782 12744
rect 10838 12688 12530 12744
rect 12586 12688 12591 12744
rect 10777 12686 12591 12688
rect 10777 12683 10843 12686
rect 12525 12683 12591 12686
rect 20161 12746 20227 12749
rect 22461 12746 22527 12749
rect 20161 12744 22527 12746
rect 20161 12688 20166 12744
rect 20222 12688 22466 12744
rect 22522 12688 22527 12744
rect 20161 12686 22527 12688
rect 20161 12683 20227 12686
rect 22461 12683 22527 12686
rect 24761 12746 24827 12749
rect 26325 12746 26391 12749
rect 24761 12744 26391 12746
rect 24761 12688 24766 12744
rect 24822 12688 26330 12744
rect 26386 12688 26391 12744
rect 24761 12686 26391 12688
rect 24761 12683 24827 12686
rect 26325 12683 26391 12686
rect 17125 12610 17191 12613
rect 20897 12610 20963 12613
rect 17125 12608 20963 12610
rect 17125 12552 17130 12608
rect 17186 12552 20902 12608
rect 20958 12552 20963 12608
rect 17125 12550 20963 12552
rect 17125 12547 17191 12550
rect 20897 12547 20963 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 17309 12474 17375 12477
rect 21173 12474 21239 12477
rect 17309 12472 21239 12474
rect 17309 12416 17314 12472
rect 17370 12416 21178 12472
rect 21234 12416 21239 12472
rect 17309 12414 21239 12416
rect 17309 12411 17375 12414
rect 21173 12411 21239 12414
rect 25589 12474 25655 12477
rect 27705 12474 27771 12477
rect 28073 12474 28139 12477
rect 25589 12472 28139 12474
rect 25589 12416 25594 12472
rect 25650 12416 27710 12472
rect 27766 12416 28078 12472
rect 28134 12416 28139 12472
rect 25589 12414 28139 12416
rect 25589 12411 25655 12414
rect 27705 12411 27771 12414
rect 28073 12411 28139 12414
rect 11605 12338 11671 12341
rect 11470 12336 11671 12338
rect 11470 12280 11610 12336
rect 11666 12280 11671 12336
rect 11470 12278 11671 12280
rect 11145 11794 11211 11797
rect 11470 11794 11530 12278
rect 11605 12275 11671 12278
rect 11789 12338 11855 12341
rect 12249 12338 12315 12341
rect 11789 12336 12315 12338
rect 11789 12280 11794 12336
rect 11850 12280 12254 12336
rect 12310 12280 12315 12336
rect 11789 12278 12315 12280
rect 11789 12275 11855 12278
rect 12249 12275 12315 12278
rect 19241 12338 19307 12341
rect 20253 12338 20319 12341
rect 27061 12338 27127 12341
rect 19241 12336 27127 12338
rect 19241 12280 19246 12336
rect 19302 12280 20258 12336
rect 20314 12280 27066 12336
rect 27122 12280 27127 12336
rect 19241 12278 27127 12280
rect 19241 12275 19307 12278
rect 20253 12275 20319 12278
rect 27061 12275 27127 12278
rect 15694 12140 15700 12204
rect 15764 12202 15770 12204
rect 25773 12202 25839 12205
rect 15764 12200 25839 12202
rect 15764 12144 25778 12200
rect 25834 12144 25839 12200
rect 15764 12142 25839 12144
rect 15764 12140 15770 12142
rect 25773 12139 25839 12142
rect 14273 12066 14339 12069
rect 19241 12066 19307 12069
rect 14273 12064 19307 12066
rect 14273 12008 14278 12064
rect 14334 12008 19246 12064
rect 19302 12008 19307 12064
rect 14273 12006 19307 12008
rect 14273 12003 14339 12006
rect 19241 12003 19307 12006
rect 22921 12066 22987 12069
rect 27245 12066 27311 12069
rect 22921 12064 27311 12066
rect 22921 12008 22926 12064
rect 22982 12008 27250 12064
rect 27306 12008 27311 12064
rect 22921 12006 27311 12008
rect 22921 12003 22987 12006
rect 27245 12003 27311 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 25313 11930 25379 11933
rect 25865 11930 25931 11933
rect 25313 11928 25931 11930
rect 25313 11872 25318 11928
rect 25374 11872 25870 11928
rect 25926 11872 25931 11928
rect 25313 11870 25931 11872
rect 25313 11867 25379 11870
rect 25865 11867 25931 11870
rect 11145 11792 11530 11794
rect 11145 11736 11150 11792
rect 11206 11736 11530 11792
rect 11145 11734 11530 11736
rect 23749 11794 23815 11797
rect 28809 11794 28875 11797
rect 23749 11792 28875 11794
rect 23749 11736 23754 11792
rect 23810 11736 28814 11792
rect 28870 11736 28875 11792
rect 23749 11734 28875 11736
rect 11145 11731 11211 11734
rect 23749 11731 23815 11734
rect 28809 11731 28875 11734
rect 200 11658 800 11688
rect 1669 11658 1735 11661
rect 200 11656 1735 11658
rect 200 11600 1674 11656
rect 1730 11600 1735 11656
rect 200 11598 1735 11600
rect 200 11568 800 11598
rect 1669 11595 1735 11598
rect 25313 11658 25379 11661
rect 27337 11658 27403 11661
rect 25313 11656 27403 11658
rect 25313 11600 25318 11656
rect 25374 11600 27342 11656
rect 27398 11600 27403 11656
rect 25313 11598 27403 11600
rect 25313 11595 25379 11598
rect 27337 11595 27403 11598
rect 36261 11658 36327 11661
rect 37200 11658 37800 11688
rect 36261 11656 37800 11658
rect 36261 11600 36266 11656
rect 36322 11600 37800 11656
rect 36261 11598 37800 11600
rect 36261 11595 36327 11598
rect 37200 11568 37800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 23013 11386 23079 11389
rect 29177 11386 29243 11389
rect 23013 11384 29243 11386
rect 23013 11328 23018 11384
rect 23074 11328 29182 11384
rect 29238 11328 29243 11384
rect 23013 11326 29243 11328
rect 23013 11323 23079 11326
rect 29177 11323 29243 11326
rect 10041 11250 10107 11253
rect 36077 11250 36143 11253
rect 10041 11248 36143 11250
rect 10041 11192 10046 11248
rect 10102 11192 36082 11248
rect 36138 11192 36143 11248
rect 10041 11190 36143 11192
rect 10041 11187 10107 11190
rect 36077 11187 36143 11190
rect 23422 11052 23428 11116
rect 23492 11114 23498 11116
rect 24669 11114 24735 11117
rect 23492 11112 24735 11114
rect 23492 11056 24674 11112
rect 24730 11056 24735 11112
rect 23492 11054 24735 11056
rect 23492 11052 23498 11054
rect 24669 11051 24735 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 26693 10842 26759 10845
rect 28717 10842 28783 10845
rect 26693 10840 28783 10842
rect 26693 10784 26698 10840
rect 26754 10784 28722 10840
rect 28778 10784 28783 10840
rect 26693 10782 28783 10784
rect 26693 10779 26759 10782
rect 28717 10779 28783 10782
rect 10501 10706 10567 10709
rect 14825 10706 14891 10709
rect 15837 10706 15903 10709
rect 10501 10704 15903 10706
rect 10501 10648 10506 10704
rect 10562 10648 14830 10704
rect 14886 10648 15842 10704
rect 15898 10648 15903 10704
rect 10501 10646 15903 10648
rect 10501 10643 10567 10646
rect 14825 10643 14891 10646
rect 15837 10643 15903 10646
rect 19241 10706 19307 10709
rect 24853 10706 24919 10709
rect 19241 10704 24919 10706
rect 19241 10648 19246 10704
rect 19302 10648 24858 10704
rect 24914 10648 24919 10704
rect 19241 10646 24919 10648
rect 19241 10643 19307 10646
rect 24853 10643 24919 10646
rect 19609 10570 19675 10573
rect 21081 10570 21147 10573
rect 19609 10568 21147 10570
rect 19609 10512 19614 10568
rect 19670 10512 21086 10568
rect 21142 10512 21147 10568
rect 19609 10510 21147 10512
rect 19609 10507 19675 10510
rect 21081 10507 21147 10510
rect 14825 10434 14891 10437
rect 15009 10434 15075 10437
rect 16021 10434 16087 10437
rect 14825 10432 16087 10434
rect 14825 10376 14830 10432
rect 14886 10376 15014 10432
rect 15070 10376 16026 10432
rect 16082 10376 16087 10432
rect 14825 10374 16087 10376
rect 14825 10371 14891 10374
rect 15009 10371 15075 10374
rect 16021 10371 16087 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 200 10296 1735 10298
rect 200 10240 1674 10296
rect 1730 10240 1735 10296
rect 200 10238 1735 10240
rect 200 10208 800 10238
rect 1669 10235 1735 10238
rect 19374 10236 19380 10300
rect 19444 10298 19450 10300
rect 19977 10298 20043 10301
rect 19444 10296 20043 10298
rect 19444 10240 19982 10296
rect 20038 10240 20043 10296
rect 19444 10238 20043 10240
rect 19444 10236 19450 10238
rect 19977 10235 20043 10238
rect 20253 10298 20319 10301
rect 21817 10298 21883 10301
rect 20253 10296 21883 10298
rect 20253 10240 20258 10296
rect 20314 10240 21822 10296
rect 21878 10240 21883 10296
rect 20253 10238 21883 10240
rect 20253 10235 20319 10238
rect 21817 10235 21883 10238
rect 36261 10298 36327 10301
rect 37200 10298 37800 10328
rect 36261 10296 37800 10298
rect 36261 10240 36266 10296
rect 36322 10240 37800 10296
rect 36261 10238 37800 10240
rect 36261 10235 36327 10238
rect 37200 10208 37800 10238
rect 14958 10100 14964 10164
rect 15028 10162 15034 10164
rect 25221 10162 25287 10165
rect 15028 10160 25287 10162
rect 15028 10104 25226 10160
rect 25282 10104 25287 10160
rect 15028 10102 25287 10104
rect 15028 10100 15034 10102
rect 25221 10099 25287 10102
rect 17677 10026 17743 10029
rect 23381 10026 23447 10029
rect 17677 10024 23447 10026
rect 17677 9968 17682 10024
rect 17738 9968 23386 10024
rect 23442 9968 23447 10024
rect 17677 9966 23447 9968
rect 17677 9963 17743 9966
rect 23381 9963 23447 9966
rect 14549 9890 14615 9893
rect 18321 9890 18387 9893
rect 14549 9888 18387 9890
rect 14549 9832 14554 9888
rect 14610 9832 18326 9888
rect 18382 9832 18387 9888
rect 14549 9830 18387 9832
rect 14549 9827 14615 9830
rect 18321 9827 18387 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 13997 9754 14063 9757
rect 22093 9756 22159 9757
rect 15142 9754 15148 9756
rect 13997 9752 15148 9754
rect 13997 9696 14002 9752
rect 14058 9696 15148 9752
rect 13997 9694 15148 9696
rect 13997 9691 14063 9694
rect 15142 9692 15148 9694
rect 15212 9692 15218 9756
rect 22093 9752 22140 9756
rect 22204 9754 22210 9756
rect 25773 9754 25839 9757
rect 27337 9754 27403 9757
rect 22093 9696 22098 9752
rect 22093 9692 22140 9696
rect 22204 9694 22250 9754
rect 25773 9752 27403 9754
rect 25773 9696 25778 9752
rect 25834 9696 27342 9752
rect 27398 9696 27403 9752
rect 25773 9694 27403 9696
rect 22204 9692 22210 9694
rect 22093 9691 22159 9692
rect 25773 9691 25839 9694
rect 27337 9691 27403 9694
rect 15653 9618 15719 9621
rect 16665 9618 16731 9621
rect 15653 9616 16731 9618
rect 15653 9560 15658 9616
rect 15714 9560 16670 9616
rect 16726 9560 16731 9616
rect 15653 9558 16731 9560
rect 15653 9555 15719 9558
rect 16665 9555 16731 9558
rect 25681 9618 25747 9621
rect 27797 9618 27863 9621
rect 25681 9616 27863 9618
rect 25681 9560 25686 9616
rect 25742 9560 27802 9616
rect 27858 9560 27863 9616
rect 25681 9558 27863 9560
rect 25681 9555 25747 9558
rect 27797 9555 27863 9558
rect 17033 9482 17099 9485
rect 18873 9482 18939 9485
rect 17033 9480 18939 9482
rect 17033 9424 17038 9480
rect 17094 9424 18878 9480
rect 18934 9424 18939 9480
rect 17033 9422 18939 9424
rect 17033 9419 17099 9422
rect 18873 9419 18939 9422
rect 23841 9482 23907 9485
rect 26785 9482 26851 9485
rect 23841 9480 26851 9482
rect 23841 9424 23846 9480
rect 23902 9424 26790 9480
rect 26846 9424 26851 9480
rect 23841 9422 26851 9424
rect 23841 9419 23907 9422
rect 26785 9419 26851 9422
rect 10961 9346 11027 9349
rect 13997 9346 14063 9349
rect 18597 9346 18663 9349
rect 10961 9344 18663 9346
rect 10961 9288 10966 9344
rect 11022 9288 14002 9344
rect 14058 9288 18602 9344
rect 18658 9288 18663 9344
rect 10961 9286 18663 9288
rect 10961 9283 11027 9286
rect 13997 9283 14063 9286
rect 18597 9283 18663 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 14733 8802 14799 8805
rect 16849 8802 16915 8805
rect 14733 8800 16915 8802
rect 14733 8744 14738 8800
rect 14794 8744 16854 8800
rect 16910 8744 16915 8800
rect 14733 8742 16915 8744
rect 14733 8739 14799 8742
rect 16849 8739 16915 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 15929 8666 15995 8669
rect 17769 8666 17835 8669
rect 15929 8664 17835 8666
rect 15929 8608 15934 8664
rect 15990 8608 17774 8664
rect 17830 8608 17835 8664
rect 15929 8606 17835 8608
rect 15929 8603 15995 8606
rect 17769 8603 17835 8606
rect 19977 8666 20043 8669
rect 22737 8666 22803 8669
rect 19977 8664 22803 8666
rect 19977 8608 19982 8664
rect 20038 8608 22742 8664
rect 22798 8608 22803 8664
rect 19977 8606 22803 8608
rect 19977 8603 20043 8606
rect 22737 8603 22803 8606
rect 13997 8530 14063 8533
rect 21633 8530 21699 8533
rect 13997 8528 21699 8530
rect 13997 8472 14002 8528
rect 14058 8472 21638 8528
rect 21694 8472 21699 8528
rect 13997 8470 21699 8472
rect 13997 8467 14063 8470
rect 21633 8467 21699 8470
rect 21817 8530 21883 8533
rect 25865 8530 25931 8533
rect 27705 8530 27771 8533
rect 21817 8528 27771 8530
rect 21817 8472 21822 8528
rect 21878 8472 25870 8528
rect 25926 8472 27710 8528
rect 27766 8472 27771 8528
rect 21817 8470 27771 8472
rect 21817 8467 21883 8470
rect 25865 8467 25931 8470
rect 27705 8467 27771 8470
rect 1853 8394 1919 8397
rect 23105 8394 23171 8397
rect 1853 8392 23171 8394
rect 1853 8336 1858 8392
rect 1914 8336 23110 8392
rect 23166 8336 23171 8392
rect 1853 8334 23171 8336
rect 1853 8331 1919 8334
rect 23105 8331 23171 8334
rect 27654 8332 27660 8396
rect 27724 8394 27730 8396
rect 28533 8394 28599 8397
rect 27724 8392 28599 8394
rect 27724 8336 28538 8392
rect 28594 8336 28599 8392
rect 27724 8334 28599 8336
rect 27724 8332 27730 8334
rect 28533 8331 28599 8334
rect 200 8258 800 8288
rect 1577 8258 1643 8261
rect 200 8256 1643 8258
rect 200 8200 1582 8256
rect 1638 8200 1643 8256
rect 200 8198 1643 8200
rect 200 8168 800 8198
rect 1577 8195 1643 8198
rect 36261 8258 36327 8261
rect 37200 8258 37800 8288
rect 36261 8256 37800 8258
rect 36261 8200 36266 8256
rect 36322 8200 37800 8256
rect 36261 8198 37800 8200
rect 36261 8195 36327 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 37200 8168 37800 8198
rect 34930 8127 35246 8128
rect 22093 8122 22159 8125
rect 28073 8122 28139 8125
rect 22093 8120 28139 8122
rect 22093 8064 22098 8120
rect 22154 8064 28078 8120
rect 28134 8064 28139 8120
rect 22093 8062 28139 8064
rect 22093 8059 22159 8062
rect 28073 8059 28139 8062
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 22737 7578 22803 7581
rect 27470 7578 27476 7580
rect 22737 7576 27476 7578
rect 22737 7520 22742 7576
rect 22798 7520 27476 7576
rect 22737 7518 27476 7520
rect 22737 7515 22803 7518
rect 27470 7516 27476 7518
rect 27540 7516 27546 7580
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 22001 6898 22067 6901
rect 26233 6898 26299 6901
rect 22001 6896 26299 6898
rect 22001 6840 22006 6896
rect 22062 6840 26238 6896
rect 26294 6840 26299 6896
rect 22001 6838 26299 6840
rect 22001 6835 22067 6838
rect 26233 6835 26299 6838
rect 35801 6898 35867 6901
rect 37200 6898 37800 6928
rect 35801 6896 37800 6898
rect 35801 6840 35806 6896
rect 35862 6840 37800 6896
rect 35801 6838 37800 6840
rect 35801 6835 35867 6838
rect 37200 6808 37800 6838
rect 23749 6762 23815 6765
rect 30741 6762 30807 6765
rect 23749 6760 30807 6762
rect 23749 6704 23754 6760
rect 23810 6704 30746 6760
rect 30802 6704 30807 6760
rect 23749 6702 30807 6704
rect 23749 6699 23815 6702
rect 30741 6699 30807 6702
rect 23933 6626 23999 6629
rect 26693 6626 26759 6629
rect 23933 6624 26759 6626
rect 23933 6568 23938 6624
rect 23994 6568 26698 6624
rect 26754 6568 26759 6624
rect 23933 6566 26759 6568
rect 23933 6563 23999 6566
rect 26693 6563 26759 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 13721 6354 13787 6357
rect 27797 6354 27863 6357
rect 13721 6352 27863 6354
rect 13721 6296 13726 6352
rect 13782 6296 27802 6352
rect 27858 6296 27863 6352
rect 13721 6294 27863 6296
rect 13721 6291 13787 6294
rect 27797 6291 27863 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 16297 5810 16363 5813
rect 24669 5810 24735 5813
rect 16297 5808 24735 5810
rect 16297 5752 16302 5808
rect 16358 5752 24674 5808
rect 24730 5752 24735 5808
rect 16297 5750 24735 5752
rect 16297 5747 16363 5750
rect 24669 5747 24735 5750
rect 25129 5810 25195 5813
rect 25957 5810 26023 5813
rect 25129 5808 26023 5810
rect 25129 5752 25134 5808
rect 25190 5752 25962 5808
rect 26018 5752 26023 5808
rect 25129 5750 26023 5752
rect 25129 5747 25195 5750
rect 25957 5747 26023 5750
rect 13629 5674 13695 5677
rect 23422 5674 23428 5676
rect 13629 5672 23428 5674
rect 13629 5616 13634 5672
rect 13690 5616 23428 5672
rect 13629 5614 23428 5616
rect 13629 5611 13695 5614
rect 23422 5612 23428 5614
rect 23492 5612 23498 5676
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 24393 5402 24459 5405
rect 28073 5402 28139 5405
rect 24393 5400 28139 5402
rect 24393 5344 24398 5400
rect 24454 5344 28078 5400
rect 28134 5344 28139 5400
rect 24393 5342 28139 5344
rect 24393 5339 24459 5342
rect 28073 5339 28139 5342
rect 16481 5266 16547 5269
rect 27654 5266 27660 5268
rect 16481 5264 27660 5266
rect 16481 5208 16486 5264
rect 16542 5208 27660 5264
rect 16481 5206 27660 5208
rect 16481 5203 16547 5206
rect 27654 5204 27660 5206
rect 27724 5204 27730 5268
rect 15561 5130 15627 5133
rect 27981 5130 28047 5133
rect 15561 5128 28047 5130
rect 15561 5072 15566 5128
rect 15622 5072 27986 5128
rect 28042 5072 28047 5128
rect 15561 5070 28047 5072
rect 15561 5067 15627 5070
rect 27981 5067 28047 5070
rect 22829 4994 22895 4997
rect 26233 4994 26299 4997
rect 22829 4992 26299 4994
rect 22829 4936 22834 4992
rect 22890 4936 26238 4992
rect 26294 4936 26299 4992
rect 22829 4934 26299 4936
rect 22829 4931 22895 4934
rect 26233 4931 26299 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1577 4858 1643 4861
rect 200 4856 1643 4858
rect 200 4800 1582 4856
rect 1638 4800 1643 4856
rect 200 4798 1643 4800
rect 200 4768 800 4798
rect 1577 4795 1643 4798
rect 13169 4858 13235 4861
rect 18781 4858 18847 4861
rect 13169 4856 18847 4858
rect 13169 4800 13174 4856
rect 13230 4800 18786 4856
rect 18842 4800 18847 4856
rect 13169 4798 18847 4800
rect 13169 4795 13235 4798
rect 18781 4795 18847 4798
rect 25078 4796 25084 4860
rect 25148 4858 25154 4860
rect 26693 4858 26759 4861
rect 25148 4856 26759 4858
rect 25148 4800 26698 4856
rect 26754 4800 26759 4856
rect 25148 4798 26759 4800
rect 25148 4796 25154 4798
rect 26693 4795 26759 4798
rect 36353 4858 36419 4861
rect 37200 4858 37800 4888
rect 36353 4856 37800 4858
rect 36353 4800 36358 4856
rect 36414 4800 37800 4856
rect 36353 4798 37800 4800
rect 36353 4795 36419 4798
rect 37200 4768 37800 4798
rect 12985 4722 13051 4725
rect 18229 4722 18295 4725
rect 12985 4720 18295 4722
rect 12985 4664 12990 4720
rect 13046 4664 18234 4720
rect 18290 4664 18295 4720
rect 12985 4662 18295 4664
rect 12985 4659 13051 4662
rect 18229 4659 18295 4662
rect 24301 4722 24367 4725
rect 25957 4722 26023 4725
rect 24301 4720 26023 4722
rect 24301 4664 24306 4720
rect 24362 4664 25962 4720
rect 26018 4664 26023 4720
rect 24301 4662 26023 4664
rect 24301 4659 24367 4662
rect 25957 4659 26023 4662
rect 19609 4586 19675 4589
rect 20989 4586 21055 4589
rect 19609 4584 21055 4586
rect 19609 4528 19614 4584
rect 19670 4528 20994 4584
rect 21050 4528 21055 4584
rect 19609 4526 21055 4528
rect 19609 4523 19675 4526
rect 20989 4523 21055 4526
rect 24117 4586 24183 4589
rect 24853 4586 24919 4589
rect 26969 4586 27035 4589
rect 24117 4584 27035 4586
rect 24117 4528 24122 4584
rect 24178 4528 24858 4584
rect 24914 4528 26974 4584
rect 27030 4528 27035 4584
rect 24117 4526 27035 4528
rect 24117 4523 24183 4526
rect 24853 4523 24919 4526
rect 26969 4523 27035 4526
rect 20437 4450 20503 4453
rect 25957 4450 26023 4453
rect 28717 4450 28783 4453
rect 20437 4448 28783 4450
rect 20437 4392 20442 4448
rect 20498 4392 25962 4448
rect 26018 4392 28722 4448
rect 28778 4392 28783 4448
rect 20437 4390 28783 4392
rect 20437 4387 20503 4390
rect 25957 4387 26023 4390
rect 28717 4387 28783 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 21909 4314 21975 4317
rect 26601 4314 26667 4317
rect 21909 4312 26667 4314
rect 21909 4256 21914 4312
rect 21970 4256 26606 4312
rect 26662 4256 26667 4312
rect 21909 4254 26667 4256
rect 21909 4251 21975 4254
rect 26601 4251 26667 4254
rect 18505 4178 18571 4181
rect 30373 4178 30439 4181
rect 18505 4176 30439 4178
rect 18505 4120 18510 4176
rect 18566 4120 30378 4176
rect 30434 4120 30439 4176
rect 18505 4118 30439 4120
rect 18505 4115 18571 4118
rect 30373 4115 30439 4118
rect 15142 3980 15148 4044
rect 15212 4042 15218 4044
rect 35893 4042 35959 4045
rect 15212 4040 35959 4042
rect 15212 3984 35898 4040
rect 35954 3984 35959 4040
rect 15212 3982 35959 3984
rect 15212 3980 15218 3982
rect 35893 3979 35959 3982
rect 23289 3906 23355 3909
rect 30741 3906 30807 3909
rect 23289 3904 30807 3906
rect 23289 3848 23294 3904
rect 23350 3848 30746 3904
rect 30802 3848 30807 3904
rect 23289 3846 30807 3848
rect 23289 3843 23355 3846
rect 30741 3843 30807 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 23381 3770 23447 3773
rect 28257 3770 28323 3773
rect 23381 3768 28323 3770
rect 23381 3712 23386 3768
rect 23442 3712 28262 3768
rect 28318 3712 28323 3768
rect 23381 3710 28323 3712
rect 23381 3707 23447 3710
rect 28257 3707 28323 3710
rect 13537 3634 13603 3637
rect 22461 3636 22527 3637
rect 22461 3634 22508 3636
rect 13537 3632 22508 3634
rect 22572 3634 22578 3636
rect 28993 3634 29059 3637
rect 22572 3632 29059 3634
rect 13537 3576 13542 3632
rect 13598 3576 22466 3632
rect 22572 3576 28998 3632
rect 29054 3576 29059 3632
rect 13537 3574 22508 3576
rect 13537 3571 13603 3574
rect 22461 3572 22508 3574
rect 22572 3574 29059 3576
rect 22572 3572 22578 3574
rect 22461 3571 22527 3572
rect 28993 3571 29059 3574
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 11789 3498 11855 3501
rect 14273 3498 14339 3501
rect 11789 3496 14339 3498
rect 11789 3440 11794 3496
rect 11850 3440 14278 3496
rect 14334 3440 14339 3496
rect 11789 3438 14339 3440
rect 11789 3435 11855 3438
rect 14273 3435 14339 3438
rect 18965 3498 19031 3501
rect 19333 3498 19399 3501
rect 18965 3496 19399 3498
rect 18965 3440 18970 3496
rect 19026 3440 19338 3496
rect 19394 3440 19399 3496
rect 18965 3438 19399 3440
rect 18965 3435 19031 3438
rect 19333 3435 19399 3438
rect 21725 3498 21791 3501
rect 25037 3498 25103 3501
rect 21725 3496 25103 3498
rect 21725 3440 21730 3496
rect 21786 3440 25042 3496
rect 25098 3440 25103 3496
rect 21725 3438 25103 3440
rect 21725 3435 21791 3438
rect 25037 3435 25103 3438
rect 36261 3498 36327 3501
rect 37200 3498 37800 3528
rect 36261 3496 37800 3498
rect 36261 3440 36266 3496
rect 36322 3440 37800 3496
rect 36261 3438 37800 3440
rect 36261 3435 36327 3438
rect 37200 3408 37800 3438
rect 21081 3362 21147 3365
rect 28441 3362 28507 3365
rect 21081 3360 28507 3362
rect 21081 3304 21086 3360
rect 21142 3304 28446 3360
rect 28502 3304 28507 3360
rect 21081 3302 28507 3304
rect 21081 3299 21147 3302
rect 28441 3299 28507 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 15009 3228 15075 3229
rect 14958 3164 14964 3228
rect 15028 3226 15075 3228
rect 15028 3224 15120 3226
rect 15070 3168 15120 3224
rect 15028 3166 15120 3168
rect 15028 3164 15075 3166
rect 15009 3163 15075 3164
rect 2405 3090 2471 3093
rect 18270 3090 18276 3092
rect 2405 3088 18276 3090
rect 2405 3032 2410 3088
rect 2466 3032 18276 3088
rect 2405 3030 18276 3032
rect 2405 3027 2471 3030
rect 18270 3028 18276 3030
rect 18340 3028 18346 3092
rect 18873 3090 18939 3093
rect 22185 3090 22251 3093
rect 18873 3088 22251 3090
rect 18873 3032 18878 3088
rect 18934 3032 22190 3088
rect 22246 3032 22251 3088
rect 18873 3030 22251 3032
rect 18873 3027 18939 3030
rect 22185 3027 22251 3030
rect 22461 3090 22527 3093
rect 26141 3090 26207 3093
rect 22461 3088 26207 3090
rect 22461 3032 22466 3088
rect 22522 3032 26146 3088
rect 26202 3032 26207 3088
rect 22461 3030 26207 3032
rect 22461 3027 22527 3030
rect 26141 3027 26207 3030
rect 27613 3090 27679 3093
rect 28993 3090 29059 3093
rect 27613 3088 29059 3090
rect 27613 3032 27618 3088
rect 27674 3032 28998 3088
rect 29054 3032 29059 3088
rect 27613 3030 29059 3032
rect 27613 3027 27679 3030
rect 28993 3027 29059 3030
rect 12065 2954 12131 2957
rect 12709 2954 12775 2957
rect 12065 2952 12775 2954
rect 12065 2896 12070 2952
rect 12126 2896 12714 2952
rect 12770 2896 12775 2952
rect 12065 2894 12775 2896
rect 12065 2891 12131 2894
rect 12709 2891 12775 2894
rect 13445 2954 13511 2957
rect 16573 2954 16639 2957
rect 13445 2952 16639 2954
rect 13445 2896 13450 2952
rect 13506 2896 16578 2952
rect 16634 2896 16639 2952
rect 13445 2894 16639 2896
rect 13445 2891 13511 2894
rect 16573 2891 16639 2894
rect 12433 2818 12499 2821
rect 14457 2818 14523 2821
rect 12433 2816 14523 2818
rect 12433 2760 12438 2816
rect 12494 2760 14462 2816
rect 14518 2760 14523 2816
rect 12433 2758 14523 2760
rect 12433 2755 12499 2758
rect 14457 2755 14523 2758
rect 24393 2818 24459 2821
rect 24669 2818 24735 2821
rect 27797 2818 27863 2821
rect 24393 2816 27863 2818
rect 24393 2760 24398 2816
rect 24454 2760 24674 2816
rect 24730 2760 27802 2816
rect 27858 2760 27863 2816
rect 24393 2758 27863 2760
rect 24393 2755 24459 2758
rect 24669 2755 24735 2758
rect 27797 2755 27863 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 13629 2682 13695 2685
rect 22134 2682 22140 2684
rect 13629 2680 22140 2682
rect 13629 2624 13634 2680
rect 13690 2624 22140 2680
rect 13629 2622 22140 2624
rect 13629 2619 13695 2622
rect 22134 2620 22140 2622
rect 22204 2620 22210 2684
rect 10869 2546 10935 2549
rect 21398 2546 21404 2548
rect 10869 2544 21404 2546
rect 10869 2488 10874 2544
rect 10930 2488 21404 2544
rect 10869 2486 21404 2488
rect 10869 2483 10935 2486
rect 21398 2484 21404 2486
rect 21468 2484 21474 2548
rect 10777 2410 10843 2413
rect 20846 2410 20852 2412
rect 10777 2408 20852 2410
rect 10777 2352 10782 2408
rect 10838 2352 20852 2408
rect 10777 2350 20852 2352
rect 10777 2347 10843 2350
rect 20846 2348 20852 2350
rect 20916 2348 20922 2412
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 2773 1458 2839 1461
rect 200 1456 2839 1458
rect 200 1400 2778 1456
rect 2834 1400 2839 1456
rect 200 1398 2839 1400
rect 200 1368 800 1398
rect 2773 1395 2839 1398
rect 36261 1458 36327 1461
rect 37200 1458 37800 1488
rect 36261 1456 37800 1458
rect 36261 1400 36266 1456
rect 36322 1400 37800 1456
rect 36261 1398 37800 1400
rect 36261 1395 36327 1398
rect 37200 1368 37800 1398
rect 35985 98 36051 101
rect 37200 98 37800 128
rect 35985 96 37800 98
rect 35985 40 35990 96
rect 36046 40 37800 96
rect 35985 38 37800 40
rect 35985 35 36051 38
rect 37200 8 37800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 15700 37088 15764 37092
rect 15700 37032 15714 37088
rect 15714 37032 15764 37088
rect 15700 37028 15764 37032
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 27476 36544 27540 36548
rect 27476 36488 27490 36544
rect 27490 36488 27540 36544
rect 27476 36484 27540 36488
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 25084 20844 25148 20908
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 20852 17640 20916 17644
rect 20852 17584 20866 17640
rect 20866 17584 20916 17640
rect 20852 17580 20916 17584
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 19380 16144 19444 16148
rect 19380 16088 19394 16144
rect 19394 16088 19444 16144
rect 19380 16084 19444 16088
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 21404 15676 21468 15740
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19380 14240 19444 14244
rect 19380 14184 19394 14240
rect 19394 14184 19444 14240
rect 19380 14180 19444 14184
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 22508 13636 22572 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 18276 12820 18340 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 15700 12140 15764 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 23428 11052 23492 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19380 10236 19444 10300
rect 14964 10100 15028 10164
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 15148 9692 15212 9756
rect 22140 9752 22204 9756
rect 22140 9696 22154 9752
rect 22154 9696 22204 9752
rect 22140 9692 22204 9696
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 27660 8332 27724 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 27476 7516 27540 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 23428 5612 23492 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 27660 5204 27724 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 25084 4796 25148 4860
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 15148 3980 15212 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 22508 3632 22572 3636
rect 22508 3576 22522 3632
rect 22522 3576 22572 3632
rect 22508 3572 22572 3576
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 14964 3224 15028 3228
rect 14964 3168 15014 3224
rect 15014 3168 15028 3224
rect 14964 3164 15028 3168
rect 18276 3028 18340 3092
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 22140 2620 22204 2684
rect 21404 2484 21468 2548
rect 20852 2348 20916 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 15699 37092 15765 37093
rect 15699 37028 15700 37092
rect 15764 37028 15765 37092
rect 15699 37027 15765 37028
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 15702 12205 15762 37027
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 27475 36548 27541 36549
rect 27475 36484 27476 36548
rect 27540 36484 27541 36548
rect 27475 36483 27541 36484
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 25083 20908 25149 20909
rect 25083 20844 25084 20908
rect 25148 20844 25149 20908
rect 25083 20843 25149 20844
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 20851 17644 20917 17645
rect 20851 17580 20852 17644
rect 20916 17580 20917 17644
rect 20851 17579 20917 17580
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19379 16148 19445 16149
rect 19379 16084 19380 16148
rect 19444 16084 19445 16148
rect 19379 16083 19445 16084
rect 19382 14245 19442 16083
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19379 14244 19445 14245
rect 19379 14180 19380 14244
rect 19444 14180 19445 14244
rect 19379 14179 19445 14180
rect 18275 12884 18341 12885
rect 18275 12820 18276 12884
rect 18340 12820 18341 12884
rect 18275 12819 18341 12820
rect 15699 12204 15765 12205
rect 15699 12140 15700 12204
rect 15764 12140 15765 12204
rect 15699 12139 15765 12140
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 14963 10164 15029 10165
rect 14963 10100 14964 10164
rect 15028 10100 15029 10164
rect 14963 10099 15029 10100
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 14966 3229 15026 10099
rect 15147 9756 15213 9757
rect 15147 9692 15148 9756
rect 15212 9692 15213 9756
rect 15147 9691 15213 9692
rect 15150 4045 15210 9691
rect 15147 4044 15213 4045
rect 15147 3980 15148 4044
rect 15212 3980 15213 4044
rect 15147 3979 15213 3980
rect 14963 3228 15029 3229
rect 14963 3164 14964 3228
rect 15028 3164 15029 3228
rect 14963 3163 15029 3164
rect 18278 3093 18338 12819
rect 19382 10301 19442 14179
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19379 10300 19445 10301
rect 19379 10236 19380 10300
rect 19444 10236 19445 10300
rect 19379 10235 19445 10236
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 18275 3092 18341 3093
rect 18275 3028 18276 3092
rect 18340 3028 18341 3092
rect 18275 3027 18341 3028
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 20854 2413 20914 17579
rect 21403 15740 21469 15741
rect 21403 15676 21404 15740
rect 21468 15676 21469 15740
rect 21403 15675 21469 15676
rect 21406 2549 21466 15675
rect 22507 13700 22573 13701
rect 22507 13636 22508 13700
rect 22572 13636 22573 13700
rect 22507 13635 22573 13636
rect 22139 9756 22205 9757
rect 22139 9692 22140 9756
rect 22204 9692 22205 9756
rect 22139 9691 22205 9692
rect 22142 2685 22202 9691
rect 22510 3637 22570 13635
rect 23427 11116 23493 11117
rect 23427 11052 23428 11116
rect 23492 11052 23493 11116
rect 23427 11051 23493 11052
rect 23430 5677 23490 11051
rect 23427 5676 23493 5677
rect 23427 5612 23428 5676
rect 23492 5612 23493 5676
rect 23427 5611 23493 5612
rect 25086 4861 25146 20843
rect 27478 7581 27538 36483
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 27659 8396 27725 8397
rect 27659 8332 27660 8396
rect 27724 8332 27725 8396
rect 27659 8331 27725 8332
rect 27475 7580 27541 7581
rect 27475 7516 27476 7580
rect 27540 7516 27541 7580
rect 27475 7515 27541 7516
rect 27662 5269 27722 8331
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 27659 5268 27725 5269
rect 27659 5204 27660 5268
rect 27724 5204 27725 5268
rect 27659 5203 27725 5204
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 25083 4860 25149 4861
rect 25083 4796 25084 4860
rect 25148 4796 25149 4860
rect 25083 4795 25149 4796
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 22507 3636 22573 3637
rect 22507 3572 22508 3636
rect 22572 3572 22573 3636
rect 22507 3571 22573 3572
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 22139 2684 22205 2685
rect 22139 2620 22140 2684
rect 22204 2620 22205 2684
rect 22139 2619 22205 2620
rect 21403 2548 21469 2549
rect 21403 2484 21404 2548
rect 21468 2484 21469 2548
rect 21403 2483 21469 2484
rect 20851 2412 20917 2413
rect 20851 2348 20852 2412
rect 20916 2348 20917 2412
rect 20851 2347 20917 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 9476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1667941163
transform 1 0 30360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1667941163
transform -1 0 9476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A
timestamp 1667941163
transform -1 0 32476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform -1 0 32200 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1667941163
transform 1 0 30912 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1667941163
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform 1 0 31464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1667941163
transform -1 0 31740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A
timestamp 1667941163
transform -1 0 9752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform -1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform 1 0 17940 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1667941163
transform -1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform -1 0 30452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 31648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1667941163
transform -1 0 28520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform -1 0 30452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform -1 0 31096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A
timestamp 1667941163
transform -1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform -1 0 10672 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform 1 0 14996 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1667941163
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1667941163
transform 1 0 22172 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1667941163
transform -1 0 20976 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1667941163
transform -1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform -1 0 28520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1667941163
transform -1 0 10120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1667941163
transform -1 0 10672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1667941163
transform 1 0 21344 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1667941163
transform -1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1667941163
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1667941163
transform -1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform -1 0 7360 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1667941163
transform -1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1667941163
transform -1 0 31004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1667941163
transform 1 0 26128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1667941163
transform -1 0 31556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform 1 0 9844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1667941163
transform -1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform -1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform -1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1667941163
transform -1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform -1 0 31096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1667941163
transform -1 0 27968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform 1 0 29716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform -1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform 1 0 20240 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1667941163
transform -1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1667941163
transform -1 0 30544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform -1 0 23276 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1667941163
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform -1 0 21252 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform -1 0 19596 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform -1 0 27968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1667941163
transform -1 0 26128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1667941163
transform -1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1667941163
transform 1 0 16560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1667941163
transform -1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1667941163
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1667941163
transform -1 0 30452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1667941163
transform -1 0 13984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1667941163
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1667941163
transform -1 0 30544 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1667941163
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1667941163
transform 1 0 28888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1667941163
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1667941163
transform -1 0 30636 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1667941163
transform -1 0 29900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1667941163
transform 1 0 10672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1667941163
transform -1 0 24564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1667941163
transform 1 0 25576 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1667941163
transform 1 0 31556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1667941163
transform -1 0 17848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1667941163
transform 1 0 8280 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1667941163
transform -1 0 27968 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1667941163
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1667941163
transform 1 0 23092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1667941163
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A
timestamp 1667941163
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1667941163
transform -1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1667941163
transform 1 0 8004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1667941163
transform 1 0 9476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1667941163
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1667941163
transform 1 0 31464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1667941163
transform 1 0 9936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1667941163
transform 1 0 31556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A
timestamp 1667941163
transform -1 0 8280 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1667941163
transform -1 0 35696 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1667941163
transform -1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__A
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__A
timestamp 1667941163
transform 1 0 21160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__A
timestamp 1667941163
transform 1 0 18676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1667941163
transform -1 0 9476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1667941163
transform -1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__A
timestamp 1667941163
transform 1 0 23920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A
timestamp 1667941163
transform 1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1667941163
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A
timestamp 1667941163
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__D
timestamp 1667941163
transform -1 0 23276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__D
timestamp 1667941163
transform -1 0 14536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__D
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__D
timestamp 1667941163
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__D
timestamp 1667941163
transform -1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__D
timestamp 1667941163
transform -1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__D
timestamp 1667941163
transform -1 0 26956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__RESET_B
timestamp 1667941163
transform -1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__D
timestamp 1667941163
transform -1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__D
timestamp 1667941163
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__D
timestamp 1667941163
transform -1 0 29164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__D
timestamp 1667941163
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__RESET_B
timestamp 1667941163
transform -1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__D
timestamp 1667941163
transform 1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__D
timestamp 1667941163
transform -1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__D
timestamp 1667941163
transform -1 0 28980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__D
timestamp 1667941163
transform -1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__D
timestamp 1667941163
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__D
timestamp 1667941163
transform -1 0 19688 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__D
timestamp 1667941163
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__D
timestamp 1667941163
transform -1 0 17480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__D
timestamp 1667941163
transform -1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__D
timestamp 1667941163
transform -1 0 26956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__D
timestamp 1667941163
transform -1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__D
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__D
timestamp 1667941163
transform -1 0 28980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__D
timestamp 1667941163
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__D
timestamp 1667941163
transform -1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__D
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__D
timestamp 1667941163
transform 1 0 28244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__RESET_B
timestamp 1667941163
transform -1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__RESET_B
timestamp 1667941163
transform -1 0 11592 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__D
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__RESET_B
timestamp 1667941163
transform -1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__A
timestamp 1667941163
transform -1 0 30084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__A
timestamp 1667941163
transform -1 0 24748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__A
timestamp 1667941163
transform -1 0 27968 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__A
timestamp 1667941163
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__A
timestamp 1667941163
transform -1 0 29900 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__A
timestamp 1667941163
transform 1 0 2392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__A
timestamp 1667941163
transform 1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__A
timestamp 1667941163
transform 1 0 9936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__A
timestamp 1667941163
transform 1 0 30912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__A
timestamp 1667941163
transform -1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__A
timestamp 1667941163
transform -1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__A
timestamp 1667941163
transform -1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__A
timestamp 1667941163
transform -1 0 30820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__A
timestamp 1667941163
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A
timestamp 1667941163
transform 1 0 20424 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__A
timestamp 1667941163
transform -1 0 22816 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__A
timestamp 1667941163
transform 1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__A
timestamp 1667941163
transform 1 0 26496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__A
timestamp 1667941163
transform -1 0 21620 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__A
timestamp 1667941163
transform 1 0 12696 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__A
timestamp 1667941163
transform 1 0 31648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1667941163
transform -1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__A
timestamp 1667941163
transform -1 0 21988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A
timestamp 1667941163
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__A
timestamp 1667941163
transform -1 0 33120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A
timestamp 1667941163
transform -1 0 10028 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A
timestamp 1667941163
transform -1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__A
timestamp 1667941163
transform 1 0 27784 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A
timestamp 1667941163
transform -1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__A
timestamp 1667941163
transform 1 0 31188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1667941163
transform 1 0 9844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__744__A
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__759__A
timestamp 1667941163
transform 1 0 32016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__765__A
timestamp 1667941163
transform 1 0 22172 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1667941163
transform 1 0 20424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_prog_clk_A
timestamp 1667941163
transform -1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_prog_clk_A
timestamp 1667941163
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_prog_clk_A
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_prog_clk_A
timestamp 1667941163
transform -1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_prog_clk_A
timestamp 1667941163
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_prog_clk_A
timestamp 1667941163
transform -1 0 30636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_prog_clk_A
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_prog_clk_A
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform 1 0 26496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 12604 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform 1 0 16192 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 35696 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 35696 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 19412 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 36432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 35144 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 36432 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 1748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 1748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 32476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 36432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 35052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 1748 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 1748 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 33764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 35788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 35696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 27508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 1748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 34500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 35696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 1748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 4232 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 35788 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1667941163
transform 1 0 35512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1667941163
transform -1 0 15824 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1667941163
transform 1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform 1 0 18492 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1667941163
transform 1 0 2300 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1667941163
transform 1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1667941163
transform -1 0 2484 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1667941163
transform -1 0 34960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1667941163
transform 1 0 35880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1667941163
transform -1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1667941163
transform 1 0 3496 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1667941163
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1667941163
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1667941163
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1667941163
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1667941163
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1667941163
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_341
timestamp 1667941163
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1667941163
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_356
timestamp 1667941163
transform 1 0 33856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1667941163
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_384
timestamp 1667941163
transform 1 0 36432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3128 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1667941163
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1667941163
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1667941163
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1667941163
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1667941163
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_138
timestamp 1667941163
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_144
timestamp 1667941163
transform 1 0 14352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1667941163
transform 1 0 17204 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp 1667941163
transform 1 0 17940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1667941163
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1667941163
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1667941163
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1667941163
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_303
timestamp 1667941163
transform 1 0 28980 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_321
timestamp 1667941163
transform 1 0 30636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_328
timestamp 1667941163
transform 1 0 31280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_355
timestamp 1667941163
transform 1 0 33764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1667941163
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_369
timestamp 1667941163
transform 1 0 35052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_376
timestamp 1667941163
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1667941163
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1667941163
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1667941163
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_154
timestamp 1667941163
transform 1 0 15272 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1667941163
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1667941163
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1667941163
transform 1 0 21804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1667941163
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1667941163
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_299
timestamp 1667941163
transform 1 0 28612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1667941163
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1667941163
transform 1 0 30084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_327
timestamp 1667941163
transform 1 0 31188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1667941163
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 1667941163
transform 1 0 32200 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_372
timestamp 1667941163
transform 1 0 35328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_384
timestamp 1667941163
transform 1 0 36432 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1667941163
transform 1 0 9476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1667941163
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1667941163
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1667941163
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_138
timestamp 1667941163
transform 1 0 13800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1667941163
transform 1 0 18676 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1667941163
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_303
timestamp 1667941163
transform 1 0 28980 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1667941163
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_315
timestamp 1667941163
transform 1 0 30084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1667941163
transform 1 0 30820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1667941163
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_377
timestamp 1667941163
transform 1 0 35788 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_380
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_89
timestamp 1667941163
transform 1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1667941163
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1667941163
transform 1 0 10488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_108
timestamp 1667941163
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1667941163
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1667941163
transform 1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1667941163
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1667941163
transform 1 0 18308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_191
timestamp 1667941163
transform 1 0 18676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1667941163
transform 1 0 19596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_222
timestamp 1667941163
transform 1 0 21528 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1667941163
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_283
timestamp 1667941163
transform 1 0 27140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1667941163
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_297
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1667941163
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_325
timestamp 1667941163
transform 1 0 31004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1667941163
transform 1 0 32108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1667941163
transform 1 0 33212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1667941163
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_381
timestamp 1667941163
transform 1 0 36156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_384
timestamp 1667941163
transform 1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_89
timestamp 1667941163
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_101
timestamp 1667941163
transform 1 0 10396 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_107
timestamp 1667941163
transform 1 0 10948 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1667941163
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1667941163
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_177
timestamp 1667941163
transform 1 0 17388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_183
timestamp 1667941163
transform 1 0 17940 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_186
timestamp 1667941163
transform 1 0 18216 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_247
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1667941163
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_285
timestamp 1667941163
transform 1 0 27324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_291
timestamp 1667941163
transform 1 0 27876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_299
timestamp 1667941163
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_384
timestamp 1667941163
transform 1 0 36432 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_90
timestamp 1667941163
transform 1 0 9384 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_102
timestamp 1667941163
transform 1 0 10488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_110
timestamp 1667941163
transform 1 0 11224 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1667941163
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1667941163
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_151
timestamp 1667941163
transform 1 0 14996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1667941163
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_184
timestamp 1667941163
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1667941163
transform 1 0 18308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1667941163
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_201
timestamp 1667941163
transform 1 0 19596 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1667941163
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_239
timestamp 1667941163
transform 1 0 23092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1667941163
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_275
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_281
timestamp 1667941163
transform 1 0 26956 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_287
timestamp 1667941163
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1667941163
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_315
timestamp 1667941163
transform 1 0 30084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_327
timestamp 1667941163
transform 1 0 31188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_331
timestamp 1667941163
transform 1 0 31556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_335
timestamp 1667941163
transform 1 0 31924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_347
timestamp 1667941163
transform 1 0 33028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1667941163
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_385
timestamp 1667941163
transform 1 0 36524 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_76
timestamp 1667941163
transform 1 0 8096 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_82
timestamp 1667941163
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_94
timestamp 1667941163
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_97
timestamp 1667941163
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1667941163
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1667941163
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1667941163
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_173
timestamp 1667941163
transform 1 0 17020 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_197
timestamp 1667941163
transform 1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1667941163
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_250
timestamp 1667941163
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_254
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_285
timestamp 1667941163
transform 1 0 27324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_292
timestamp 1667941163
transform 1 0 27968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_300
timestamp 1667941163
transform 1 0 28704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_312
timestamp 1667941163
transform 1 0 29808 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_319
timestamp 1667941163
transform 1 0 30452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 1667941163
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_104
timestamp 1667941163
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_110
timestamp 1667941163
transform 1 0 11224 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1667941163
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1667941163
transform 1 0 17020 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_179
timestamp 1667941163
transform 1 0 17572 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_231
timestamp 1667941163
transform 1 0 22356 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1667941163
transform 1 0 23276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_275
timestamp 1667941163
transform 1 0 26404 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_281
timestamp 1667941163
transform 1 0 26956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1667941163
transform 1 0 27600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1667941163
transform 1 0 28244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1667941163
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_314
timestamp 1667941163
transform 1 0 29992 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_326
timestamp 1667941163
transform 1 0 31096 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_338
timestamp 1667941163
transform 1 0 32200 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_347
timestamp 1667941163
transform 1 0 33028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1667941163
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 1667941163
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_117
timestamp 1667941163
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1667941163
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1667941163
transform 1 0 14168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1667941163
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1667941163
transform 1 0 17848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_185
timestamp 1667941163
transform 1 0 18124 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_191
timestamp 1667941163
transform 1 0 18676 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_213
timestamp 1667941163
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1667941163
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1667941163
transform 1 0 22172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1667941163
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_241
timestamp 1667941163
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_268
timestamp 1667941163
transform 1 0 25760 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_274
timestamp 1667941163
transform 1 0 26312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_300
timestamp 1667941163
transform 1 0 28704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_307
timestamp 1667941163
transform 1 0 29348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_314
timestamp 1667941163
transform 1 0 29992 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1667941163
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1667941163
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_376
timestamp 1667941163
transform 1 0 35696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_384
timestamp 1667941163
transform 1 0 36432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_7
timestamp 1667941163
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1667941163
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_60
timestamp 1667941163
transform 1 0 6624 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_66
timestamp 1667941163
transform 1 0 7176 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1667941163
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1667941163
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_117
timestamp 1667941163
transform 1 0 11868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1667941163
transform 1 0 14536 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_175
timestamp 1667941163
transform 1 0 17204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_184
timestamp 1667941163
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_222
timestamp 1667941163
transform 1 0 21528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_246
timestamp 1667941163
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_276
timestamp 1667941163
transform 1 0 26496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_284
timestamp 1667941163
transform 1 0 27232 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_288
timestamp 1667941163
transform 1 0 27600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_294
timestamp 1667941163
transform 1 0 28152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_298
timestamp 1667941163
transform 1 0 28520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1667941163
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_318
timestamp 1667941163
transform 1 0 30360 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_330
timestamp 1667941163
transform 1 0 31464 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_342
timestamp 1667941163
transform 1 0 32568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_354
timestamp 1667941163
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1667941163
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_385
timestamp 1667941163
transform 1 0 36524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1667941163
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1667941163
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1667941163
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1667941163
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1667941163
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1667941163
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1667941163
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_120
timestamp 1667941163
transform 1 0 12144 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_128
timestamp 1667941163
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1667941163
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1667941163
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_173
timestamp 1667941163
transform 1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1667941163
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1667941163
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_214
timestamp 1667941163
transform 1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1667941163
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_231
timestamp 1667941163
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_260
timestamp 1667941163
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_266
timestamp 1667941163
transform 1 0 25576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1667941163
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_287
timestamp 1667941163
transform 1 0 27508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_297
timestamp 1667941163
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_303
timestamp 1667941163
transform 1 0 28980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1667941163
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_323
timestamp 1667941163
transform 1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1667941163
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_379
timestamp 1667941163
transform 1 0 35972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 1667941163
transform 1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp 1667941163
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_104
timestamp 1667941163
transform 1 0 10672 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1667941163
transform 1 0 11224 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1667941163
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1667941163
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1667941163
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1667941163
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1667941163
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1667941163
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_244
timestamp 1667941163
transform 1 0 23552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1667941163
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_278
timestamp 1667941163
transform 1 0 26680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1667941163
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_317
timestamp 1667941163
transform 1 0 30268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_324
timestamp 1667941163
transform 1 0 30912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_328
timestamp 1667941163
transform 1 0 31280 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_350
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1667941163
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_385
timestamp 1667941163
transform 1 0 36524 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1667941163
transform 1 0 9476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1667941163
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_124
timestamp 1667941163
transform 1 0 12512 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_130
timestamp 1667941163
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_134
timestamp 1667941163
transform 1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1667941163
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_173
timestamp 1667941163
transform 1 0 17020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_200
timestamp 1667941163
transform 1 0 19504 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1667941163
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1667941163
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 1667941163
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_255
timestamp 1667941163
transform 1 0 24564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1667941163
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1667941163
transform 1 0 28704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_307
timestamp 1667941163
transform 1 0 29348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_313
timestamp 1667941163
transform 1 0 29900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_323
timestamp 1667941163
transform 1 0 30820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_377
timestamp 1667941163
transform 1 0 35788 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_381
timestamp 1667941163
transform 1 0 36156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1667941163
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_96
timestamp 1667941163
transform 1 0 9936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1667941163
transform 1 0 10488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1667941163
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1667941163
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1667941163
transform 1 0 12512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1667941163
transform 1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1667941163
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_175
timestamp 1667941163
transform 1 0 17204 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_183
timestamp 1667941163
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1667941163
transform 1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1667941163
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1667941163
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_241
timestamp 1667941163
transform 1 0 23276 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1667941163
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_278
timestamp 1667941163
transform 1 0 26680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_285
timestamp 1667941163
transform 1 0 27324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_292
timestamp 1667941163
transform 1 0 27968 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1667941163
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 1667941163
transform 1 0 30544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1667941163
transform 1 0 31188 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_385
timestamp 1667941163
transform 1 0 36524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1667941163
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1667941163
transform 1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_91
timestamp 1667941163
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1667941163
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1667941163
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_124
timestamp 1667941163
transform 1 0 12512 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1667941163
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1667941163
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1667941163
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1667941163
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1667941163
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1667941163
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_263
timestamp 1667941163
transform 1 0 25300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_270
timestamp 1667941163
transform 1 0 25944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1667941163
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_292
timestamp 1667941163
transform 1 0 27968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_302
timestamp 1667941163
transform 1 0 28888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1667941163
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1667941163
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_326
timestamp 1667941163
transform 1 0 31096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1667941163
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1667941163
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_384
timestamp 1667941163
transform 1 0 36432 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1667941163
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1667941163
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_113
timestamp 1667941163
transform 1 0 11500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_119
timestamp 1667941163
transform 1 0 12052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1667941163
transform 1 0 12420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1667941163
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1667941163
transform 1 0 14720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1667941163
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1667941163
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_222
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1667941163
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1667941163
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_243
timestamp 1667941163
transform 1 0 23460 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_272
timestamp 1667941163
transform 1 0 26128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_279
timestamp 1667941163
transform 1 0 26772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_286
timestamp 1667941163
transform 1 0 27416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_300
timestamp 1667941163
transform 1 0 28704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_320
timestamp 1667941163
transform 1 0 30544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_326
timestamp 1667941163
transform 1 0 31096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1667941163
transform 1 0 31648 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1667941163
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1667941163
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1667941163
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_385
timestamp 1667941163
transform 1 0 36524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_21
timestamp 1667941163
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_33
timestamp 1667941163
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1667941163
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1667941163
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1667941163
transform 1 0 8188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_83
timestamp 1667941163
transform 1 0 8740 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_124
timestamp 1667941163
transform 1 0 12512 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_139
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_154
timestamp 1667941163
transform 1 0 15272 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_162
timestamp 1667941163
transform 1 0 16008 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1667941163
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_183
timestamp 1667941163
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1667941163
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_197
timestamp 1667941163
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_203
timestamp 1667941163
transform 1 0 19780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1667941163
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1667941163
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_236
timestamp 1667941163
transform 1 0 22816 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_257
timestamp 1667941163
transform 1 0 24748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_264
timestamp 1667941163
transform 1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_271
timestamp 1667941163
transform 1 0 26036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1667941163
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1667941163
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_314
timestamp 1667941163
transform 1 0 29992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_320
timestamp 1667941163
transform 1 0 30544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_326
timestamp 1667941163
transform 1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1667941163
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_376
timestamp 1667941163
transform 1 0 35696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_384
timestamp 1667941163
transform 1 0 36432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_10
timestamp 1667941163
transform 1 0 2024 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1667941163
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1667941163
transform 1 0 7360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1667941163
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_92
timestamp 1667941163
transform 1 0 9568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1667941163
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1667941163
transform 1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_113
timestamp 1667941163
transform 1 0 11500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1667941163
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1667941163
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_155
timestamp 1667941163
transform 1 0 15364 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_161
timestamp 1667941163
transform 1 0 15916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_171
timestamp 1667941163
transform 1 0 16836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_184
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_190
timestamp 1667941163
transform 1 0 18584 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_217
timestamp 1667941163
transform 1 0 21068 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_227
timestamp 1667941163
transform 1 0 21988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1667941163
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1667941163
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_279
timestamp 1667941163
transform 1 0 26772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1667941163
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_326
timestamp 1667941163
transform 1 0 31096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_332
timestamp 1667941163
transform 1 0 31648 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_338
timestamp 1667941163
transform 1 0 32200 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_350
timestamp 1667941163
transform 1 0 33304 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1667941163
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_385
timestamp 1667941163
transform 1 0 36524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1667941163
transform 1 0 2392 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_20
timestamp 1667941163
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_32
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_44
timestamp 1667941163
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1667941163
transform 1 0 8188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1667941163
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1667941163
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1667941163
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1667941163
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1667941163
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1667941163
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1667941163
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1667941163
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_189
timestamp 1667941163
transform 1 0 18492 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_195
timestamp 1667941163
transform 1 0 19044 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_199
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1667941163
transform 1 0 20884 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_238
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1667941163
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_252
timestamp 1667941163
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_259
timestamp 1667941163
transform 1 0 24932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_263
timestamp 1667941163
transform 1 0 25300 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1667941163
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1667941163
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_307
timestamp 1667941163
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_314
timestamp 1667941163
transform 1 0 29992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_321
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_328
timestamp 1667941163
transform 1 0 31280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1667941163
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_341
timestamp 1667941163
transform 1 0 32476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_353
timestamp 1667941163
transform 1 0 33580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_365
timestamp 1667941163
transform 1 0 34684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_377
timestamp 1667941163
transform 1 0 35788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1667941163
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_90
timestamp 1667941163
transform 1 0 9384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_110
timestamp 1667941163
transform 1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_123
timestamp 1667941163
transform 1 0 12420 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_152
timestamp 1667941163
transform 1 0 15088 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1667941163
transform 1 0 16468 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_188
timestamp 1667941163
transform 1 0 18400 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_212
timestamp 1667941163
transform 1 0 20608 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_225
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_238
timestamp 1667941163
transform 1 0 23000 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1667941163
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1667941163
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_299
timestamp 1667941163
transform 1 0 28612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1667941163
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_327
timestamp 1667941163
transform 1 0 31188 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_385
timestamp 1667941163
transform 1 0 36524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_77
timestamp 1667941163
transform 1 0 8188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_88
timestamp 1667941163
transform 1 0 9200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_94
timestamp 1667941163
transform 1 0 9752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_101
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_119
timestamp 1667941163
transform 1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1667941163
transform 1 0 13248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1667941163
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1667941163
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_214
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_218
timestamp 1667941163
transform 1 0 21160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_241
timestamp 1667941163
transform 1 0 23276 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_255
timestamp 1667941163
transform 1 0 24564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_268
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1667941163
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_292
timestamp 1667941163
transform 1 0 27968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_312
timestamp 1667941163
transform 1 0 29808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_319
timestamp 1667941163
transform 1 0 30452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_325
timestamp 1667941163
transform 1 0 31004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1667941163
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_377
timestamp 1667941163
transform 1 0 35788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_384
timestamp 1667941163
transform 1 0 36432 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1667941163
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_92
timestamp 1667941163
transform 1 0 9568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_98
timestamp 1667941163
transform 1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_104
timestamp 1667941163
transform 1 0 10672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1667941163
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1667941163
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1667941163
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_151
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1667941163
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_201
timestamp 1667941163
transform 1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_214
timestamp 1667941163
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_229
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_243
timestamp 1667941163
transform 1 0 23460 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_268
timestamp 1667941163
transform 1 0 25760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_294
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1667941163
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_385
timestamp 1667941163
transform 1 0 36524 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1667941163
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_104
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1667941163
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 1667941163
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_155
timestamp 1667941163
transform 1 0 15364 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1667941163
transform 1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1667941163
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1667941163
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1667941163
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_262
timestamp 1667941163
transform 1 0 25208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1667941163
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_285
timestamp 1667941163
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1667941163
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_307
timestamp 1667941163
transform 1 0 29348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1667941163
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1667941163
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_377
timestamp 1667941163
transform 1 0 35788 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_382
timestamp 1667941163
transform 1 0 36248 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_40
timestamp 1667941163
transform 1 0 4784 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_52
timestamp 1667941163
transform 1 0 5888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_64
timestamp 1667941163
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1667941163
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1667941163
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1667941163
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1667941163
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1667941163
transform 1 0 11868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_146
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1667941163
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1667941163
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_203
timestamp 1667941163
transform 1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_210
timestamp 1667941163
transform 1 0 20424 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1667941163
transform 1 0 20976 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1667941163
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1667941163
transform 1 0 23092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1667941163
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_264
timestamp 1667941163
transform 1 0 25392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_290
timestamp 1667941163
transform 1 0 27784 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1667941163
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_328
timestamp 1667941163
transform 1 0 31280 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_340
timestamp 1667941163
transform 1 0 32384 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_352
timestamp 1667941163
transform 1 0 33488 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_385
timestamp 1667941163
transform 1 0 36524 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_16
timestamp 1667941163
transform 1 0 2576 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_22
timestamp 1667941163
transform 1 0 3128 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_34
timestamp 1667941163
transform 1 0 4232 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_46
timestamp 1667941163
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_101
timestamp 1667941163
transform 1 0 10396 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_104
timestamp 1667941163
transform 1 0 10672 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 1667941163
transform 1 0 12696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_133
timestamp 1667941163
transform 1 0 13340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_151
timestamp 1667941163
transform 1 0 14996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_188
timestamp 1667941163
transform 1 0 18400 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_210
timestamp 1667941163
transform 1 0 20424 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_214
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_241
timestamp 1667941163
transform 1 0 23276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_262
timestamp 1667941163
transform 1 0 25208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_290
timestamp 1667941163
transform 1 0 27784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_299
timestamp 1667941163
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_313
timestamp 1667941163
transform 1 0 29900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_319
timestamp 1667941163
transform 1 0 30452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_325
timestamp 1667941163
transform 1 0 31004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_379
timestamp 1667941163
transform 1 0 35972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_384
timestamp 1667941163
transform 1 0 36432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_7
timestamp 1667941163
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1667941163
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1667941163
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1667941163
transform 1 0 12052 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1667941163
transform 1 0 12696 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1667941163
transform 1 0 14536 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1667941163
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_172
timestamp 1667941163
transform 1 0 16928 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_183
timestamp 1667941163
transform 1 0 17940 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1667941163
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_228
timestamp 1667941163
transform 1 0 22080 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1667941163
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1667941163
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1667941163
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1667941163
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_297
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1667941163
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_313
timestamp 1667941163
transform 1 0 29900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_319
timestamp 1667941163
transform 1 0 30452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_323
timestamp 1667941163
transform 1 0 30820 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_326
timestamp 1667941163
transform 1 0 31096 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_338
timestamp 1667941163
transform 1 0 32200 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_350
timestamp 1667941163
transform 1 0 33304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1667941163
transform 1 0 36524 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1667941163
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1667941163
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1667941163
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1667941163
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1667941163
transform 1 0 9568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_98
timestamp 1667941163
transform 1 0 10120 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1667941163
transform 1 0 10856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 1667941163
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1667941163
transform 1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1667941163
transform 1 0 13524 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1667941163
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1667941163
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1667941163
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_200
timestamp 1667941163
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_208
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1667941163
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1667941163
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1667941163
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_266
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1667941163
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_307
timestamp 1667941163
transform 1 0 29348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_313
timestamp 1667941163
transform 1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1667941163
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_379
timestamp 1667941163
transform 1 0 35972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_384
timestamp 1667941163
transform 1 0 36432 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_103
timestamp 1667941163
transform 1 0 10580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1667941163
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_113
timestamp 1667941163
transform 1 0 11500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_124
timestamp 1667941163
transform 1 0 12512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1667941163
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1667941163
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1667941163
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_185
timestamp 1667941163
transform 1 0 18124 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1667941163
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1667941163
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_228
timestamp 1667941163
transform 1 0 22080 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1667941163
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_268
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_274
timestamp 1667941163
transform 1 0 26312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_291
timestamp 1667941163
transform 1 0 27876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1667941163
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_313
timestamp 1667941163
transform 1 0 29900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_325
timestamp 1667941163
transform 1 0 31004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_337
timestamp 1667941163
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_349
timestamp 1667941163
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1667941163
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1667941163
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1667941163
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_134
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1667941163
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_175
timestamp 1667941163
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1667941163
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1667941163
transform 1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1667941163
transform 1 0 19412 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1667941163
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_231
timestamp 1667941163
transform 1 0 22356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1667941163
transform 1 0 23644 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1667941163
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1667941163
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_263
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1667941163
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_304
timestamp 1667941163
transform 1 0 29072 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_316
timestamp 1667941163
transform 1 0 30176 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1667941163
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_7
timestamp 1667941163
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1667941163
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_150
timestamp 1667941163
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1667941163
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_161
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_172
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_180
timestamp 1667941163
transform 1 0 17664 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_201
timestamp 1667941163
transform 1 0 19596 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_210
timestamp 1667941163
transform 1 0 20424 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_216
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1667941163
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_230
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_234
timestamp 1667941163
transform 1 0 22632 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_238
timestamp 1667941163
transform 1 0 23000 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1667941163
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1667941163
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_262
timestamp 1667941163
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_279
timestamp 1667941163
transform 1 0 26772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_286
timestamp 1667941163
transform 1 0 27416 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1667941163
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1667941163
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1667941163
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1667941163
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1667941163
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1667941163
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1667941163
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_183
timestamp 1667941163
transform 1 0 17940 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_200
timestamp 1667941163
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_206
timestamp 1667941163
transform 1 0 20056 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_216
timestamp 1667941163
transform 1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1667941163
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1667941163
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_269
timestamp 1667941163
transform 1 0 25852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1667941163
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_292
timestamp 1667941163
transform 1 0 27968 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_304
timestamp 1667941163
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1667941163
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_342
timestamp 1667941163
transform 1 0 32568 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_348
timestamp 1667941163
transform 1 0 33120 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_360
timestamp 1667941163
transform 1 0 34224 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_372
timestamp 1667941163
transform 1 0 35328 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_384
timestamp 1667941163
transform 1 0 36432 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1667941163
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1667941163
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1667941163
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_182
timestamp 1667941163
transform 1 0 17848 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_188
timestamp 1667941163
transform 1 0 18400 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_203
timestamp 1667941163
transform 1 0 19780 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1667941163
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_216
timestamp 1667941163
transform 1 0 20976 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1667941163
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_227
timestamp 1667941163
transform 1 0 21988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 1667941163
transform 1 0 22356 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_244
timestamp 1667941163
transform 1 0 23552 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_264
timestamp 1667941163
transform 1 0 25392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_290
timestamp 1667941163
transform 1 0 27784 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1667941163
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_385
timestamp 1667941163
transform 1 0 36524 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_10
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_16
timestamp 1667941163
transform 1 0 2576 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_28
timestamp 1667941163
transform 1 0 3680 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_40
timestamp 1667941163
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1667941163
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_152
timestamp 1667941163
transform 1 0 15088 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1667941163
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1667941163
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1667941163
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1667941163
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1667941163
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1667941163
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_245
timestamp 1667941163
transform 1 0 23644 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_253
timestamp 1667941163
transform 1 0 24380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_258
timestamp 1667941163
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1667941163
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1667941163
transform 1 0 26128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_316
timestamp 1667941163
transform 1 0 30176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1667941163
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp 1667941163
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_186
timestamp 1667941163
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1667941163
transform 1 0 20700 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_223
timestamp 1667941163
transform 1 0 21620 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_231
timestamp 1667941163
transform 1 0 22356 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1667941163
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1667941163
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1667941163
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_266
timestamp 1667941163
transform 1 0 25576 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_272
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_284
timestamp 1667941163
transform 1 0 27232 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_296
timestamp 1667941163
transform 1 0 28336 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_384
timestamp 1667941163
transform 1 0 36432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1667941163
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_19
timestamp 1667941163
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1667941163
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 1667941163
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1667941163
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1667941163
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_231
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_238
timestamp 1667941163
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1667941163
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_251
timestamp 1667941163
transform 1 0 24196 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_259
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_262
timestamp 1667941163
transform 1 0 25208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1667941163
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_158
timestamp 1667941163
transform 1 0 15640 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_170
timestamp 1667941163
transform 1 0 16744 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_182
timestamp 1667941163
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_212
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_224
timestamp 1667941163
transform 1 0 21712 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_239
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_385
timestamp 1667941163
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1667941163
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1667941163
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1667941163
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_214
timestamp 1667941163
transform 1 0 20792 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_229
timestamp 1667941163
transform 1 0 22172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_241
timestamp 1667941163
transform 1 0 23276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_253
timestamp 1667941163
transform 1 0 24380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_265
timestamp 1667941163
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1667941163
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1667941163
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_292
timestamp 1667941163
transform 1 0 27968 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_304
timestamp 1667941163
transform 1 0 29072 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_316
timestamp 1667941163
transform 1 0 30176 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_328
timestamp 1667941163
transform 1 0 31280 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_379
timestamp 1667941163
transform 1 0 35972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_384
timestamp 1667941163
transform 1 0 36432 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_201
timestamp 1667941163
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_208
timestamp 1667941163
transform 1 0 20240 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_223
timestamp 1667941163
transform 1 0 21620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_235
timestamp 1667941163
transform 1 0 22724 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1667941163
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_385
timestamp 1667941163
transform 1 0 36524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_7
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_19
timestamp 1667941163
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_31
timestamp 1667941163
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_43
timestamp 1667941163
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_245
timestamp 1667941163
transform 1 0 23644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_255
timestamp 1667941163
transform 1 0 24564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_267
timestamp 1667941163
transform 1 0 25668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_373
timestamp 1667941163
transform 1 0 35420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_384
timestamp 1667941163
transform 1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_267
timestamp 1667941163
transform 1 0 25668 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_272
timestamp 1667941163
transform 1 0 26128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_385
timestamp 1667941163
transform 1 0 36524 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_262
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_268
timestamp 1667941163
transform 1 0 25760 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_280
timestamp 1667941163
transform 1 0 26864 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_292
timestamp 1667941163
transform 1 0 27968 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1667941163
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_384
timestamp 1667941163
transform 1 0 36432 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_72
timestamp 1667941163
transform 1 0 7728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1667941163
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_120
timestamp 1667941163
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1667941163
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_314
timestamp 1667941163
transform 1 0 29992 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_326
timestamp 1667941163
transform 1 0 31096 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_338
timestamp 1667941163
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_350
timestamp 1667941163
transform 1 0 33304 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_385
timestamp 1667941163
transform 1 0 36524 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_9
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_134
timestamp 1667941163
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_140
timestamp 1667941163
transform 1 0 13984 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_152
timestamp 1667941163
transform 1 0 15088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1667941163
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_211
timestamp 1667941163
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_376
timestamp 1667941163
transform 1 0 35696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_384
timestamp 1667941163
transform 1 0 36432 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_385
timestamp 1667941163
transform 1 0 36524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_7
timestamp 1667941163
transform 1 0 1748 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_19
timestamp 1667941163
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_31
timestamp 1667941163
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_43
timestamp 1667941163
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_381
timestamp 1667941163
transform 1 0 36156 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_384
timestamp 1667941163
transform 1 0 36432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1667941163
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_257
timestamp 1667941163
transform 1 0 24748 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_269
timestamp 1667941163
transform 1 0 25852 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_281
timestamp 1667941163
transform 1 0 26956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_293
timestamp 1667941163
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1667941163
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_370
timestamp 1667941163
transform 1 0 35144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_376
timestamp 1667941163
transform 1 0 35696 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_384
timestamp 1667941163
transform 1 0 36432 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_311
timestamp 1667941163
transform 1 0 29716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_315
timestamp 1667941163
transform 1 0 30084 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_321
timestamp 1667941163
transform 1 0 30636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1667941163
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_385
timestamp 1667941163
transform 1 0 36524 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_7
timestamp 1667941163
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_19
timestamp 1667941163
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_31
timestamp 1667941163
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_43
timestamp 1667941163
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_309
timestamp 1667941163
transform 1 0 29532 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_315
timestamp 1667941163
transform 1 0 30084 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_327
timestamp 1667941163
transform 1 0 31188 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1667941163
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_373
timestamp 1667941163
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_376
timestamp 1667941163
transform 1 0 35696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_384
timestamp 1667941163
transform 1 0 36432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1667941163
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_19
timestamp 1667941163
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1667941163
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_43
timestamp 1667941163
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1667941163
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_236
timestamp 1667941163
transform 1 0 22816 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_248
timestamp 1667941163
transform 1 0 23920 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_260
timestamp 1667941163
transform 1 0 25024 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1667941163
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_381
timestamp 1667941163
transform 1 0 36156 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_384
timestamp 1667941163
transform 1 0 36432 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1667941163
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_373
timestamp 1667941163
transform 1 0 35420 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_384
timestamp 1667941163
transform 1 0 36432 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_385
timestamp 1667941163
transform 1 0 36524 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_381
timestamp 1667941163
transform 1 0 36156 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_384
timestamp 1667941163
transform 1 0 36432 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1667941163
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1667941163
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_213
timestamp 1667941163
transform 1 0 20700 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_217
timestamp 1667941163
transform 1 0 21068 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_223
timestamp 1667941163
transform 1 0 21620 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_235
timestamp 1667941163
transform 1 0 22724 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_247
timestamp 1667941163
transform 1 0 23828 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_373
timestamp 1667941163
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_384
timestamp 1667941163
transform 1 0 36432 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1667941163
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_13
timestamp 1667941163
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_25
timestamp 1667941163
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_37
timestamp 1667941163
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_49
timestamp 1667941163
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_286
timestamp 1667941163
transform 1 0 27416 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_292
timestamp 1667941163
transform 1 0 27968 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_304
timestamp 1667941163
transform 1 0 29072 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_316
timestamp 1667941163
transform 1 0 30176 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1667941163
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_377
timestamp 1667941163
transform 1 0 35788 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_381
timestamp 1667941163
transform 1 0 36156 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_370
timestamp 1667941163
transform 1 0 35144 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_384
timestamp 1667941163
transform 1 0 36432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_17
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_25
timestamp 1667941163
transform 1 0 3404 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_28
timestamp 1667941163
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_40
timestamp 1667941163
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1667941163
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_74
timestamp 1667941163
transform 1 0 7912 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_80
timestamp 1667941163
transform 1 0 8464 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_92
timestamp 1667941163
transform 1 0 9568 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_104
timestamp 1667941163
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_122
timestamp 1667941163
transform 1 0 12328 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_128
timestamp 1667941163
transform 1 0 12880 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_140
timestamp 1667941163
transform 1 0 13984 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_152
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1667941163
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_191
timestamp 1667941163
transform 1 0 18676 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_199
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_211
timestamp 1667941163
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_310
timestamp 1667941163
transform 1 0 29624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_314
timestamp 1667941163
transform 1 0 29992 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_320
timestamp 1667941163
transform 1 0 30544 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1667941163
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1667941163
transform 1 0 34684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_368
timestamp 1667941163
transform 1 0 34960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_376
timestamp 1667941163
transform 1 0 35696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_384
timestamp 1667941163
transform 1 0 36432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_21
timestamp 1667941163
transform 1 0 3036 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_50
timestamp 1667941163
transform 1 0 5704 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_160
timestamp 1667941163
transform 1 0 15824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1667941163
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_239
timestamp 1667941163
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1667941163
transform 1 0 26036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_275
timestamp 1667941163
transform 1 0 26404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_323
timestamp 1667941163
transform 1 0 30820 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_329
timestamp 1667941163
transform 1 0 31372 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_345
timestamp 1667941163
transform 1 0 32844 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 36892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 36892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 36892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 36892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 36892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 36892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 36892 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 36892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 36892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 36892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 36892 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 36892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 36892 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 36892 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 36892 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 36892 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 36892 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 36892 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 36892 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 36892 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 36892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 36892 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _236_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 29992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29808 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 25944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 26772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 29992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform -1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 30452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform -1 0 27600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform -1 0 29348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform -1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _248_
timestamp 1667941163
transform 1 0 32476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform -1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 26680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform -1 0 30084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform -1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 27968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 27968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 28704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform -1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform 1 0 35052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform -1 0 12144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 11224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 10580 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform -1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform -1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform 1 0 11684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform 1 0 20056 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 30728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 31280 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform 1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform 1 0 13800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform -1 0 29348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform -1 0 31188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform 1 0 29716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform 1 0 11224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform -1 0 17940 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 27048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform -1 0 19228 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform -1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 29256 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform -1 0 28704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform 1 0 27140 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 29072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform -1 0 29992 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 27784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform 1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 21160 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform -1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform 1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform -1 0 23000 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform -1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform 1 0 26496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform -1 0 27416 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform 1 0 30176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform -1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform 1 0 16928 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform 1 0 21252 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform 1 0 17112 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform -1 0 21436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform -1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform -1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform 1 0 12328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform -1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform -1 0 11224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform 1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform -1 0 13156 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform 1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 10120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform 1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform -1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform -1 0 9936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform -1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform 1 0 14444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform 1 0 22632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform 1 0 26312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform -1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform -1 0 29808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform -1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 20516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform 1 0 12880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform -1 0 19412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform -1 0 26680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform -1 0 26496 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform -1 0 26220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform 1 0 29624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform 1 0 19504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform 1 0 11960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform -1 0 22264 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform -1 0 13800 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform -1 0 19872 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform 1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform -1 0 12420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 21160 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform -1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform -1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform 1 0 27784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform -1 0 20424 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform 1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform 1 0 16652 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform -1 0 12696 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform 1 0 28520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1667941163
transform 1 0 22356 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1667941163
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform -1 0 26404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform -1 0 19044 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1667941163
transform 1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1667941163
transform -1 0 26772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform 1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform -1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1667941163
transform 1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform -1 0 23736 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform 1 0 13156 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform 1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform -1 0 29992 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform 1 0 29716 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1667941163
transform -1 0 25024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 20240 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform -1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1667941163
transform -1 0 30084 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform -1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform 1 0 11224 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform 1 0 23736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 17664 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform -1 0 25208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform -1 0 12144 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform 1 0 20240 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform -1 0 27416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1667941163
transform -1 0 29992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _428_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 7912 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform -1 0 23552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 31188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform -1 0 28060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1667941163
transform 1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform 1 0 10396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform 1 0 9936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform -1 0 31096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1667941163
transform -1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform 1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform -1 0 28796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform -1 0 11316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 1667941163
transform 1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform -1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform -1 0 7728 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1667941163
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _455_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 30820 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _456_
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform -1 0 29348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform -1 0 23920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform -1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform -1 0 26128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform 1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform -1 0 27600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1667941163
transform -1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1667941163
transform -1 0 28704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1667941163
transform -1 0 23276 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _467_
timestamp 1667941163
transform -1 0 29256 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1667941163
transform -1 0 18952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1667941163
transform -1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1667941163
transform -1 0 18952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1667941163
transform -1 0 17296 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1667941163
transform -1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1667941163
transform -1 0 20332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1667941163
transform 1 0 19872 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1667941163
transform -1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1667941163
transform -1 0 22264 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1667941163
transform -1 0 24932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _478_
timestamp 1667941163
transform -1 0 29900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1667941163
transform -1 0 24104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1667941163
transform -1 0 27416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1667941163
transform -1 0 25576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1667941163
transform -1 0 25484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1667941163
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 1667941163
transform -1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _485_
timestamp 1667941163
transform -1 0 24840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1667941163
transform -1 0 25392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1667941163
transform -1 0 27416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1667941163
transform -1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _489_
timestamp 1667941163
transform -1 0 29808 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 1667941163
transform -1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1667941163
transform -1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1667941163
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _493_
timestamp 1667941163
transform 1 0 13064 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1667941163
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _495_
timestamp 1667941163
transform -1 0 23644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1667941163
transform 1 0 18032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _497_
timestamp 1667941163
transform 1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1667941163
transform 1 0 14444 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _499_
timestamp 1667941163
transform 1 0 14720 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _500_
timestamp 1667941163
transform 1 0 29716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _501_
timestamp 1667941163
transform -1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1667941163
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1667941163
transform -1 0 29808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 1667941163
transform -1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1667941163
transform -1 0 28060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1667941163
transform -1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1667941163
transform -1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 1667941163
transform -1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1667941163
transform 1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _510_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27048 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _511_
timestamp 1667941163
transform 1 0 24564 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform 1 0 21896 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _513_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _514_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _515_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20700 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _517_
timestamp 1667941163
transform -1 0 26404 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _519_
timestamp 1667941163
transform 1 0 14904 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _520_
timestamp 1667941163
transform -1 0 17020 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1667941163
transform -1 0 22908 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp 1667941163
transform 1 0 11960 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _523_
timestamp 1667941163
transform -1 0 14076 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform -1 0 16376 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _525_
timestamp 1667941163
transform -1 0 16376 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _526_
timestamp 1667941163
transform -1 0 23092 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _527_
timestamp 1667941163
transform -1 0 26680 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp 1667941163
transform -1 0 11592 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp 1667941163
transform 1 0 11960 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _531_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _532_
timestamp 1667941163
transform 1 0 23368 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _533_
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 1667941163
transform 1 0 19688 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _535_
timestamp 1667941163
transform 1 0 22172 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _537_
timestamp 1667941163
transform -1 0 16376 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _538_
timestamp 1667941163
transform 1 0 15640 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _539_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _540_
timestamp 1667941163
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _541_
timestamp 1667941163
transform -1 0 13800 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _542_
timestamp 1667941163
transform -1 0 26404 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _543_
timestamp 1667941163
transform -1 0 20148 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _544_
timestamp 1667941163
transform -1 0 21528 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _545_
timestamp 1667941163
transform -1 0 17664 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _546_
timestamp 1667941163
transform -1 0 21804 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _547_
timestamp 1667941163
transform -1 0 23828 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _548_
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _549_
timestamp 1667941163
transform 1 0 17388 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _550_
timestamp 1667941163
transform 1 0 16008 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _551_
timestamp 1667941163
transform 1 0 16008 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _552_
timestamp 1667941163
transform -1 0 28980 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _553_
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _554_
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _555_
timestamp 1667941163
transform 1 0 15088 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _556_
timestamp 1667941163
transform -1 0 16376 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _557_
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _558_
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _559_
timestamp 1667941163
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _560_
timestamp 1667941163
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _561_
timestamp 1667941163
transform 1 0 15088 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _562_
timestamp 1667941163
transform 1 0 23644 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _563_
timestamp 1667941163
transform 1 0 18952 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _564_
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _565_
timestamp 1667941163
transform -1 0 23828 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _566_
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _567_
timestamp 1667941163
transform -1 0 24564 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _568_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _569_
timestamp 1667941163
transform 1 0 20516 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _570_
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _571_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _572_
timestamp 1667941163
transform 1 0 22264 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _573_
timestamp 1667941163
transform 1 0 19044 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _574_
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _575_
timestamp 1667941163
transform 1 0 24472 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _576_
timestamp 1667941163
transform 1 0 11960 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _577_
timestamp 1667941163
transform 1 0 12328 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _578_
timestamp 1667941163
transform -1 0 16376 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _579_
timestamp 1667941163
transform 1 0 14444 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _580_
timestamp 1667941163
transform 1 0 14444 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _581_
timestamp 1667941163
transform -1 0 24104 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _594_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 29532 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _595_
timestamp 1667941163
transform -1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 1667941163
transform -1 0 36156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _597_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _598_
timestamp 1667941163
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _599_
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _600_
timestamp 1667941163
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _601_
timestamp 1667941163
transform -1 0 29348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _602_
timestamp 1667941163
transform -1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _603_
timestamp 1667941163
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _604_
timestamp 1667941163
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _605_
timestamp 1667941163
transform -1 0 31372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _606_
timestamp 1667941163
transform -1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _607_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _608_
timestamp 1667941163
transform 1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _609_
timestamp 1667941163
transform 1 0 31188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _610_
timestamp 1667941163
transform -1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _611_
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _612_
timestamp 1667941163
transform -1 0 22264 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _613_
timestamp 1667941163
transform -1 0 36156 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _614_
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _615_
timestamp 1667941163
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _616_
timestamp 1667941163
transform -1 0 26128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _617_
timestamp 1667941163
transform -1 0 27416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _618_
timestamp 1667941163
transform -1 0 21068 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _619_
timestamp 1667941163
transform 1 0 12052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _620_
timestamp 1667941163
transform 1 0 30360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _621_
timestamp 1667941163
transform -1 0 18400 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _622_
timestamp 1667941163
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _623_
timestamp 1667941163
transform -1 0 21528 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _624_
timestamp 1667941163
transform -1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _625_
timestamp 1667941163
transform -1 0 32568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _626_
timestamp 1667941163
transform 1 0 1748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _627_
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _628_
timestamp 1667941163
transform -1 0 36248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _629_
timestamp 1667941163
transform -1 0 14536 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _630_
timestamp 1667941163
transform -1 0 27416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _631_
timestamp 1667941163
transform -1 0 9568 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _632_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform 1 0 19872 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform 1 0 14904 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _635_
timestamp 1667941163
transform 1 0 13984 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform 1 0 26956 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _636__92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform 1 0 25760 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _638_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27876 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _639_
timestamp 1667941163
transform 1 0 23184 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform -1 0 18308 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 25392 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _643_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _644_
timestamp 1667941163
transform -1 0 25760 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform 1 0 17848 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform -1 0 20424 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _647_
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _648__93
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform -1 0 23000 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _649_
timestamp 1667941163
transform 1 0 22264 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform -1 0 23000 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _651_
timestamp 1667941163
transform 1 0 18584 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _652_
timestamp 1667941163
transform 1 0 22448 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _653_
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _654_
timestamp 1667941163
transform 1 0 17572 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _655_
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _656_
timestamp 1667941163
transform -1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform -1 0 16928 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform -1 0 19504 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _659__94
timestamp 1667941163
transform 1 0 15364 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _659_
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _660_
timestamp 1667941163
transform 1 0 24380 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _661_
timestamp 1667941163
transform 1 0 14904 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _662_
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform -1 0 15732 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _665_
timestamp 1667941163
transform -1 0 21620 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform -1 0 25392 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _667_
timestamp 1667941163
transform -1 0 20240 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _668_
timestamp 1667941163
transform 1 0 17204 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _669_
timestamp 1667941163
transform -1 0 20700 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform -1 0 27784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform -1 0 23920 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _671__95
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform -1 0 22816 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _673_
timestamp 1667941163
transform 1 0 15640 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform -1 0 26588 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _675_
timestamp 1667941163
transform -1 0 25760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _676_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform -1 0 26128 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform -1 0 20792 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _679_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _680_
timestamp 1667941163
transform 1 0 17296 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _681_
timestamp 1667941163
transform -1 0 27416 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform -1 0 28888 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _683_
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _683__96
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform 1 0 14444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _685_
timestamp 1667941163
transform 1 0 12604 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform 1 0 20976 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _688_
timestamp 1667941163
transform 1 0 23368 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform 1 0 14536 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 12788 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform -1 0 26220 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform -1 0 10948 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform 1 0 9200 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform -1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _695_
timestamp 1667941163
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _695__97
timestamp 1667941163
transform 1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform -1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform 1 0 10672 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform 1 0 11592 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform -1 0 11224 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform 1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform -1 0 11224 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _704_
timestamp 1667941163
transform 1 0 14168 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _705_
timestamp 1667941163
transform -1 0 18952 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform -1 0 25392 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _707__98
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _708_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13524 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _709_
timestamp 1667941163
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _710_
timestamp 1667941163
transform 1 0 12420 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _711_
timestamp 1667941163
transform -1 0 17480 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _712_
timestamp 1667941163
transform -1 0 13800 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _713_
timestamp 1667941163
transform -1 0 25208 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _714_
timestamp 1667941163
transform -1 0 14444 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _715_
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _716_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _717_
timestamp 1667941163
transform 1 0 27784 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _718_
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _719_
timestamp 1667941163
transform 1 0 22172 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _719__99
timestamp 1667941163
transform -1 0 22264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _720_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _721_
timestamp 1667941163
transform 1 0 21068 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _722_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _723_
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _724_
timestamp 1667941163
transform 1 0 27324 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _725_
timestamp 1667941163
transform 1 0 25576 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _726_
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _727_
timestamp 1667941163
transform -1 0 21160 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _728_
timestamp 1667941163
transform 1 0 25300 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _729_
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _730_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _731__100
timestamp 1667941163
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _731_
timestamp 1667941163
transform 1 0 23184 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _732_
timestamp 1667941163
transform -1 0 24472 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _733_
timestamp 1667941163
transform 1 0 16836 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _734_
timestamp 1667941163
transform 1 0 17296 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _735_
timestamp 1667941163
transform 1 0 16100 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _736_
timestamp 1667941163
transform 1 0 22816 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _737_
timestamp 1667941163
transform 1 0 22264 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _738_
timestamp 1667941163
transform 1 0 22264 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _739_
timestamp 1667941163
transform -1 0 23552 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _740_
timestamp 1667941163
transform 1 0 28336 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _741_
timestamp 1667941163
transform 1 0 28336 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _742_
timestamp 1667941163
transform -1 0 29348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _743__101
timestamp 1667941163
transform -1 0 28704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _743_
timestamp 1667941163
transform -1 0 28612 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _744_
timestamp 1667941163
transform -1 0 26956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _745_
timestamp 1667941163
transform 1 0 15364 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _746_
timestamp 1667941163
transform -1 0 28428 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _747_
timestamp 1667941163
transform -1 0 27232 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _748_
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _749_
timestamp 1667941163
transform 1 0 28244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _750_
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _751_
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _752_
timestamp 1667941163
transform 1 0 27324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _753_
timestamp 1667941163
transform 1 0 31372 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _754_
timestamp 1667941163
transform -1 0 30544 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _755__102
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _755_
timestamp 1667941163
transform -1 0 25392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _756_
timestamp 1667941163
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _757_
timestamp 1667941163
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _758_
timestamp 1667941163
transform 1 0 22172 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _759_
timestamp 1667941163
transform 1 0 29716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _760_
timestamp 1667941163
transform -1 0 30820 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _761_
timestamp 1667941163
transform 1 0 17204 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _762_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _763_
timestamp 1667941163
transform -1 0 30544 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _764_
timestamp 1667941163
transform -1 0 15180 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _765_
timestamp 1667941163
transform -1 0 23184 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _766_
timestamp 1667941163
transform -1 0 20884 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _767_
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _767__103
timestamp 1667941163
transform -1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _768_
timestamp 1667941163
transform -1 0 20792 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _769_
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _770_
timestamp 1667941163
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _771_
timestamp 1667941163
transform -1 0 13708 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _772_
timestamp 1667941163
transform -1 0 12512 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _773_
timestamp 1667941163
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _774_
timestamp 1667941163
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _775_
timestamp 1667941163
transform 1 0 11776 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21436 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1667941163
transform -1 0 18952 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1667941163
transform -1 0 13800 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1667941163
transform 1 0 11960 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1667941163
transform -1 0 23828 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1667941163
transform -1 0 28980 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1667941163
transform 1 0 17388 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1667941163
transform -1 0 26404 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform -1 0 36432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform -1 0 2484 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform -1 0 36432 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1667941163
transform -1 0 36432 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 35512 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1667941163
transform -1 0 36432 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform -1 0 36432 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1667941163
transform -1 0 30636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform -1 0 36432 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1667941163
transform 1 0 32936 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 36156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform -1 0 36432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1667941163
transform -1 0 27140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform -1 0 36432 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 29716 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 36156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 36064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 14904 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 36064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform 1 0 22724 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform 1 0 36064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform 1 0 36064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform -1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 36064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 36064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform -1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform -1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform -1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 36064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 32936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 1932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 35328 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 36064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 10856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform -1 0 18952 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform -1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform -1 0 3496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 27508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform -1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform -1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 36064 0 -1 19584
box -38 -48 406 592
<< labels >>
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 0 nsew signal tristate
flabel metal3 s 37200 25848 37800 25968 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 1 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 2 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
port 3 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 37200 10208 37800 10328 0 FreeSans 480 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 37200 27888 37800 28008 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 37200 31288 37800 31408 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 37200 34688 37800 34808 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 37200 36048 37800 36168 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 37200 32648 37800 32768 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal3 s 37200 4768 37800 4888 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal3 s 37200 29248 37800 29368 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal3 s 37200 8 37800 128 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal3 s 37200 17008 37800 17128 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal3 s 37200 20408 37800 20528 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal3 s 37200 8168 37800 8288 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal3 s 37200 15648 37800 15768 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal3 s 37200 13608 37800 13728 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal3 s 37200 6808 37800 6928 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal3 s 37200 1368 37800 1488 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal3 s 37200 11568 37800 11688 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal3 s 37200 38088 37800 38208 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal3 s 37200 3408 37800 3528 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal3 s 37200 22448 37800 22568 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal3 s 37200 23808 37800 23928 0 FreeSans 480 0 0 0 pReset
port 82 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 prog_clk
port 83 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 84 nsew signal tristate
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_
port 85 nsew signal tristate
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_
port 86 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_
port 87 nsew signal tristate
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_
port 88 nsew signal tristate
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_
port 89 nsew signal tristate
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_
port 90 nsew signal tristate
flabel metal3 s 37200 19048 37800 19168 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_
port 91 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 92 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 92 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 93 nsew ground bidirectional
rlabel metal1 18998 37536 18998 37536 0 vccd1
rlabel metal1 18998 36992 18998 36992 0 vssd1
rlabel metal2 29210 8194 29210 8194 0 _000_
rlabel metal1 27738 7174 27738 7174 0 _001_
rlabel metal1 23605 7786 23605 7786 0 _002_
rlabel metal1 21298 11016 21298 11016 0 _003_
rlabel metal1 24656 11254 24656 11254 0 _004_
rlabel metal1 20286 7480 20286 7480 0 _005_
rlabel metal1 25990 4631 25990 4631 0 _006_
rlabel metal2 25530 6494 25530 6494 0 _007_
rlabel metal1 26503 11798 26503 11798 0 _008_
rlabel metal1 17855 6766 17855 6766 0 _009_
rlabel metal1 18814 10200 18814 10200 0 _010_
rlabel metal1 28244 7990 28244 7990 0 _011_
rlabel metal1 14129 6766 14129 6766 0 _012_
rlabel metal1 13485 5270 13485 5270 0 _013_
rlabel metal1 16705 6358 16705 6358 0 _014_
rlabel metal1 18768 9078 18768 9078 0 _015_
rlabel metal1 20562 9894 20562 9894 0 _016_
rlabel metal1 28014 8602 28014 8602 0 _017_
rlabel metal1 13577 2346 13577 2346 0 _018_
rlabel metal2 18998 12517 18998 12517 0 _019_
rlabel metal1 21114 7208 21114 7208 0 _020_
rlabel metal1 26135 8942 26135 8942 0 _021_
rlabel metal2 25438 10166 25438 10166 0 _022_
rlabel metal2 23230 9044 23230 9044 0 _023_
rlabel metal1 21114 4699 21114 4699 0 _024_
rlabel metal1 24065 3434 24065 3434 0 _025_
rlabel metal1 13577 5610 13577 5610 0 _026_
rlabel metal2 15042 3145 15042 3145 0 _027_
rlabel metal2 17066 6052 17066 6052 0 _028_
rlabel metal1 21029 2346 21029 2346 0 _029_
rlabel metal1 13807 3502 13807 3502 0 _030_
rlabel metal1 20884 9350 20884 9350 0 _031_
rlabel metal1 23085 2414 23085 2414 0 _032_
rlabel metal1 14766 10778 14766 10778 0 _033_
rlabel metal1 18945 7786 18945 7786 0 _034_
rlabel metal2 16330 5695 16330 5695 0 _035_
rlabel metal1 18584 9894 18584 9894 0 _036_
rlabel metal2 17986 6868 17986 6868 0 _037_
rlabel metal2 20746 10506 20746 10506 0 _038_
rlabel metal1 15502 9078 15502 9078 0 _039_
rlabel metal1 18453 8942 18453 8942 0 _040_
rlabel metal1 17763 3434 17763 3434 0 _041_
rlabel metal1 28941 4182 28941 4182 0 _042_
rlabel metal1 28895 2346 28895 2346 0 _043_
rlabel metal1 27876 9350 27876 9350 0 _044_
rlabel metal1 17257 10030 17257 10030 0 _045_
rlabel metal2 20654 9894 20654 9894 0 _046_
rlabel metal1 25162 9350 25162 9350 0 _047_
rlabel via2 18538 4165 18538 4165 0 _048_
rlabel metal2 22034 9265 22034 9265 0 _049_
rlabel via2 19274 10693 19274 10693 0 _050_
rlabel metal1 17165 7786 17165 7786 0 _051_
rlabel metal1 26128 11322 26128 11322 0 _052_
rlabel metal2 24794 6222 24794 6222 0 _053_
rlabel metal1 27278 2550 27278 2550 0 _054_
rlabel metal1 23283 4182 23283 4182 0 _055_
rlabel metal1 26680 7922 26680 7922 0 _056_
rlabel metal1 28014 9146 28014 9146 0 _057_
rlabel metal1 26641 7786 26641 7786 0 _058_
rlabel metal2 21942 8466 21942 8466 0 _059_
rlabel metal1 32407 3094 32407 3094 0 _060_
rlabel metal1 31142 3468 31142 3468 0 _061_
rlabel metal1 24065 4590 24065 4590 0 _062_
rlabel metal2 21850 5576 21850 5576 0 _063_
rlabel metal1 21144 3026 21144 3026 0 _064_
rlabel metal1 29762 3910 29762 3910 0 _065_
rlabel metal1 14129 4182 14129 4182 0 _066_
rlabel via2 13754 6307 13754 6307 0 _067_
rlabel metal2 15594 4641 15594 4641 0 _068_
rlabel via2 16514 5253 16514 5253 0 _069_
rlabel metal2 32062 6698 32062 6698 0 _070_
rlabel metal2 31602 3162 31602 3162 0 _071_
rlabel metal1 32154 3536 32154 3536 0 _072_
rlabel metal1 28842 7854 28842 7854 0 _073_
rlabel metal1 18906 11084 18906 11084 0 _074_
rlabel metal2 28842 7582 28842 7582 0 _075_
rlabel metal1 20930 9554 20930 9554 0 _076_
rlabel metal2 22770 11169 22770 11169 0 _077_
rlabel metal1 29164 9554 29164 9554 0 _078_
rlabel metal2 31786 3842 31786 3842 0 _079_
rlabel metal2 23598 15912 23598 15912 0 _080_
rlabel metal2 19642 20264 19642 20264 0 _081_
rlabel metal1 14996 17238 14996 17238 0 _082_
rlabel metal1 14766 18326 14766 18326 0 _083_
rlabel metal2 27186 20026 27186 20026 0 _084_
rlabel metal2 25990 19992 25990 19992 0 _085_
rlabel metal1 29808 12954 29808 12954 0 _086_
rlabel metal1 25760 14042 25760 14042 0 _087_
rlabel metal2 21482 18088 21482 18088 0 _088_
rlabel metal2 18078 17646 18078 17646 0 _089_
rlabel metal2 25622 18462 25622 18462 0 _090_
rlabel metal1 29164 13362 29164 13362 0 _091_
rlabel metal1 25530 14280 25530 14280 0 _092_
rlabel metal1 18124 15402 18124 15402 0 _093_
rlabel metal1 20148 15062 20148 15062 0 _094_
rlabel metal1 13938 16150 13938 16150 0 _095_
rlabel metal2 22770 17544 22770 17544 0 _096_
rlabel metal2 25346 13872 25346 13872 0 _097_
rlabel metal2 22770 20638 22770 20638 0 _098_
rlabel metal2 16974 18904 16974 18904 0 _099_
rlabel metal1 27140 12750 27140 12750 0 _100_
rlabel metal2 24978 17918 24978 17918 0 _101_
rlabel metal1 17296 18326 17296 18326 0 _102_
rlabel metal2 20286 18462 20286 18462 0 _103_
rlabel metal1 14720 16490 14720 16490 0 _104_
rlabel metal1 16836 16422 16836 16422 0 _105_
rlabel metal2 19274 17374 19274 17374 0 _106_
rlabel metal1 15180 20570 15180 20570 0 _107_
rlabel metal2 22494 15538 22494 15538 0 _108_
rlabel metal2 15134 15674 15134 15674 0 _109_
rlabel metal1 16744 18938 16744 18938 0 _110_
rlabel metal2 15502 18088 15502 18088 0 _111_
rlabel metal1 15548 18326 15548 18326 0 _112_
rlabel metal2 21022 22882 21022 22882 0 _113_
rlabel metal1 24656 12614 24656 12614 0 _114_
rlabel metal1 19872 22406 19872 22406 0 _115_
rlabel metal2 12098 13226 12098 13226 0 _116_
rlabel metal2 19826 12512 19826 12512 0 _117_
rlabel metal2 27554 15674 27554 15674 0 _118_
rlabel metal1 25484 17306 25484 17306 0 _119_
rlabel metal1 22356 14042 22356 14042 0 _120_
rlabel via1 13662 14773 13662 14773 0 _121_
rlabel metal1 24380 13498 24380 13498 0 _122_
rlabel metal1 25990 13974 25990 13974 0 _123_
rlabel metal2 19366 11968 19366 11968 0 _124_
rlabel metal2 25898 18904 25898 18904 0 _125_
rlabel metal1 20378 14314 20378 14314 0 _126_
rlabel metal1 19136 12954 19136 12954 0 _127_
rlabel metal1 19090 9486 19090 9486 0 _128_
rlabel metal1 27186 13192 27186 13192 0 _129_
rlabel metal1 29486 10710 29486 10710 0 _130_
rlabel metal1 15502 11560 15502 11560 0 _131_
rlabel metal1 13846 9962 13846 9962 0 _132_
rlabel metal1 12834 8840 12834 8840 0 _133_
rlabel metal1 21022 13192 21022 13192 0 _134_
rlabel metal1 15778 12920 15778 12920 0 _135_
rlabel metal2 23598 14093 23598 14093 0 _136_
rlabel metal1 14030 9622 14030 9622 0 _137_
rlabel metal2 13018 10642 13018 10642 0 _138_
rlabel metal1 26036 12886 26036 12886 0 _139_
rlabel metal1 10856 8058 10856 8058 0 _140_
rlabel metal1 9338 5882 9338 5882 0 _141_
rlabel metal1 19320 11322 19320 11322 0 _142_
rlabel metal2 8050 11560 8050 11560 0 _143_
rlabel metal1 15594 11322 15594 11322 0 _144_
rlabel metal1 12627 12886 12627 12886 0 _145_
rlabel metal2 10902 11322 10902 11322 0 _146_
rlabel metal1 11822 13192 11822 13192 0 _147_
rlabel metal1 10764 6970 10764 6970 0 _148_
rlabel metal2 9798 5032 9798 5032 0 _149_
rlabel metal1 10994 13192 10994 13192 0 _150_
rlabel metal1 10902 13838 10902 13838 0 _151_
rlabel metal2 14398 14824 14398 14824 0 _152_
rlabel metal1 19826 9146 19826 9146 0 _153_
rlabel metal1 25162 19720 25162 19720 0 _154_
rlabel metal1 20194 19482 20194 19482 0 _155_
rlabel metal2 13294 17612 13294 17612 0 _156_
rlabel metal1 13156 16626 13156 16626 0 _157_
rlabel metal2 12650 14654 12650 14654 0 _158_
rlabel via2 17250 15419 17250 15419 0 _159_
rlabel metal1 13708 15062 13708 15062 0 _160_
rlabel metal1 24978 19448 24978 19448 0 _161_
rlabel metal2 13386 16558 13386 16558 0 _162_
rlabel metal1 13202 14280 13202 14280 0 _163_
rlabel metal1 27370 14008 27370 14008 0 _164_
rlabel metal1 27646 10778 27646 10778 0 _165_
rlabel metal1 17112 15062 17112 15062 0 _166_
rlabel metal2 21390 13056 21390 13056 0 _167_
rlabel metal1 17112 16150 17112 16150 0 _168_
rlabel metal2 21298 14994 21298 14994 0 _169_
rlabel metal1 19642 17544 19642 17544 0 _170_
rlabel metal1 22678 14008 22678 14008 0 _171_
rlabel metal1 30222 13974 30222 13974 0 _172_
rlabel metal1 24886 14586 24886 14586 0 _173_
rlabel metal1 17664 15130 17664 15130 0 _174_
rlabel metal1 21068 16762 21068 16762 0 _175_
rlabel metal1 26082 16150 26082 16150 0 _176_
rlabel metal1 25484 11866 25484 11866 0 _177_
rlabel metal2 23506 16796 23506 16796 0 _178_
rlabel metal2 21482 19550 21482 19550 0 _179_
rlabel metal1 24242 16184 24242 16184 0 _180_
rlabel metal1 17066 13192 17066 13192 0 _181_
rlabel metal1 17296 17578 17296 17578 0 _182_
rlabel metal1 16284 17306 16284 17306 0 _183_
rlabel metal1 21620 12342 21620 12342 0 _184_
rlabel metal2 22862 21794 22862 21794 0 _185_
rlabel metal1 22448 15402 22448 15402 0 _186_
rlabel metal1 23322 19720 23322 19720 0 _187_
rlabel metal1 28244 13974 28244 13974 0 _188_
rlabel metal2 28566 13260 28566 13260 0 _189_
rlabel metal1 29486 14994 29486 14994 0 _190_
rlabel metal2 28382 16252 28382 16252 0 _191_
rlabel metal2 30498 14892 30498 14892 0 _192_
rlabel metal1 15594 14280 15594 14280 0 _193_
rlabel metal1 28658 16218 28658 16218 0 _194_
rlabel metal2 27002 16728 27002 16728 0 _195_
rlabel metal1 27416 10234 27416 10234 0 _196_
rlabel metal1 28106 17714 28106 17714 0 _197_
rlabel metal1 16790 14280 16790 14280 0 _198_
rlabel metal2 18354 14552 18354 14552 0 _199_
rlabel metal1 29164 11866 29164 11866 0 _200_
rlabel metal2 31786 7378 31786 7378 0 _201_
rlabel metal1 30314 9928 30314 9928 0 _202_
rlabel metal1 27416 11526 27416 11526 0 _203_
rlabel metal1 16146 13838 16146 13838 0 _204_
rlabel metal2 12466 11934 12466 11934 0 _205_
rlabel metal1 23644 12886 23644 12886 0 _206_
rlabel metal2 29854 11730 29854 11730 0 _207_
rlabel metal1 30728 4794 30728 4794 0 _208_
rlabel metal1 14628 9486 14628 9486 0 _209_
rlabel metal1 14490 13192 14490 13192 0 _210_
rlabel metal1 30728 12954 30728 12954 0 _211_
rlabel metal1 15226 12886 15226 12886 0 _212_
rlabel metal2 27278 11951 27278 11951 0 _213_
rlabel metal1 20102 12886 20102 12886 0 _214_
rlabel metal1 16008 11866 16008 11866 0 _215_
rlabel metal1 20378 12410 20378 12410 0 _216_
rlabel metal1 13052 13226 13052 13226 0 _217_
rlabel metal1 11270 12614 11270 12614 0 _218_
rlabel metal2 13478 13158 13478 13158 0 _219_
rlabel metal2 12006 9112 12006 9112 0 _220_
rlabel metal2 11454 6120 11454 6120 0 _221_
rlabel metal2 11454 9384 11454 9384 0 _222_
rlabel metal1 11868 10234 11868 10234 0 _223_
rlabel metal1 34776 37094 34776 37094 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
rlabel metal3 36532 25908 36532 25908 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
rlabel metal2 36110 1520 36110 1520 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal1 14996 3366 14996 3366 0 bottom_grid_top_width_0_height_0_subtile_0__pin_clk_0_
rlabel metal1 26496 37434 26496 37434 0 ccff_head
rlabel metal2 36294 10353 36294 10353 0 ccff_tail
rlabel metal1 13018 37230 13018 37230 0 chanx_left_in[0]
rlabel metal1 16767 37230 16767 37230 0 chanx_left_in[10]
rlabel metal2 36294 27999 36294 27999 0 chanx_left_in[11]
rlabel metal2 2438 37723 2438 37723 0 chanx_left_in[12]
rlabel metal2 35834 31569 35834 31569 0 chanx_left_in[13]
rlabel metal1 19412 37298 19412 37298 0 chanx_left_in[14]
rlabel via2 36386 34731 36386 34731 0 chanx_left_in[15]
rlabel via2 1610 4811 1610 4811 0 chanx_left_in[16]
rlabel metal1 2576 2414 2576 2414 0 chanx_left_in[17]
rlabel via2 35558 36125 35558 36125 0 chanx_left_in[18]
rlabel metal2 36386 32623 36386 32623 0 chanx_left_in[1]
rlabel metal2 1702 32759 1702 32759 0 chanx_left_in[2]
rlabel via2 36386 4811 36386 4811 0 chanx_left_in[3]
rlabel metal1 1518 36822 1518 36822 0 chanx_left_in[4]
rlabel metal2 1610 20689 1610 20689 0 chanx_left_in[5]
rlabel metal1 31464 2482 31464 2482 0 chanx_left_in[6]
rlabel metal2 1610 19023 1610 19023 0 chanx_left_in[7]
rlabel via2 36386 29291 36386 29291 0 chanx_left_in[8]
rlabel metal2 36018 1547 36018 1547 0 chanx_left_in[9]
rlabel metal1 22770 37094 22770 37094 0 chanx_left_out[0]
rlabel metal1 2668 36890 2668 36890 0 chanx_left_out[10]
rlabel via2 36294 17051 36294 17051 0 chanx_left_out[11]
rlabel metal3 1188 15708 1188 15708 0 chanx_left_out[12]
rlabel metal2 7774 1520 7774 1520 0 chanx_left_out[13]
rlabel metal2 36294 20621 36294 20621 0 chanx_left_out[14]
rlabel metal1 14950 37094 14950 37094 0 chanx_left_out[15]
rlabel metal2 36294 8279 36294 8279 0 chanx_left_out[16]
rlabel metal1 24656 37094 24656 37094 0 chanx_left_out[17]
rlabel metal1 36846 36890 36846 36890 0 chanx_left_out[18]
rlabel metal2 34178 823 34178 823 0 chanx_left_out[1]
rlabel metal1 18170 37094 18170 37094 0 chanx_left_out[2]
rlabel metal2 30958 1520 30958 1520 0 chanx_left_out[3]
rlabel metal3 1188 3468 1188 3468 0 chanx_left_out[4]
rlabel metal2 10994 1520 10994 1520 0 chanx_left_out[5]
rlabel metal3 1188 27948 1188 27948 0 chanx_left_out[6]
rlabel metal2 36294 15793 36294 15793 0 chanx_left_out[7]
rlabel metal2 4554 1520 4554 1520 0 chanx_left_out[8]
rlabel metal3 1188 13668 1188 13668 0 chanx_left_out[9]
rlabel via2 1610 31365 1610 31365 0 chanx_right_in[0]
rlabel metal3 1142 6868 1142 6868 0 chanx_right_in[10]
rlabel via2 1610 29291 1610 29291 0 chanx_right_in[11]
rlabel metal1 6578 37230 6578 37230 0 chanx_right_in[12]
rlabel metal1 3312 2278 3312 2278 0 chanx_right_in[13]
rlabel metal2 9706 1761 9706 1761 0 chanx_right_in[14]
rlabel metal1 32936 2414 32936 2414 0 chanx_right_in[15]
rlabel metal2 36386 13787 36386 13787 0 chanx_right_in[16]
rlabel metal3 36532 6868 36532 6868 0 chanx_right_in[17]
rlabel metal2 24518 823 24518 823 0 chanx_right_in[18]
rlabel metal3 1188 36108 1188 36108 0 chanx_right_in[1]
rlabel metal2 36294 2227 36294 2227 0 chanx_right_in[2]
rlabel metal2 1610 8143 1610 8143 0 chanx_right_in[3]
rlabel metal2 36294 11679 36294 11679 0 chanx_right_in[4]
rlabel via2 1610 23851 1610 23851 0 chanx_right_in[5]
rlabel metal1 30084 3026 30084 3026 0 chanx_right_in[6]
rlabel metal2 1702 17119 1702 17119 0 chanx_right_in[7]
rlabel metal1 9798 37230 9798 37230 0 chanx_right_in[8]
rlabel metal1 4692 37230 4692 37230 0 chanx_right_in[9]
rlabel metal1 18170 2822 18170 2822 0 chanx_right_out[0]
rlabel metal2 46 1792 46 1792 0 chanx_right_out[10]
rlabel metal1 23092 3706 23092 3706 0 chanx_right_out[11]
rlabel metal1 11454 37094 11454 37094 0 chanx_right_out[12]
rlabel metal1 21758 37094 21758 37094 0 chanx_right_out[13]
rlabel metal2 33028 37094 33028 37094 0 chanx_right_out[14]
rlabel metal2 1702 26061 1702 26061 0 chanx_right_out[15]
rlabel metal3 1188 22508 1188 22508 0 chanx_right_out[16]
rlabel metal2 1334 1520 1334 1520 0 chanx_right_out[17]
rlabel metal1 36248 37094 36248 37094 0 chanx_right_out[18]
rlabel metal1 28198 37094 28198 37094 0 chanx_right_out[1]
rlabel metal2 16238 2788 16238 2788 0 chanx_right_out[2]
rlabel metal2 35558 37519 35558 37519 0 chanx_right_out[3]
rlabel metal2 36294 3417 36294 3417 0 chanx_right_out[4]
rlabel metal3 1188 10268 1188 10268 0 chanx_right_out[5]
rlabel via2 36294 22491 36294 22491 0 chanx_right_out[6]
rlabel metal2 6486 1520 6486 1520 0 chanx_right_out[7]
rlabel metal2 12926 1520 12926 1520 0 chanx_right_out[8]
rlabel metal1 19044 3366 19044 3366 0 chanx_right_out[9]
rlabel metal1 9016 3094 9016 3094 0 clknet_0_prog_clk
rlabel metal1 11776 2482 11776 2482 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15870 2482 15870 2482 0 clknet_3_1__leaf_prog_clk
rlabel metal1 14720 6834 14720 6834 0 clknet_3_2__leaf_prog_clk
rlabel metal1 14030 7378 14030 7378 0 clknet_3_3__leaf_prog_clk
rlabel metal1 22034 6324 22034 6324 0 clknet_3_4__leaf_prog_clk
rlabel metal2 24610 5712 24610 5712 0 clknet_3_5__leaf_prog_clk
rlabel metal1 21068 7922 21068 7922 0 clknet_3_6__leaf_prog_clk
rlabel metal1 23184 10642 23184 10642 0 clknet_3_7__leaf_prog_clk
rlabel metal1 18814 18258 18814 18258 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal1 15410 19822 15410 19822 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal1 14674 18700 14674 18700 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal1 24932 7718 24932 7718 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal1 26680 13906 26680 13906 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal1 29532 12818 29532 12818 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal3 19044 12580 19044 12580 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel via1 15219 6970 15219 6970 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal2 16974 6392 16974 6392 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel metal1 26404 12614 26404 12614 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal1 25300 5882 25300 5882 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal1 28474 14382 28474 14382 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal1 23000 22406 23000 22406 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal1 18952 17646 18952 17646 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal1 13202 16082 13202 16082 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal1 14490 6222 14490 6222 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal1 11904 6970 11904 6970 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal1 13662 6834 13662 6834 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal2 16146 13974 16146 13974 0 mem_bottom_ipin_3.DFFR_0_.Q
rlabel metal1 29670 16116 29670 16116 0 mem_bottom_ipin_3.DFFR_1_.Q
rlabel metal2 14950 7344 14950 7344 0 mem_bottom_ipin_3.DFFR_2_.Q
rlabel metal1 13708 7514 13708 7514 0 mem_bottom_ipin_3.DFFR_3_.Q
rlabel metal1 11960 2346 11960 2346 0 mem_bottom_ipin_3.DFFR_4_.Q
rlabel metal1 18952 12206 18952 12206 0 mem_bottom_ipin_3.DFFR_5_.Q
rlabel metal1 18952 1938 18952 1938 0 mem_bottom_ipin_4.DFFR_0_.Q
rlabel metal2 21942 10948 21942 10948 0 mem_bottom_ipin_4.DFFR_1_.Q
rlabel metal2 12742 2873 12742 2873 0 mem_bottom_ipin_4.DFFR_2_.Q
rlabel metal2 13570 3808 13570 3808 0 mem_bottom_ipin_4.DFFR_3_.Q
rlabel metal1 20056 4658 20056 4658 0 mem_bottom_ipin_4.DFFR_4_.Q
rlabel metal1 18124 4726 18124 4726 0 mem_bottom_ipin_4.DFFR_5_.Q
rlabel metal1 21068 7786 21068 7786 0 mem_bottom_ipin_5.DFFR_0_.Q
rlabel metal1 14076 11118 14076 11118 0 mem_bottom_ipin_5.DFFR_1_.Q
rlabel metal1 18078 8364 18078 8364 0 mem_bottom_ipin_5.DFFR_2_.Q
rlabel metal1 19550 2516 19550 2516 0 mem_bottom_ipin_5.DFFR_3_.Q
rlabel metal1 12098 3570 12098 3570 0 mem_bottom_ipin_5.DFFR_4_.Q
rlabel metal1 13754 3400 13754 3400 0 mem_bottom_ipin_5.DFFR_5_.Q
rlabel metal1 21252 19278 21252 19278 0 mem_bottom_ipin_6.DFFR_0_.Q
rlabel metal1 13570 18258 13570 18258 0 mem_bottom_ipin_6.DFFR_1_.Q
rlabel metal1 19964 19346 19964 19346 0 mem_bottom_ipin_6.DFFR_2_.Q
rlabel metal1 21574 11254 21574 11254 0 mem_bottom_ipin_6.DFFR_3_.Q
rlabel metal1 20332 4998 20332 4998 0 mem_bottom_ipin_6.DFFR_4_.Q
rlabel metal1 19826 8942 19826 8942 0 mem_bottom_ipin_6.DFFR_5_.Q
rlabel metal1 17204 14994 17204 14994 0 mem_bottom_ipin_7.DFFR_0_.Q
rlabel metal1 16284 14994 16284 14994 0 mem_bottom_ipin_7.DFFR_1_.Q
rlabel metal1 17388 10098 17388 10098 0 mem_bottom_ipin_7.DFFR_2_.Q
rlabel metal1 26772 2346 26772 2346 0 mem_bottom_ipin_7.DFFR_3_.Q
rlabel metal1 30498 14382 30498 14382 0 mem_bottom_ipin_7.DFFR_4_.Q
rlabel metal1 20654 5100 20654 5100 0 mem_bottom_ipin_7.DFFR_5_.Q
rlabel metal2 21298 18700 21298 18700 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal1 16100 19346 16100 19346 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal1 21160 19822 21160 19822 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal1 19274 10608 19274 10608 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal1 21436 10438 21436 10438 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 20884 6868 20884 6868 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal2 24886 8092 24886 8092 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal1 30176 15470 30176 15470 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal2 20838 14875 20838 14875 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal1 26726 5338 26726 5338 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal1 14674 2346 14674 2346 0 mem_top_ipin_1.DFFR_4_.Q
rlabel metal1 28520 4590 28520 4590 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal2 21482 2992 21482 2992 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal2 20148 12308 20148 12308 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal1 21068 4114 21068 4114 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal1 30774 4624 30774 4624 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal2 29762 7684 29762 7684 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal2 28566 3876 28566 3876 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal1 19182 6630 19182 6630 0 mem_top_ipin_3.DFFR_0_.Q
rlabel via2 12926 12869 12926 12869 0 mem_top_ipin_3.DFFR_1_.Q
rlabel metal1 16054 4216 16054 4216 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal1 13248 6222 13248 6222 0 mem_top_ipin_3.DFFR_3_.Q
rlabel metal1 14030 6154 14030 6154 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal2 20194 18020 20194 18020 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal1 20056 20366 20056 20366 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal2 17342 15538 17342 15538 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel via1 19366 15997 19366 15997 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 13708 27914 13708 27914 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal2 13110 16830 13110 16830 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal1 27692 27302 27692 27302 0 mux_bottom_ipin_0.INVTX1_6_.out
rlabel metal2 25254 20332 25254 20332 0 mux_bottom_ipin_0.INVTX1_7_.out
rlabel metal1 21528 20502 21528 20502 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 21206 17204 21206 17204 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 26910 18190 26910 18190 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 29072 36754 29072 36754 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 23506 26282 23506 26282 0 mux_bottom_ipin_1.INVTX1_2_.out
rlabel metal2 17250 20026 17250 20026 0 mux_bottom_ipin_1.INVTX1_3_.out
rlabel metal1 15594 17714 15594 17714 0 mux_bottom_ipin_1.INVTX1_4_.out
rlabel metal1 21804 15538 21804 15538 0 mux_bottom_ipin_1.INVTX1_5_.out
rlabel metal1 24380 23494 24380 23494 0 mux_bottom_ipin_1.INVTX1_6_.out
rlabel metal1 14490 3570 14490 3570 0 mux_bottom_ipin_1.INVTX1_7_.out
rlabel metal2 22218 19312 22218 19312 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20148 14858 20148 14858 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20562 16014 20562 16014 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 30268 30226 30268 30226 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 16698 16762 16698 16762 0 mux_bottom_ipin_2.INVTX1_2_.out
rlabel metal2 28290 15606 28290 15606 0 mux_bottom_ipin_2.INVTX1_3_.out
rlabel metal2 24334 15538 24334 15538 0 mux_bottom_ipin_2.INVTX1_4_.out
rlabel metal1 14030 15402 14030 15402 0 mux_bottom_ipin_2.INVTX1_5_.out
rlabel metal1 20930 27846 20930 27846 0 mux_bottom_ipin_2.INVTX1_6_.out
rlabel metal2 20746 17374 20746 17374 0 mux_bottom_ipin_2.INVTX1_7_.out
rlabel metal1 18676 19278 18676 19278 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15778 15470 15778 15470 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19366 23018 19366 23018 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 13294 27438 13294 27438 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 26036 12750 26036 12750 0 mux_bottom_ipin_3.INVTX1_2_.out
rlabel metal1 22908 9146 22908 9146 0 mux_bottom_ipin_3.INVTX1_3_.out
rlabel metal1 32292 12070 32292 12070 0 mux_bottom_ipin_3.INVTX1_4_.out
rlabel metal1 13984 13362 13984 13362 0 mux_bottom_ipin_3.INVTX1_5_.out
rlabel metal1 26956 22406 26956 22406 0 mux_bottom_ipin_3.INVTX1_6_.out
rlabel metal1 27738 15402 27738 15402 0 mux_bottom_ipin_3.INVTX1_7_.out
rlabel metal1 25392 13838 25392 13838 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20056 14314 20056 14314 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 25714 18836 25714 18836 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 8096 36754 8096 36754 0 mux_bottom_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 15456 12750 15456 12750 0 mux_bottom_ipin_4.INVTX1_2_.out
rlabel metal1 10488 11186 10488 11186 0 mux_bottom_ipin_4.INVTX1_3_.out
rlabel metal1 14076 13838 14076 13838 0 mux_bottom_ipin_4.INVTX1_4_.out
rlabel metal2 12742 10336 12742 10336 0 mux_bottom_ipin_4.INVTX1_5_.out
rlabel metal1 16008 12274 16008 12274 0 mux_bottom_ipin_4.INVTX1_6_.out
rlabel metal2 28750 10370 28750 10370 0 mux_bottom_ipin_4.INVTX1_7_.out
rlabel metal1 18906 12920 18906 12920 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16652 12750 16652 12750 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal3 26864 12444 26864 12444 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 18446 13294 18446 13294 0 mux_bottom_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 12742 13872 12742 13872 0 mux_bottom_ipin_5.INVTX1_2_.out
rlabel metal1 12466 13804 12466 13804 0 mux_bottom_ipin_5.INVTX1_3_.out
rlabel metal1 20470 13838 20470 13838 0 mux_bottom_ipin_5.INVTX1_4_.out
rlabel metal1 12765 13362 12765 13362 0 mux_bottom_ipin_5.INVTX1_5_.out
rlabel metal2 9706 4148 9706 4148 0 mux_bottom_ipin_5.INVTX1_6_.out
rlabel metal2 20746 13090 20746 13090 0 mux_bottom_ipin_5.INVTX1_7_.out
rlabel metal2 11362 9350 11362 9350 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 13018 12716 13018 12716 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15686 11832 15686 11832 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 10166 9588 10166 9588 0 mux_bottom_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 14582 14518 14582 14518 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13478 16864 13478 16864 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 18814 19006 18814 19006 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 7912 27438 7912 27438 0 mux_bottom_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel via2 23966 14909 23966 14909 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 21850 15368 21850 15368 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 21988 13498 21988 13498 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 28106 14994 28106 14994 0 mux_bottom_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 18078 17544 18078 17544 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18423 13430 18423 13430 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 23598 20604 23598 20604 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 25921 29478 25921 29478 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27554 14892 27554 14892 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16652 14518 16652 14518 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 27922 17000 27922 17000 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 29118 17986 29118 17986 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 29854 13464 29854 13464 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20102 12342 20102 12342 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 29992 9962 29992 9962 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 32154 8840 32154 8840 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 12788 12070 12788 12070 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 11454 9554 11454 9554 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 12466 6120 12466 6120 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 14352 12750 14352 12750 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel via3 27485 36516 27485 36516 0 net1
rlabel metal2 2530 2822 2530 2822 0 net10
rlabel metal2 23322 19822 23322 19822 0 net100
rlabel metal1 28612 16082 28612 16082 0 net101
rlabel metal1 26220 12682 26220 12682 0 net102
rlabel metal1 15686 14008 15686 14008 0 net103
rlabel metal2 34546 31552 34546 31552 0 net11
rlabel metal1 25438 26350 25438 26350 0 net12
rlabel metal1 2070 32810 2070 32810 0 net13
rlabel metal1 36156 5202 36156 5202 0 net14
rlabel metal1 2254 36618 2254 36618 0 net15
rlabel metal2 1886 18735 1886 18735 0 net16
rlabel metal1 29624 2482 29624 2482 0 net17
rlabel metal1 8786 17850 8786 17850 0 net18
rlabel metal1 32936 29546 32936 29546 0 net19
rlabel metal1 12880 37298 12880 37298 0 net2
rlabel metal1 32522 2992 32522 2992 0 net20
rlabel metal1 20194 23154 20194 23154 0 net21
rlabel metal1 2622 20230 2622 20230 0 net22
rlabel metal1 1978 29546 1978 29546 0 net23
rlabel metal1 5750 15674 5750 15674 0 net24
rlabel metal1 4876 2550 4876 2550 0 net25
rlabel via2 10810 2363 10810 2363 0 net26
rlabel metal2 28428 2516 28428 2516 0 net27
rlabel metal1 35972 9554 35972 9554 0 net28
rlabel metal1 24564 29478 24564 29478 0 net29
rlabel metal1 16928 37298 16928 37298 0 net3
rlabel metal1 29900 31110 29900 31110 0 net30
rlabel metal1 4393 36074 4393 36074 0 net31
rlabel metal1 25622 20502 25622 20502 0 net32
rlabel via2 1886 8347 1886 8347 0 net33
rlabel metal2 36110 11407 36110 11407 0 net34
rlabel metal1 4738 24106 4738 24106 0 net35
rlabel metal1 20286 15470 20286 15470 0 net36
rlabel metal1 2254 17034 2254 17034 0 net37
rlabel metal1 12926 15504 12926 15504 0 net38
rlabel metal1 2553 12818 2553 12818 0 net39
rlabel metal1 35742 27914 35742 27914 0 net4
rlabel metal1 36202 15096 36202 15096 0 net40
rlabel metal1 35006 37230 35006 37230 0 net41
rlabel metal2 36110 23460 36110 23460 0 net42
rlabel metal2 35374 3026 35374 3026 0 net43
rlabel metal1 14996 3502 14996 3502 0 net44
rlabel metal1 36110 10676 36110 10676 0 net45
rlabel metal1 22494 32538 22494 32538 0 net46
rlabel metal1 2162 36754 2162 36754 0 net47
rlabel metal1 33925 17170 33925 17170 0 net48
rlabel metal2 1886 15878 1886 15878 0 net49
rlabel metal1 2162 37196 2162 37196 0 net5
rlabel metal1 8648 2414 8648 2414 0 net50
rlabel metal2 35926 20162 35926 20162 0 net51
rlabel via2 15686 37077 15686 37077 0 net52
rlabel metal2 36110 8908 36110 8908 0 net53
rlabel metal1 24288 29818 24288 29818 0 net54
rlabel metal1 36018 36686 36018 36686 0 net55
rlabel metal1 34592 2414 34592 2414 0 net56
rlabel metal1 18492 37230 18492 37230 0 net57
rlabel metal1 31280 3910 31280 3910 0 net58
rlabel metal2 7866 4794 7866 4794 0 net59
rlabel metal1 24104 23698 24104 23698 0 net6
rlabel metal1 10488 2414 10488 2414 0 net60
rlabel metal2 2392 21420 2392 21420 0 net61
rlabel metal1 33925 16082 33925 16082 0 net62
rlabel metal1 5152 2414 5152 2414 0 net63
rlabel metal1 2024 12954 2024 12954 0 net64
rlabel metal2 9614 7548 9614 7548 0 net65
rlabel metal2 2438 3213 2438 3213 0 net66
rlabel metal1 30544 12614 30544 12614 0 net67
rlabel metal2 12098 37060 12098 37060 0 net68
rlabel metal1 21528 35258 21528 35258 0 net69
rlabel metal1 19872 37230 19872 37230 0 net7
rlabel metal2 27370 37026 27370 37026 0 net70
rlabel metal1 2162 26350 2162 26350 0 net71
rlabel metal1 2254 19686 2254 19686 0 net72
rlabel metal2 1886 2618 1886 2618 0 net73
rlabel metal2 36110 36516 36110 36516 0 net74
rlabel metal1 27922 35802 27922 35802 0 net75
rlabel metal2 15088 14382 15088 14382 0 net76
rlabel metal1 35144 36754 35144 36754 0 net77
rlabel via2 35926 3995 35926 3995 0 net78
rlabel metal2 1886 11356 1886 11356 0 net79
rlabel metal1 27600 22610 27600 22610 0 net8
rlabel metal1 34316 22610 34316 22610 0 net80
rlabel metal2 6578 5066 6578 5066 0 net81
rlabel metal2 7406 2176 7406 2176 0 net82
rlabel metal1 19274 3536 19274 3536 0 net83
rlabel metal1 30452 36890 30452 36890 0 net84
rlabel metal1 29992 37230 29992 37230 0 net85
rlabel metal1 3496 37230 3496 37230 0 net86
rlabel metal2 7682 37060 7682 37060 0 net87
rlabel metal2 26542 4420 26542 4420 0 net88
rlabel metal2 8786 11254 8786 11254 0 net89
rlabel metal2 2714 12920 2714 12920 0 net9
rlabel metal2 7590 31314 7590 31314 0 net90
rlabel metal2 36110 17510 36110 17510 0 net91
rlabel metal1 27140 19482 27140 19482 0 net92
rlabel metal1 23184 16626 23184 16626 0 net93
rlabel metal2 15318 21726 15318 21726 0 net94
rlabel metal2 24058 18530 24058 18530 0 net95
rlabel metal2 18538 10336 18538 10336 0 net96
rlabel metal1 8004 10778 8004 10778 0 net97
rlabel metal1 21022 20570 21022 20570 0 net98
rlabel metal1 22264 11866 22264 11866 0 net99
rlabel metal2 36386 24021 36386 24021 0 pReset
rlabel metal1 20930 5542 20930 5542 0 prog_clk
rlabel metal1 31096 37094 31096 37094 0 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 29762 37094 29762 37094 0 top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 3266 38158 3266 38158 0 top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 7912 37094 7912 37094 0 top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 27048 3706 27048 3706 0 top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal3 1188 11628 1188 11628 0 top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal3 1188 34748 1188 34748 0 top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_
rlabel via2 36294 19125 36294 19125 0 top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 38000 40000
<< end >>
